//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1273,
    new_n1274, new_n1275, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n211), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n221), .A2(new_n208), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT64), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n216), .B(new_n225), .C1(new_n223), .C2(new_n222), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G58), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G97), .B(G107), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  AND2_X1   g0043(.A1(G1), .A2(G13), .ZN(new_n244));
  NAND2_X1  g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G274), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AND2_X1   g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(new_n212), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n255), .A2(G226), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G223), .A3(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G77), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G222), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n258), .B1(new_n259), .B2(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n244), .A2(KEYINPUT66), .A3(new_n245), .ZN(new_n264));
  AOI21_X1  g0064(.A(KEYINPUT66), .B1(new_n244), .B2(new_n245), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI211_X1 g0066(.A(new_n249), .B(new_n256), .C1(new_n263), .C2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G179), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G20), .A2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G150), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n206), .A2(G33), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT8), .B(G58), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n270), .B(new_n272), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n212), .ZN(new_n277));
  INV_X1    g0077(.A(G50), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n275), .A2(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n276), .A2(new_n212), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n279), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT67), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n283), .A2(new_n284), .B1(new_n205), .B2(G20), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n280), .A2(new_n277), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n281), .B1(new_n288), .B2(new_n278), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n269), .B(new_n289), .C1(G169), .C2(new_n267), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT10), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT9), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g0094(.A(new_n294), .B(KEYINPUT68), .Z(new_n295));
  NAND2_X1  g0095(.A1(new_n267), .A2(G190), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(new_n267), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(new_n293), .B2(new_n289), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n292), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n295), .A2(new_n299), .A3(new_n292), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n291), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G58), .ZN(new_n304));
  INV_X1    g0104(.A(G68), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(G20), .B1(new_n306), .B2(new_n201), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n271), .A2(G159), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OR2_X1    g0109(.A1(KEYINPUT3), .A2(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(KEYINPUT3), .A2(G33), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n310), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT71), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  NOR2_X1   g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n317), .A2(KEYINPUT71), .A3(KEYINPUT7), .A4(new_n206), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT7), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n257), .B2(G20), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n314), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n309), .B1(new_n321), .B2(G68), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n282), .B1(new_n322), .B2(KEYINPUT16), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT16), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n305), .B1(new_n320), .B2(new_n312), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(new_n309), .ZN(new_n326));
  INV_X1    g0126(.A(new_n274), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n288), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n274), .A2(new_n279), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n323), .A2(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n264), .A2(new_n265), .ZN(new_n331));
  OAI211_X1 g0131(.A(G223), .B(new_n260), .C1(new_n315), .C2(new_n316), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT72), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT72), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n257), .A2(new_n334), .A3(G223), .A4(new_n260), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g0136(.A(G226), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G87), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n331), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n246), .A2(G232), .A3(new_n248), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT73), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT73), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n246), .A2(new_n344), .A3(G232), .A4(new_n248), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n249), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(G169), .B1(new_n341), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n249), .B1(new_n343), .B2(new_n345), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n339), .B1(new_n335), .B2(new_n333), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n350), .B(G179), .C1(new_n351), .C2(new_n331), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT18), .B1(new_n330), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n297), .B1(new_n341), .B2(new_n348), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n350), .B(new_n356), .C1(new_n351), .C2(new_n331), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n321), .A2(G68), .ZN(new_n359));
  INV_X1    g0159(.A(new_n309), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(KEYINPUT16), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(new_n277), .A3(new_n326), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n328), .A2(new_n329), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n358), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT17), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n362), .A2(new_n363), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT18), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n349), .A2(new_n352), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n330), .A2(KEYINPUT17), .A3(new_n358), .ZN(new_n371));
  AND4_X1   g0171(.A1(new_n354), .A2(new_n366), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n271), .A2(G50), .B1(G20), .B2(new_n305), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n259), .B2(new_n273), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n277), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT11), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n280), .A2(new_n305), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT12), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n374), .A2(KEYINPUT11), .A3(new_n277), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n286), .B(G68), .C1(G1), .C2(new_n206), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n377), .A2(new_n379), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n382), .A2(KEYINPUT69), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(KEYINPUT69), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT13), .ZN(new_n386));
  INV_X1    g0186(.A(new_n247), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(new_n254), .B1(new_n255), .B2(G238), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G97), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n229), .A2(G1698), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(G226), .B2(G1698), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n389), .B1(new_n391), .B2(new_n317), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n266), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n386), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n388), .A2(new_n386), .A3(new_n393), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G200), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n385), .B(new_n398), .C1(new_n397), .C2(new_n356), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n395), .A2(G179), .A3(new_n396), .ZN(new_n401));
  INV_X1    g0201(.A(new_n396), .ZN(new_n402));
  OAI21_X1  g0202(.A(G169), .B1(new_n402), .B2(new_n394), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n401), .B1(new_n403), .B2(KEYINPUT14), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT70), .ZN(new_n405));
  INV_X1    g0205(.A(G169), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n395), .B2(new_n396), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT14), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n403), .A2(KEYINPUT70), .A3(KEYINPUT14), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n404), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n385), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n400), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n327), .A2(new_n271), .B1(G20), .B2(G77), .ZN(new_n415));
  XOR2_X1   g0215(.A(KEYINPUT15), .B(G87), .Z(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n415), .B1(new_n273), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n277), .ZN(new_n419));
  OAI21_X1  g0219(.A(G77), .B1(new_n206), .B2(G1), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n419), .B1(G77), .B2(new_n279), .C1(new_n283), .C2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n257), .A2(G238), .A3(G1698), .ZN(new_n422));
  INV_X1    g0222(.A(G107), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n422), .B1(new_n423), .B2(new_n257), .C1(new_n261), .C2(new_n229), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n266), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n249), .B1(G244), .B2(new_n255), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n421), .B1(G190), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n297), .B2(new_n428), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n406), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n421), .B(new_n431), .C1(G179), .C2(new_n427), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n303), .A2(new_n372), .A3(new_n414), .A4(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n253), .A2(G1), .ZN(new_n436));
  AND2_X1   g0236(.A1(KEYINPUT5), .A2(G41), .ZN(new_n437));
  NOR2_X1   g0237(.A1(KEYINPUT5), .A2(G41), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n439), .A2(G270), .A3(new_n246), .ZN(new_n440));
  XNOR2_X1  g0240(.A(KEYINPUT5), .B(G41), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n441), .A2(new_n246), .A3(G274), .A4(new_n436), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT79), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n440), .A2(KEYINPUT79), .A3(new_n442), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(G264), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT80), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n257), .A2(KEYINPUT80), .A3(G264), .A4(G1698), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n317), .A2(G303), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n257), .A2(G257), .A3(new_n260), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n454), .A2(KEYINPUT81), .A3(new_n266), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n447), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT81), .B1(new_n454), .B2(new_n266), .ZN(new_n457));
  OAI21_X1  g0257(.A(G200), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G33), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n282), .B(new_n279), .C1(G1), .C2(new_n459), .ZN(new_n460));
  MUX2_X1   g0260(.A(new_n279), .B(new_n460), .S(G116), .Z(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  INV_X1    g0262(.A(G97), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n206), .C1(G33), .C2(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n277), .C1(new_n206), .C2(G116), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT20), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n454), .A2(new_n266), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT81), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n472), .A2(G190), .A3(new_n455), .A4(new_n447), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n458), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n455), .A3(new_n447), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n406), .B1(new_n461), .B2(new_n467), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT21), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n456), .A2(new_n457), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(G179), .A3(new_n468), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n475), .A2(KEYINPUT21), .A3(new_n476), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n474), .A2(new_n479), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n206), .B(G87), .C1(new_n315), .C2(new_n316), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT82), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT22), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(KEYINPUT22), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n257), .A2(new_n206), .A3(G87), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G116), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT83), .B1(new_n490), .B2(G20), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT83), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(new_n206), .A3(G33), .A4(G116), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI22_X1  g0294(.A1(new_n206), .A2(G107), .B1(KEYINPUT84), .B2(KEYINPUT23), .ZN(new_n495));
  AND2_X1   g0295(.A1(KEYINPUT84), .A2(KEYINPUT23), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n423), .A2(G20), .ZN(new_n497));
  OAI22_X1  g0297(.A1(new_n495), .A2(new_n496), .B1(KEYINPUT23), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n489), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT85), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT85), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n489), .A2(new_n502), .A3(new_n499), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(KEYINPUT24), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n502), .B1(new_n489), .B2(new_n499), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT24), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n282), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n280), .A2(KEYINPUT25), .A3(new_n423), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT25), .B1(new_n280), .B2(new_n423), .ZN(new_n511));
  OAI22_X1  g0311(.A1(new_n510), .A2(new_n511), .B1(new_n460), .B2(new_n423), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(G257), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n514));
  OAI211_X1 g0314(.A(G250), .B(new_n260), .C1(new_n315), .C2(new_n316), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G294), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n441), .A2(new_n436), .B1(new_n244), .B2(new_n245), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n517), .A2(new_n266), .B1(new_n518), .B2(G264), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n442), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n297), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n356), .A3(new_n442), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n508), .A2(new_n513), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n512), .B1(new_n504), .B2(new_n507), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n520), .A2(new_n406), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(G179), .B2(new_n520), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n271), .A2(G77), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT74), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n271), .A2(KEYINPUT74), .A3(G77), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT6), .ZN(new_n534));
  AND2_X1   g0334(.A1(G97), .A2(G107), .ZN(new_n535));
  NOR2_X1   g0335(.A1(G97), .A2(G107), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n423), .A2(KEYINPUT6), .A3(G97), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n533), .B1(new_n539), .B2(G20), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT7), .B1(new_n317), .B2(new_n206), .ZN(new_n541));
  INV_X1    g0341(.A(new_n312), .ZN(new_n542));
  OAI21_X1  g0342(.A(G107), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n282), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n280), .A2(new_n463), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n460), .B2(new_n463), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT75), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n534), .A2(new_n463), .A3(G107), .ZN(new_n548));
  XNOR2_X1  g0348(.A(G97), .B(G107), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n534), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n532), .B(new_n531), .C1(new_n550), .C2(new_n206), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n423), .B1(new_n320), .B2(new_n312), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n277), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT75), .ZN(new_n554));
  INV_X1    g0354(.A(new_n546), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n439), .A2(new_n246), .ZN(new_n557));
  INV_X1    g0357(.A(G257), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n442), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(G244), .B(new_n260), .C1(new_n315), .C2(new_n316), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT4), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(KEYINPUT76), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(KEYINPUT76), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n257), .A2(G244), .A3(new_n260), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n562), .A2(new_n462), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  AOI211_X1 g0366(.A(G190), .B(new_n559), .C1(new_n266), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n266), .ZN(new_n568));
  INV_X1    g0368(.A(new_n559), .ZN(new_n569));
  AOI21_X1  g0369(.A(G200), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n547), .B(new_n556), .C1(new_n567), .C2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n416), .A2(new_n279), .ZN(new_n572));
  INV_X1    g0372(.A(G87), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n460), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g0374(.A(KEYINPUT78), .B(G87), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n536), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT19), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n206), .B1(new_n389), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n257), .A2(new_n206), .A3(G68), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n577), .B1(new_n273), .B2(new_n463), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI211_X1 g0382(.A(new_n572), .B(new_n574), .C1(new_n582), .C2(new_n277), .ZN(new_n583));
  INV_X1    g0383(.A(G238), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n260), .ZN(new_n585));
  INV_X1    g0385(.A(G244), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G1698), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n585), .B(new_n587), .C1(new_n315), .C2(new_n316), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n490), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT77), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT77), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(new_n591), .A3(new_n490), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n266), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G250), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n251), .A2(new_n594), .A3(new_n436), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n595), .B1(new_n436), .B2(new_n387), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G200), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n583), .B(new_n598), .C1(new_n356), .C2(new_n597), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n553), .A2(new_n555), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n559), .B1(new_n566), .B2(new_n266), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n406), .ZN(new_n602));
  AOI211_X1 g0402(.A(new_n268), .B(new_n559), .C1(new_n266), .C2(new_n566), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n572), .B1(new_n582), .B2(new_n277), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n460), .B2(new_n417), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n597), .A2(new_n406), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n593), .A2(new_n268), .A3(new_n596), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n571), .A2(new_n599), .A3(new_n604), .A4(new_n609), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n483), .A2(new_n528), .A3(new_n610), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n435), .A2(new_n611), .ZN(G372));
  INV_X1    g0412(.A(new_n432), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n412), .A2(new_n413), .B1(new_n399), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n366), .A2(new_n371), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n354), .B(new_n370), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT88), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n616), .A2(new_n617), .B1(new_n301), .B2(new_n302), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n291), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n508), .A2(new_n513), .ZN(new_n621));
  INV_X1    g0421(.A(new_n527), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT86), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT86), .B1(new_n525), .B2(new_n527), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT87), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n524), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n610), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n626), .A2(new_n627), .A3(KEYINPUT87), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n630), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n599), .A2(new_n609), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n602), .A2(new_n603), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n547), .A2(new_n556), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n609), .B1(new_n640), .B2(KEYINPUT26), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  INV_X1    g0442(.A(new_n604), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n636), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n634), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n435), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n620), .A2(new_n647), .ZN(G369));
  INV_X1    g0448(.A(new_n627), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n469), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n649), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n483), .B2(new_n657), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n528), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n525), .B2(new_n656), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n525), .A2(new_n527), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n663), .B1(new_n665), .B2(new_n656), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n627), .A2(new_n655), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n662), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n624), .A2(new_n625), .A3(new_n656), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT89), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(KEYINPUT89), .A3(new_n670), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n667), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n209), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n576), .A2(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n214), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n609), .B(KEYINPUT93), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n627), .A2(new_n665), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(new_n632), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n642), .B1(new_n635), .B2(new_n604), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT94), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n636), .A2(KEYINPUT26), .A3(new_n638), .A4(new_n639), .ZN(new_n690));
  OAI211_X1 g0490(.A(KEYINPUT94), .B(new_n642), .C1(new_n635), .C2(new_n604), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n655), .B1(new_n686), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT29), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n655), .B1(new_n634), .B2(new_n645), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n695), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G330), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT92), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n472), .A2(G179), .A3(new_n455), .A4(new_n447), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n593), .A2(new_n519), .A3(new_n596), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT90), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n593), .A2(KEYINPUT90), .A3(new_n519), .A4(new_n596), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT30), .B1(new_n705), .B2(new_n601), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT91), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n601), .B1(new_n597), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(G179), .B1(new_n519), .B2(new_n442), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n593), .A2(KEYINPUT91), .A3(new_n596), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n708), .A2(new_n475), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n699), .B1(new_n706), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n700), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n703), .A2(new_n704), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n601), .A2(KEYINPUT30), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n706), .A2(new_n699), .A3(new_n712), .ZN(new_n719));
  OAI211_X1 g0519(.A(KEYINPUT31), .B(new_n655), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n711), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n655), .B1(new_n706), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n611), .A2(new_n656), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n698), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n697), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n683), .B1(new_n728), .B2(G1), .ZN(G364));
  INV_X1    g0529(.A(G13), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n205), .B1(new_n731), .B2(G45), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n678), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n661), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(G330), .B2(new_n659), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n677), .A2(new_n317), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G355), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(G116), .B2(new_n209), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n677), .A2(new_n257), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n253), .B2(new_n215), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n239), .A2(new_n253), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n739), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n244), .B1(new_n206), .B2(G169), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n745), .A2(KEYINPUT95), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(KEYINPUT95), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n734), .B1(new_n744), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n206), .A2(new_n268), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT98), .Z(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n356), .A2(G179), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n206), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n758), .A2(G326), .B1(G294), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT99), .Z(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n755), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n206), .A2(G179), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n764), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G311), .A2(new_n765), .B1(new_n768), .B2(G329), .ZN(new_n769));
  INV_X1    g0569(.A(G322), .ZN(new_n770));
  NOR4_X1   g0570(.A1(new_n206), .A2(new_n268), .A3(new_n356), .A4(G200), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n769), .B(new_n317), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G283), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n766), .A2(new_n356), .A3(G200), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n766), .A2(G190), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(G303), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n755), .A2(new_n356), .A3(G200), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n780), .A2(KEYINPUT97), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(KEYINPUT97), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(KEYINPUT33), .B(G317), .Z(new_n784));
  OAI21_X1  g0584(.A(new_n779), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n765), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n259), .A2(new_n786), .B1(new_n772), .B2(new_n304), .ZN(new_n787));
  INV_X1    g0587(.A(new_n756), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G50), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT32), .ZN(new_n790));
  INV_X1    g0590(.A(G159), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n767), .A2(new_n791), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n789), .B1(new_n790), .B2(new_n792), .C1(new_n463), .C2(new_n760), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n787), .B(new_n793), .C1(new_n790), .C2(new_n792), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n305), .B2(new_n783), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n257), .B1(new_n775), .B2(new_n423), .C1(new_n575), .C2(new_n776), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT96), .Z(new_n797));
  OAI22_X1  g0597(.A1(new_n763), .A2(new_n785), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n754), .B1(new_n798), .B2(new_n748), .ZN(new_n799));
  INV_X1    g0599(.A(new_n751), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n659), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n736), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  NAND2_X1  g0603(.A1(new_n613), .A2(KEYINPUT101), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT101), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n432), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n807), .A2(new_n430), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n646), .A2(new_n656), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n421), .A2(new_n655), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n804), .A2(new_n430), .A3(new_n810), .A4(new_n806), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n613), .A2(new_n655), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n809), .B1(new_n696), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n734), .B1(new_n814), .B2(new_n726), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n726), .B2(new_n814), .ZN(new_n816));
  INV_X1    g0616(.A(new_n748), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n750), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n734), .B1(new_n818), .B2(G77), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT100), .Z(new_n820));
  INV_X1    g0620(.A(G116), .ZN(new_n821));
  INV_X1    g0621(.A(G294), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n821), .A2(new_n786), .B1(new_n772), .B2(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n257), .B(new_n823), .C1(G311), .C2(new_n768), .ZN(new_n824));
  INV_X1    g0624(.A(new_n783), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(G283), .ZN(new_n826));
  INV_X1    g0626(.A(new_n776), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n761), .A2(G97), .B1(new_n827), .B2(G107), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n775), .A2(new_n573), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G303), .B2(new_n788), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n824), .A2(new_n826), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n257), .B1(new_n767), .B2(new_n832), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n278), .A2(new_n776), .B1(new_n775), .B2(new_n305), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n833), .B(new_n834), .C1(G58), .C2(new_n761), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G159), .A2(new_n765), .B1(new_n771), .B2(G143), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  INV_X1    g0637(.A(G150), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n836), .B1(new_n837), .B2(new_n756), .C1(new_n783), .C2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n835), .B1(new_n840), .B2(KEYINPUT34), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT34), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n831), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n820), .B1(new_n844), .B2(new_n748), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n813), .B2(new_n750), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n816), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G384));
  NOR2_X1   g0648(.A1(new_n731), .A2(new_n205), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT40), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n354), .A2(new_n366), .A3(new_n370), .A4(new_n371), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n361), .A2(new_n277), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n322), .A2(KEYINPUT16), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n363), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT104), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n653), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n363), .B(KEYINPUT104), .C1(new_n852), .C2(new_n853), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT105), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n851), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n860), .B1(new_n851), .B2(new_n859), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n856), .A2(new_n369), .A3(new_n858), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n864), .A2(new_n865), .A3(new_n364), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n362), .A2(new_n363), .B1(new_n349), .B2(new_n352), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n330), .B2(new_n358), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT106), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n367), .A2(new_n857), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n367), .A2(new_n369), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n873), .A2(new_n871), .A3(new_n870), .A4(new_n364), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT106), .ZN(new_n875));
  AOI22_X1  g0675(.A1(KEYINPUT37), .A2(new_n866), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n863), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT105), .B1(new_n372), .B2(new_n864), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n851), .A2(new_n859), .A3(new_n860), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n872), .A2(new_n875), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT38), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n878), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n383), .A2(new_n384), .A3(new_n655), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n399), .B1(new_n411), .B2(new_n385), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT103), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n889), .B(new_n399), .C1(new_n411), .C2(new_n385), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n887), .B(new_n404), .C1(new_n409), .C2(new_n410), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n890), .A2(new_n893), .A3(new_n813), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(KEYINPUT31), .B(new_n655), .C1(new_n706), .C2(new_n721), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT107), .B1(new_n724), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n722), .A2(new_n723), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n528), .A2(new_n610), .ZN(new_n899));
  AND4_X1   g0699(.A1(new_n479), .A2(new_n474), .A3(new_n481), .A4(new_n482), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(new_n900), .A3(new_n656), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n898), .A2(new_n901), .A3(KEYINPUT107), .A4(new_n896), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n895), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n850), .B1(new_n886), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT108), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n877), .B1(new_n863), .B2(new_n876), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n881), .A2(KEYINPUT38), .A3(new_n884), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n898), .A2(new_n901), .A3(new_n896), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT107), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n894), .B1(new_n912), .B2(new_n902), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT108), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(new_n915), .A3(new_n850), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n906), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n913), .A2(KEYINPUT109), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n912), .A2(new_n902), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(KEYINPUT109), .A3(new_n895), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n870), .B1(new_n868), .B2(new_n871), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n872), .B2(new_n875), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n372), .A2(new_n871), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n877), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n850), .B1(new_n908), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n917), .B1(new_n918), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n435), .A2(new_n919), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(G330), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n927), .B2(new_n928), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n908), .A2(new_n924), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n908), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n411), .A2(new_n385), .A3(new_n655), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n857), .B1(new_n354), .B2(new_n370), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n807), .A2(new_n655), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n696), .B2(new_n808), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n890), .A2(new_n893), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n941), .B1(new_n945), .B2(new_n909), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n620), .B1(new_n697), .B2(new_n434), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n947), .B(new_n948), .Z(new_n949));
  AOI21_X1  g0749(.A(new_n849), .B1(new_n932), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n932), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n539), .A2(KEYINPUT35), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n539), .A2(KEYINPUT35), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n952), .A2(new_n953), .A3(G116), .A4(new_n213), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT36), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n214), .A2(new_n259), .A3(new_n306), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n956), .A2(KEYINPUT102), .B1(new_n278), .B2(G68), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(KEYINPUT102), .B2(new_n956), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n958), .A2(G1), .A3(new_n730), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n951), .A2(new_n955), .A3(new_n959), .ZN(G367));
  OR2_X1    g0760(.A1(new_n583), .A2(new_n656), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n636), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n609), .B2(new_n961), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(new_n800), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n752), .B1(new_n209), .B2(new_n417), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n741), .A2(new_n235), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n734), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G283), .A2(new_n765), .B1(new_n771), .B2(G303), .ZN(new_n968));
  INV_X1    g0768(.A(G317), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n968), .B(new_n317), .C1(new_n969), .C2(new_n767), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n760), .A2(new_n423), .B1(new_n775), .B2(new_n463), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n776), .A2(new_n821), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(KEYINPUT46), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(KEYINPUT46), .ZN(new_n974));
  NOR4_X1   g0774(.A1(new_n970), .A2(new_n971), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n758), .A2(G311), .B1(new_n825), .B2(G294), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n758), .A2(G143), .B1(new_n825), .B2(G159), .ZN(new_n977));
  INV_X1    g0777(.A(new_n775), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n761), .A2(G68), .B1(new_n978), .B2(G77), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n304), .B2(new_n776), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n257), .B1(new_n772), .B2(new_n838), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n786), .A2(new_n278), .B1(new_n767), .B2(new_n837), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n975), .A2(new_n976), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(KEYINPUT47), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n817), .B1(new_n984), .B2(KEYINPUT47), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n967), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n964), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n639), .A2(new_n655), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n989), .A2(new_n604), .A3(new_n571), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n638), .A2(new_n639), .A3(new_n655), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n674), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT89), .B1(new_n669), .B2(new_n670), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT45), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n675), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n992), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n673), .A2(new_n674), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT44), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n673), .A2(KEYINPUT44), .A3(new_n674), .A4(new_n1000), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AND3_X1   g0805(.A1(new_n999), .A2(new_n667), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n667), .B1(new_n999), .B2(new_n1005), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n669), .B1(new_n666), .B2(new_n668), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(new_n660), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n727), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(KEYINPUT111), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n999), .A2(new_n1005), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n667), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n999), .A2(new_n667), .A3(new_n1005), .ZN(new_n1016));
  AND4_X1   g0816(.A1(KEYINPUT111), .A2(new_n1015), .A3(new_n1011), .A4(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n728), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n678), .B(KEYINPUT41), .Z(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n733), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n668), .A2(new_n662), .A3(new_n992), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT42), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(KEYINPUT42), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n643), .B1(new_n992), .B2(new_n664), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1023), .B(new_n1024), .C1(new_n1025), .C2(new_n655), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1026), .A2(KEYINPUT110), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n963), .B(KEYINPUT43), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(KEYINPUT110), .ZN(new_n1029));
  AND3_X1   g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n667), .A2(new_n1000), .ZN(new_n1033));
  OR3_X1    g0833(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n988), .B1(new_n1021), .B2(new_n1036), .ZN(G387));
  INV_X1    g0837(.A(new_n1011), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n727), .A2(new_n1010), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n678), .A3(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G303), .A2(new_n765), .B1(new_n771), .B2(G317), .ZN(new_n1041));
  INV_X1    g0841(.A(G311), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1041), .B1(new_n783), .B2(new_n1042), .C1(new_n757), .C2(new_n770), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT112), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n760), .A2(new_n774), .B1(new_n776), .B2(new_n822), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT49), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(KEYINPUT49), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n775), .A2(new_n821), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n257), .B(new_n1052), .C1(G326), .C2(new_n768), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n305), .A2(new_n786), .B1(new_n772), .B2(new_n278), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n317), .B(new_n1055), .C1(G150), .C2(new_n768), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n825), .A2(new_n327), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n776), .A2(new_n259), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G97), .B2(new_n978), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n416), .A2(new_n761), .B1(new_n788), .B2(G159), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n817), .B1(new_n1054), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n740), .B1(new_n232), .B2(new_n253), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n737), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n680), .B2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n680), .B(new_n253), .C1(new_n305), .C2(new_n259), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT50), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n327), .B2(new_n278), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n274), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1065), .A2(new_n1071), .B1(new_n423), .B2(new_n677), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n734), .B1(new_n1072), .B2(new_n753), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1062), .A2(KEYINPUT113), .A3(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n666), .A2(new_n800), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(KEYINPUT113), .B1(new_n1062), .B2(new_n1073), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1040), .B(new_n1079), .C1(new_n732), .C2(new_n1010), .ZN(G393));
  NAND2_X1  g0880(.A1(new_n1008), .A2(new_n733), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n992), .A2(new_n800), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT114), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n753), .B1(G97), .B2(new_n677), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n740), .A2(new_n242), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n678), .B(new_n733), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n829), .B1(G68), .B2(new_n827), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n259), .B2(new_n760), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n317), .B1(new_n768), .B2(G143), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n274), .B2(new_n786), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n772), .A2(new_n791), .B1(new_n756), .B2(new_n838), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT51), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1091), .B(new_n1093), .C1(new_n278), .C2(new_n783), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n788), .A2(G317), .B1(new_n771), .B2(G311), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT52), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n317), .B1(new_n786), .B2(new_n822), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G322), .B2(new_n768), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n423), .A2(new_n775), .B1(new_n776), .B2(new_n774), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G116), .B2(new_n761), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(new_n777), .C2(new_n783), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1094), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1102), .A2(KEYINPUT115), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n748), .B1(new_n1102), .B2(KEYINPUT115), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1083), .B(new_n1086), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1081), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n679), .B1(new_n1108), .B2(new_n1038), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1110), .A2(KEYINPUT116), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT116), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT111), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1108), .B2(new_n1038), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1008), .A2(KEYINPUT111), .A3(new_n1011), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1112), .B1(new_n1116), .B2(new_n1109), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1107), .B1(new_n1111), .B2(new_n1117), .ZN(G390));
  AOI21_X1  g0918(.A(new_n698), .B1(new_n912), .B2(new_n902), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n895), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n942), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n809), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n944), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n939), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1125), .A2(new_n1126), .B1(new_n935), .B2(new_n936), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n942), .B1(new_n693), .B2(new_n808), .ZN(new_n1128));
  OR2_X1    g0928(.A1(new_n1128), .A2(new_n944), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1129), .A2(new_n1126), .A3(new_n933), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1121), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n937), .B1(new_n945), .B2(new_n939), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n725), .A2(new_n813), .A3(new_n1124), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1129), .A2(new_n1126), .A3(new_n933), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1131), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n725), .A2(new_n813), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n944), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n1120), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n1123), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1119), .A2(new_n813), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n944), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n1128), .A3(new_n1133), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1119), .A2(new_n435), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n620), .B(new_n1145), .C1(new_n697), .C2(new_n434), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1136), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1131), .A2(new_n1147), .A3(new_n1144), .A4(new_n1135), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n678), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1131), .A2(new_n733), .A3(new_n1135), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT119), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n734), .B1(new_n818), .B2(new_n327), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n825), .A2(G137), .B1(new_n765), .B2(new_n1156), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1157), .A2(KEYINPUT117), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n257), .B1(new_n772), .B2(new_n832), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n761), .A2(G159), .B1(new_n978), .B2(G50), .ZN(new_n1160));
  INV_X1    g0960(.A(G128), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1160), .B1(new_n1161), .B2(new_n756), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1159), .B(new_n1162), .C1(G125), .C2(new_n768), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1157), .A2(KEYINPUT117), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n776), .A2(new_n838), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT53), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1158), .A2(new_n1163), .A3(new_n1164), .A4(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n783), .A2(new_n423), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n761), .A2(G77), .B1(new_n978), .B2(G68), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G283), .A2(new_n788), .B1(new_n827), .B2(G87), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n257), .B1(new_n768), .B2(G294), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G97), .A2(new_n765), .B1(new_n771), .B2(G116), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1167), .B1(new_n1168), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1174), .A2(KEYINPUT118), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1175), .A2(new_n817), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(KEYINPUT118), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1154), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n938), .B2(new_n750), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1152), .A2(new_n1153), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1153), .B1(new_n1152), .B2(new_n1179), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1151), .B1(new_n1180), .B2(new_n1181), .ZN(G378));
  INV_X1    g0982(.A(new_n947), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n915), .B1(new_n914), .B2(new_n850), .ZN(new_n1184));
  AOI211_X1 g0984(.A(KEYINPUT108), .B(KEYINPUT40), .C1(new_n909), .C2(new_n913), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(G330), .B1(new_n926), .B2(new_n918), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n289), .A2(new_n857), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n303), .B(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1186), .A2(new_n1187), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1191), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n920), .A2(new_n925), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n918), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n698), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1193), .B1(new_n917), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1183), .B1(new_n1192), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1191), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n917), .A2(new_n1196), .A3(new_n1193), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n1200), .A3(new_n947), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1198), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1191), .A2(new_n749), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n734), .B1(new_n818), .B2(G50), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(G33), .A2(G41), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT120), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G50), .B(new_n1206), .C1(new_n252), .C2(new_n317), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n978), .A2(G58), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n821), .B2(new_n756), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1058), .B(new_n1209), .C1(G68), .C2(new_n761), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n825), .A2(G97), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G41), .B(new_n257), .C1(new_n768), .C2(G283), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n416), .A2(new_n765), .B1(new_n771), .B2(G107), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT58), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1207), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n837), .A2(new_n786), .B1(new_n772), .B2(new_n1161), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G150), .B2(new_n761), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n788), .A2(G125), .B1(new_n827), .B2(new_n1156), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n783), .C2(new_n832), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(KEYINPUT59), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(KEYINPUT59), .ZN(new_n1222));
  INV_X1    g1022(.A(G124), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1206), .B1(new_n1223), .B2(new_n767), .C1(new_n791), .C2(new_n775), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT121), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1216), .B1(new_n1215), .B2(new_n1214), .C1(new_n1221), .C2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1204), .B1(new_n1227), .B2(new_n748), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1202), .A2(new_n733), .B1(new_n1203), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1150), .A2(new_n1147), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1199), .A2(new_n947), .A3(new_n1200), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n947), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1232));
  OAI211_X1 g1032(.A(KEYINPUT57), .B(new_n1230), .C1(new_n1231), .C2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n678), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1202), .B2(new_n1230), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1229), .B1(new_n1234), .B2(new_n1235), .ZN(G375));
  OAI21_X1  g1036(.A(new_n734), .B1(new_n818), .B2(G68), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n786), .A2(new_n423), .B1(new_n767), .B2(new_n777), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n257), .B(new_n1238), .C1(G283), .C2(new_n771), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n825), .A2(G116), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n761), .A2(new_n416), .B1(new_n978), .B2(G77), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G294), .A2(new_n788), .B1(new_n827), .B2(G97), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1208), .B1(new_n278), .B2(new_n760), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n257), .B1(new_n1161), .B2(new_n767), .C1(new_n786), .C2(new_n838), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(G159), .C2(new_n827), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n772), .A2(new_n837), .B1(new_n756), .B2(new_n832), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n825), .B2(new_n1156), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT123), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1246), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1248), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1251), .A2(KEYINPUT123), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1243), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1237), .B1(new_n1253), .B2(new_n748), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1124), .B2(new_n750), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1255), .B1(new_n1256), .B2(new_n732), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT122), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1256), .A2(new_n1259), .A3(new_n1146), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1140), .A2(new_n1143), .A3(new_n1146), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT122), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1148), .A2(new_n1020), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1258), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT124), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(G381));
  NOR2_X1   g1067(.A1(G381), .A2(G387), .ZN(new_n1268));
  INV_X1    g1068(.A(G375), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1151), .A2(new_n1152), .A3(new_n1179), .ZN(new_n1270));
  NOR4_X1   g1070(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .A4(new_n1271), .ZN(G407));
  NAND2_X1  g1072(.A1(new_n654), .A2(G213), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1269), .A2(new_n1270), .A3(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(G407), .A2(G213), .A3(new_n1275), .ZN(G409));
  AOI21_X1  g1076(.A(new_n727), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n732), .B1(new_n1277), .B2(new_n1019), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1036), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(G390), .A2(new_n988), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1110), .A2(KEYINPUT116), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1116), .A2(new_n1112), .A3(new_n1109), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1106), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G387), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(G393), .B(new_n802), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1281), .A2(new_n1285), .A3(new_n1286), .A4(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT125), .B1(G387), .B2(new_n1284), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1290), .A2(new_n1287), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G378), .B(new_n1229), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1202), .A2(new_n1020), .A3(new_n1230), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n733), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1203), .A2(new_n1228), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1270), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1294), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1273), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1148), .A2(KEYINPUT60), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(new_n1260), .A3(new_n1262), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1261), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n679), .B1(new_n1304), .B2(KEYINPUT60), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(G384), .B1(new_n1306), .B2(new_n1258), .ZN(new_n1307));
  AOI211_X1 g1107(.A(new_n847), .B(new_n1257), .C1(new_n1303), .C2(new_n1305), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1293), .B1(new_n1301), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1306), .A2(new_n1258), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n847), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1306), .A2(G384), .A3(new_n1258), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1274), .A2(G2897), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1315), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT61), .B1(new_n1301), .B2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1274), .B1(new_n1294), .B2(new_n1299), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1321), .A2(KEYINPUT63), .A3(new_n1309), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1292), .A2(new_n1311), .A3(new_n1320), .A4(new_n1322), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1321), .A2(new_n1309), .A3(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT61), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1326), .B1(new_n1321), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT126), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(KEYINPUT62), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1330), .B1(new_n1321), .B2(new_n1309), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1325), .A2(new_n1328), .A3(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1323), .B1(new_n1332), .B2(new_n1292), .ZN(G405));
  INV_X1    g1133(.A(KEYINPUT127), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1334), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1290), .A2(new_n1287), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1338), .A2(KEYINPUT127), .A3(new_n1288), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(G375), .A2(new_n1270), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1310), .B1(new_n1340), .B2(new_n1294), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(new_n1310), .A3(new_n1294), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  OAI211_X1 g1143(.A(new_n1335), .B(new_n1339), .C1(new_n1341), .C2(new_n1343), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1343), .A2(new_n1341), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1345), .A2(KEYINPUT127), .A3(new_n1292), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(new_n1346), .ZN(G402));
endmodule


