//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  XOR2_X1   g001(.A(KEYINPUT71), .B(G218gat), .Z(new_n203));
  AOI21_X1  g002(.A(KEYINPUT22), .B1(new_n203), .B2(G211gat), .ZN(new_n204));
  XOR2_X1   g003(.A(G197gat), .B(G204gat), .Z(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT72), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g008(.A(KEYINPUT72), .B(new_n207), .C1(new_n204), .C2(new_n205), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n209), .A2(KEYINPUT73), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT73), .B1(new_n209), .B2(new_n210), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G148gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G141gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT76), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT75), .B(G141gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G148gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n215), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n214), .A2(G141gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n221), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT74), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n223), .B1(new_n220), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n229), .B1(new_n228), .B2(new_n220), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n219), .A2(new_n224), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT29), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n213), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n218), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT76), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n215), .B(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n224), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n230), .A2(new_n227), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n206), .A2(new_n207), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n206), .A2(new_n207), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n244), .A2(KEYINPUT29), .A3(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n242), .B1(new_n246), .B2(KEYINPUT3), .ZN(new_n247));
  NAND2_X1  g046(.A1(G228gat), .A2(G233gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n236), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT29), .B1(new_n209), .B2(new_n210), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n242), .B1(new_n251), .B2(KEYINPUT3), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n248), .B1(new_n236), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n202), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n253), .ZN(new_n255));
  INV_X1    g054(.A(new_n202), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n249), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G78gat), .B(G106gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(G22gat), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n254), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n259), .B1(new_n254), .B2(new_n257), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT35), .ZN(new_n263));
  INV_X1    g062(.A(new_n213), .ZN(new_n264));
  NAND2_X1  g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT26), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n268), .B1(new_n267), .B2(new_n266), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n269), .B1(G183gat), .B2(G190gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n271));
  AOI21_X1  g070(.A(G190gat), .B1(new_n271), .B2(KEYINPUT27), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT27), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(KEYINPUT27), .B(G183gat), .Z(new_n276));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n277), .A2(G190gat), .ZN(new_n278));
  OAI22_X1  g077(.A1(new_n275), .A2(KEYINPUT28), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n270), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT25), .ZN(new_n282));
  NAND3_X1  g081(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(G183gat), .B2(G190gat), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n285), .A2(KEYINPUT64), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(KEYINPUT64), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n284), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n266), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT23), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n266), .A2(KEYINPUT23), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n292), .A3(new_n265), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n282), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n284), .A2(new_n285), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n282), .B1(new_n289), .B2(new_n290), .ZN(new_n296));
  INV_X1    g095(.A(new_n265), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n297), .A2(KEYINPUT65), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n297), .A2(KEYINPUT65), .B1(new_n266), .B2(KEYINPUT23), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n295), .A2(new_n296), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT66), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n294), .A2(new_n303), .A3(new_n300), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n281), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(G226gat), .A2(G233gat), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(KEYINPUT29), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(new_n301), .B2(new_n280), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n264), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G8gat), .B(G36gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(G64gat), .B(G92gat), .ZN(new_n313));
  XOR2_X1   g112(.A(new_n312), .B(new_n313), .Z(new_n314));
  NAND3_X1  g113(.A1(new_n301), .A2(new_n280), .A3(new_n306), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n213), .B(new_n315), .C1(new_n305), .C2(new_n309), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n311), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n314), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n310), .B1(new_n305), .B2(new_n306), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(new_n213), .ZN(new_n320));
  INV_X1    g119(.A(new_n316), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n317), .A2(new_n322), .A3(KEYINPUT30), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n320), .A2(new_n321), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT30), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(new_n314), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n262), .A2(new_n263), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT78), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n330));
  INV_X1    g129(.A(G113gat), .ZN(new_n331));
  INV_X1    g130(.A(G120gat), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT1), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G113gat), .A2(G120gat), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n330), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G127gat), .B(G134gat), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n335), .B(new_n336), .Z(new_n337));
  OAI21_X1  g136(.A(new_n329), .B1(new_n242), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n335), .B(new_n336), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n231), .A2(KEYINPUT78), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n340), .A3(KEYINPUT4), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n242), .A2(new_n337), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT5), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n242), .A2(KEYINPUT3), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(new_n233), .A3(new_n337), .ZN(new_n348));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n345), .A2(new_n346), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT4), .B1(new_n338), .B2(new_n340), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n342), .A2(new_n343), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n348), .B(new_n349), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n242), .A2(new_n337), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n340), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n349), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n346), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n353), .B1(KEYINPUT79), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n357), .A2(KEYINPUT79), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n350), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT0), .ZN(new_n362));
  XNOR2_X1  g161(.A(G57gat), .B(G85gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n357), .A2(KEYINPUT79), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n357), .A2(KEYINPUT79), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(new_n368), .A3(new_n353), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n364), .A3(new_n350), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT6), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n366), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n360), .A2(KEYINPUT6), .A3(new_n365), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT84), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n328), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G15gat), .B(G43gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(G71gat), .B(G99gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n302), .A2(new_n304), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n280), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n339), .ZN(new_n382));
  INV_X1    g181(.A(G227gat), .ZN(new_n383));
  INV_X1    g182(.A(G233gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n305), .A2(new_n337), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT33), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n379), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(KEYINPUT32), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n387), .B(KEYINPUT32), .C1(new_n388), .C2(new_n379), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n385), .B1(new_n382), .B2(new_n386), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT34), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI211_X1 g195(.A(KEYINPUT34), .B(new_n385), .C1(new_n382), .C2(new_n386), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n396), .A2(new_n397), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT70), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n400), .A2(new_n391), .A3(new_n401), .A4(new_n392), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT70), .B1(new_n393), .B2(new_n398), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n327), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n406), .B1(new_n373), .B2(new_n372), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT69), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n393), .B1(new_n408), .B2(new_n400), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n398), .A2(KEYINPUT69), .A3(new_n391), .A4(new_n392), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n407), .A2(new_n411), .A3(new_n262), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n376), .A2(new_n405), .B1(new_n412), .B2(KEYINPUT35), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT37), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n311), .A2(KEYINPUT83), .A3(new_n414), .A4(new_n316), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n316), .B(new_n414), .C1(new_n319), .C2(new_n213), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT83), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n314), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n315), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n381), .B2(new_n308), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n414), .B1(new_n421), .B2(new_n264), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n213), .B1(new_n307), .B2(new_n310), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT38), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n419), .A2(new_n424), .B1(new_n314), .B2(new_n324), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n364), .B1(new_n369), .B2(new_n350), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT84), .B1(new_n426), .B2(KEYINPUT6), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n373), .A2(new_n374), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n372), .B(new_n425), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT85), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n375), .A2(new_n431), .A3(new_n372), .A4(new_n425), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n419), .B1(new_n414), .B2(new_n324), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT38), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n430), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n262), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n349), .B1(new_n345), .B2(new_n348), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT39), .B1(new_n355), .B2(new_n356), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT39), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n439), .A2(KEYINPUT40), .A3(new_n364), .A4(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT81), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n439), .A2(new_n364), .A3(new_n441), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT40), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n447), .A2(new_n366), .A3(new_n326), .A4(new_n323), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT82), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n442), .B(KEYINPUT81), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n426), .B1(new_n446), .B2(new_n445), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n406), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n436), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT36), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n404), .A2(new_n399), .A3(new_n455), .A4(new_n402), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT36), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n456), .B(new_n457), .C1(new_n407), .C2(new_n262), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n435), .A2(new_n454), .B1(KEYINPUT80), .B2(new_n458), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n456), .A2(new_n457), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT80), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n460), .B(new_n461), .C1(new_n407), .C2(new_n262), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n413), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G29gat), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT14), .B(G29gat), .ZN(new_n467));
  INV_X1    g266(.A(G36gat), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT86), .B(G43gat), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n472));
  INV_X1    g271(.A(G50gat), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT15), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OR2_X1    g275(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n478));
  AOI21_X1  g277(.A(G50gat), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G43gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G50gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT87), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n470), .B1(new_n476), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n473), .A2(G43gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(new_n481), .A3(KEYINPUT15), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n469), .A2(new_n486), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G22gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G15gat), .ZN(new_n492));
  INV_X1    g291(.A(G15gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G22gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT16), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT89), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n492), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G1gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n501), .B(new_n497), .C1(new_n495), .C2(G1gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n502), .A3(KEYINPUT91), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT90), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT90), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n500), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(G8gat), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT93), .ZN(new_n508));
  INV_X1    g307(.A(G8gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n503), .A2(KEYINPUT90), .A3(new_n509), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n508), .B1(new_n507), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n490), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n503), .A2(KEYINPUT90), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n506), .A2(G8gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n510), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT93), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n518));
  INV_X1    g317(.A(new_n490), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n513), .A2(KEYINPUT94), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n522), .B(KEYINPUT13), .Z(new_n523));
  INV_X1    g322(.A(KEYINPUT94), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n517), .A2(new_n524), .A3(new_n518), .A4(new_n519), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n521), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n521), .A2(KEYINPUT95), .A3(new_n523), .A4(new_n525), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G197gat), .ZN(new_n532));
  XOR2_X1   g331(.A(KEYINPUT11), .B(G169gat), .Z(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n534), .B(KEYINPUT12), .Z(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT15), .B1(new_n479), .B2(new_n472), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n471), .A2(new_n473), .ZN(new_n538));
  INV_X1    g337(.A(new_n482), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n469), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n486), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n489), .B(KEYINPUT88), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT17), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n487), .A2(KEYINPUT88), .A3(KEYINPUT17), .A4(new_n489), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT92), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n516), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n507), .A2(KEYINPUT92), .A3(new_n510), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(new_n522), .A3(new_n520), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT18), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n551), .A2(new_n520), .A3(KEYINPUT18), .A4(new_n522), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n530), .A2(new_n536), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT97), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n556), .B1(new_n528), .B2(new_n529), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n561), .A3(new_n536), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n530), .A2(new_n557), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(KEYINPUT96), .A3(new_n535), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(new_n560), .B2(new_n536), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n559), .A2(new_n562), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT98), .B1(new_n463), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n435), .A2(new_n454), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n458), .A2(KEYINPUT80), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n462), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n413), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT98), .ZN(new_n574));
  INV_X1    g373(.A(new_n567), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n568), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n517), .A2(new_n518), .ZN(new_n578));
  INV_X1    g377(.A(G57gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n579), .A2(KEYINPUT99), .ZN(new_n580));
  INV_X1    g379(.A(G64gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G71gat), .A2(G78gat), .ZN(new_n583));
  OR2_X1    g382(.A1(G71gat), .A2(G78gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT9), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n579), .A2(new_n581), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n583), .B(new_n584), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT21), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n596), .B1(new_n591), .B2(new_n595), .ZN(new_n599));
  OAI21_X1  g398(.A(G127gat), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n599), .ZN(new_n601));
  INV_X1    g400(.A(G127gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(new_n602), .A3(new_n597), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n594), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n600), .A2(new_n603), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(new_n578), .A3(new_n593), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G155gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n604), .A2(new_n606), .A3(new_n611), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT100), .ZN(new_n619));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G99gat), .B(G106gat), .Z(new_n623));
  NAND2_X1  g422(.A1(G85gat), .A2(G92gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT101), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT101), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(G85gat), .A3(G92gat), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n625), .A2(new_n627), .A3(KEYINPUT102), .A4(KEYINPUT7), .ZN(new_n628));
  NAND2_X1  g427(.A1(G99gat), .A2(G106gat), .ZN(new_n629));
  INV_X1    g428(.A(G85gat), .ZN(new_n630));
  INV_X1    g429(.A(G92gat), .ZN(new_n631));
  AOI22_X1  g430(.A1(KEYINPUT8), .A2(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(new_n624), .B2(KEYINPUT7), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT7), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(new_n624), .B2(KEYINPUT101), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n635), .B1(new_n627), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n623), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n627), .ZN(new_n640));
  INV_X1    g439(.A(new_n635), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n623), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n642), .A2(new_n643), .A3(new_n628), .A4(new_n632), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(new_n644), .A3(KEYINPUT103), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n633), .A2(new_n638), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(new_n647), .A3(new_n643), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n547), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(G190gat), .B(G218gat), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n519), .A2(new_n649), .B1(KEYINPUT41), .B2(new_n617), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n651), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n653), .B1(new_n651), .B2(new_n654), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n622), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n657), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(new_n621), .A3(new_n655), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n615), .A2(new_n661), .A3(KEYINPUT104), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT104), .B1(new_n615), .B2(new_n661), .ZN(new_n663));
  INV_X1    g462(.A(G230gat), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n384), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n645), .A2(new_n591), .A3(new_n648), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT105), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n645), .A2(new_n668), .A3(new_n648), .A4(new_n591), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT10), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n592), .A2(new_n644), .A3(new_n639), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n650), .A2(new_n671), .A3(new_n591), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n665), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  AOI211_X1 g476(.A(new_n664), .B(new_n384), .C1(new_n670), .C2(new_n673), .ZN(new_n678));
  XNOR2_X1  g477(.A(G120gat), .B(G148gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n679), .B(new_n680), .Z(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n677), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n682), .B1(new_n677), .B2(new_n678), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n662), .A2(new_n663), .A3(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n577), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n372), .A2(new_n373), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g491(.A1(new_n688), .A2(new_n406), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT16), .B(G8gat), .Z(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n509), .B1(new_n688), .B2(new_n406), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT42), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(new_n693), .B2(new_n695), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(G1325gat));
  INV_X1    g500(.A(new_n688), .ZN(new_n702));
  OAI21_X1  g501(.A(G15gat), .B1(new_n702), .B2(new_n460), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n493), .A3(new_n405), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(G1326gat));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n436), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT43), .B(G22gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  INV_X1    g508(.A(new_n661), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n458), .B1(new_n435), .B2(new_n454), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n709), .B(new_n710), .C1(new_n711), .C2(new_n413), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n661), .B1(new_n571), .B2(new_n572), .ZN(new_n713));
  OAI211_X1 g512(.A(KEYINPUT107), .B(new_n712), .C1(new_n713), .C2(new_n709), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n715), .B(KEYINPUT44), .C1(new_n463), .C2(new_n661), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n567), .A2(new_n615), .A3(new_n686), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(G29gat), .B1(new_n718), .B2(new_n689), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n686), .A2(new_n615), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n710), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n574), .B1(new_n573), .B2(new_n575), .ZN(new_n723));
  AOI211_X1 g522(.A(KEYINPUT98), .B(new_n567), .C1(new_n571), .C2(new_n572), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n690), .A2(new_n464), .ZN(new_n726));
  OR3_X1    g525(.A1(new_n725), .A2(KEYINPUT106), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT106), .B1(new_n725), .B2(new_n726), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n729), .B1(new_n727), .B2(new_n728), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n719), .B1(new_n730), .B2(new_n731), .ZN(G1328gat));
  AOI21_X1  g531(.A(new_n721), .B1(new_n568), .B2(new_n576), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(new_n468), .A3(new_n406), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n734), .A2(KEYINPUT46), .ZN(new_n735));
  OAI21_X1  g534(.A(G36gat), .B1(new_n718), .B2(new_n327), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(KEYINPUT46), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(G1329gat));
  OAI21_X1  g537(.A(new_n471), .B1(new_n718), .B2(new_n460), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n405), .A2(new_n477), .A3(new_n478), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n733), .A2(KEYINPUT108), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT108), .B1(new_n733), .B2(new_n740), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n739), .B(new_n744), .C1(new_n741), .C2(new_n742), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(G1330gat));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n262), .A2(G50gat), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(new_n733), .B2(KEYINPUT110), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n725), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n714), .A2(new_n436), .A3(new_n716), .A4(new_n717), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n752), .A2(new_n754), .B1(G50gat), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n749), .B1(new_n756), .B2(KEYINPUT48), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(G50gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n750), .B1(new_n725), .B2(new_n753), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n733), .A2(KEYINPUT110), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT48), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(KEYINPUT111), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n759), .B2(new_n760), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n752), .A2(KEYINPUT112), .A3(new_n754), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n762), .B1(new_n755), .B2(G50gat), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n757), .A2(new_n763), .A3(new_n768), .ZN(G1331gat));
  OR2_X1    g568(.A1(new_n711), .A2(new_n413), .ZN(new_n770));
  INV_X1    g569(.A(new_n686), .ZN(new_n771));
  NOR4_X1   g570(.A1(new_n575), .A2(new_n663), .A3(new_n662), .A4(new_n771), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n690), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n406), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n777));
  XOR2_X1   g576(.A(KEYINPUT49), .B(G64gat), .Z(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n776), .B2(new_n778), .ZN(G1333gat));
  INV_X1    g578(.A(G71gat), .ZN(new_n780));
  INV_X1    g579(.A(new_n460), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n773), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n405), .A2(new_n780), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n773), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g584(.A1(new_n773), .A2(new_n436), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g586(.A1(new_n575), .A2(new_n615), .A3(new_n771), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n714), .A2(new_n716), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n714), .A2(KEYINPUT113), .A3(new_n716), .A4(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G85gat), .B1(new_n793), .B2(new_n689), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n575), .A2(new_n615), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n770), .A2(new_n710), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT51), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n690), .A2(new_n630), .A3(new_n686), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT114), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n794), .B1(new_n797), .B2(new_n799), .ZN(G1336gat));
  NAND3_X1  g599(.A1(new_n406), .A2(new_n631), .A3(new_n686), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n801), .B(KEYINPUT115), .Z(new_n802));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n796), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n796), .A2(new_n803), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(new_n806), .B2(KEYINPUT116), .ZN(new_n807));
  OAI21_X1  g606(.A(G92gat), .B1(new_n789), .B2(new_n327), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n807), .B(new_n808), .C1(KEYINPUT116), .C2(new_n806), .ZN(new_n809));
  INV_X1    g608(.A(new_n806), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n791), .A2(new_n406), .A3(new_n792), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n811), .B2(G92gat), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n809), .B1(new_n812), .B2(new_n813), .ZN(G1337gat));
  OAI21_X1  g613(.A(G99gat), .B1(new_n793), .B2(new_n460), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n797), .A2(new_n771), .ZN(new_n816));
  INV_X1    g615(.A(G99gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n817), .A3(new_n405), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n818), .ZN(G1338gat));
  NOR2_X1   g618(.A1(new_n262), .A2(G106gat), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822));
  OAI21_X1  g621(.A(G106gat), .B1(new_n789), .B2(new_n262), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n820), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n797), .A2(new_n771), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n791), .A2(new_n436), .A3(new_n792), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n826), .B1(new_n827), .B2(G106gat), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n824), .B1(new_n828), .B2(new_n822), .ZN(G1339gat));
  AOI21_X1  g628(.A(new_n523), .B1(new_n521), .B2(new_n525), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n522), .B1(new_n551), .B2(new_n520), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n534), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT117), .ZN(new_n833));
  INV_X1    g632(.A(new_n562), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n561), .B1(new_n560), .B2(new_n536), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n686), .B(new_n833), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n681), .B1(new_n677), .B2(new_n837), .ZN(new_n838));
  AOI211_X1 g637(.A(KEYINPUT10), .B(new_n672), .C1(new_n667), .C2(new_n669), .ZN(new_n839));
  OAI22_X1  g638(.A1(new_n839), .A2(new_n675), .B1(new_n664), .B2(new_n384), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n674), .A2(new_n676), .A3(new_n665), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n841), .A3(KEYINPUT54), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n838), .A2(new_n842), .A3(KEYINPUT55), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT55), .B1(new_n838), .B2(new_n842), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n843), .A2(new_n844), .A3(new_n683), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n661), .B(new_n836), .C1(new_n567), .C2(new_n846), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n845), .B(new_n833), .C1(new_n834), .C2(new_n835), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n615), .B1(new_n848), .B2(new_n710), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n559), .A2(new_n562), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n564), .A2(new_n566), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n687), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n689), .A2(new_n406), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n855), .A2(new_n262), .A3(new_n405), .A4(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n857), .A2(new_n331), .A3(new_n567), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n853), .B1(new_n847), .B2(new_n849), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(new_n689), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n411), .A3(new_n262), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n406), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n575), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n858), .B1(new_n863), .B2(new_n331), .ZN(G1340gat));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n332), .A3(new_n686), .ZN(new_n865));
  OAI21_X1  g664(.A(G120gat), .B1(new_n857), .B2(new_n771), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g666(.A(new_n867), .B(KEYINPUT118), .Z(G1341gat));
  NAND3_X1  g667(.A1(new_n862), .A2(new_n602), .A3(new_n615), .ZN(new_n869));
  INV_X1    g668(.A(new_n615), .ZN(new_n870));
  OAI21_X1  g669(.A(G127gat), .B1(new_n857), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1342gat));
  NAND2_X1  g671(.A1(new_n327), .A2(new_n710), .ZN(new_n873));
  OR3_X1    g672(.A1(new_n861), .A2(G134gat), .A3(new_n873), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n857), .B2(new_n661), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G1343gat));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n460), .A2(new_n436), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT121), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n567), .A2(G141gat), .ZN(new_n882));
  AND4_X1   g681(.A1(new_n327), .A2(new_n860), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n879), .B1(new_n884), .B2(KEYINPUT120), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n460), .A2(new_n856), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n859), .A2(new_n887), .A3(new_n262), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n855), .A2(KEYINPUT57), .A3(new_n436), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n887), .B1(new_n859), .B2(new_n262), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(KEYINPUT119), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n890), .A2(new_n893), .A3(new_n575), .ZN(new_n894));
  INV_X1    g693(.A(new_n217), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n884), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT122), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n896), .A2(new_n899), .A3(new_n884), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n885), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n896), .B2(new_n884), .ZN(new_n902));
  AOI211_X1 g701(.A(KEYINPUT122), .B(new_n883), .C1(new_n894), .C2(new_n895), .ZN(new_n903));
  INV_X1    g702(.A(new_n885), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n901), .A2(new_n905), .ZN(G1344gat));
  NOR2_X1   g705(.A1(new_n214), .A2(KEYINPUT59), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n893), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n771), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n891), .A2(new_n892), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n886), .A2(new_n771), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n214), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n860), .A2(new_n881), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n915), .A2(new_n406), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n917), .A2(G148gat), .A3(new_n771), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n914), .A2(KEYINPUT123), .A3(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1345gat));
  OAI21_X1  g723(.A(G155gat), .B1(new_n908), .B2(new_n870), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n870), .A2(G155gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n917), .B2(new_n926), .ZN(G1346gat));
  OAI21_X1  g726(.A(G162gat), .B1(new_n908), .B2(new_n661), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n873), .A2(G162gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n915), .B2(new_n929), .ZN(G1347gat));
  NOR2_X1   g729(.A1(new_n690), .A2(new_n327), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n931), .A2(new_n411), .A3(new_n262), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n855), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(G169gat), .B1(new_n934), .B2(new_n575), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n855), .A2(new_n262), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n405), .A2(new_n931), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n575), .A2(G169gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(G1348gat));
  INV_X1    g739(.A(new_n938), .ZN(new_n941));
  OAI21_X1  g740(.A(G176gat), .B1(new_n941), .B2(new_n771), .ZN(new_n942));
  OR3_X1    g741(.A1(new_n933), .A2(G176gat), .A3(new_n771), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT124), .ZN(G1349gat));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n946), .A2(KEYINPUT60), .ZN(new_n947));
  OAI21_X1  g746(.A(G183gat), .B1(new_n941), .B2(new_n870), .ZN(new_n948));
  OR3_X1    g747(.A1(new_n933), .A2(new_n276), .A3(new_n870), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n946), .A2(KEYINPUT60), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n950), .B(new_n951), .Z(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n941), .B2(new_n661), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT61), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n661), .A2(G190gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n933), .B2(new_n955), .ZN(G1351gat));
  INV_X1    g755(.A(new_n931), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n781), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n959), .A2(new_n859), .A3(new_n262), .ZN(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n575), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n958), .B(KEYINPUT126), .Z(new_n962));
  AOI21_X1  g761(.A(new_n962), .B1(new_n891), .B2(new_n892), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n575), .A2(G197gat), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT127), .Z(G1352gat));
  INV_X1    g765(.A(new_n960), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n967), .A2(G204gat), .A3(new_n771), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT62), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n963), .A2(new_n686), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(G204gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n971), .ZN(G1353gat));
  INV_X1    g771(.A(G211gat), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n959), .A2(new_n870), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n973), .B1(new_n910), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT63), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n973), .A3(new_n615), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1354gat));
  AOI21_X1  g777(.A(G218gat), .B1(new_n960), .B2(new_n710), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n710), .A2(new_n203), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(new_n963), .B2(new_n980), .ZN(G1355gat));
endmodule


