//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n809, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929;
  INV_X1    g000(.A(G1gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT16), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT88), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G15gat), .B(G22gat), .Z(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(G8gat), .B1(new_n207), .B2(KEYINPUT89), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n202), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(new_n205), .B2(new_n206), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n208), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT21), .ZN(new_n212));
  XOR2_X1   g011(.A(G57gat), .B(G64gat), .Z(new_n213));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214));
  INV_X1    g013(.A(G71gat), .ZN(new_n215));
  INV_X1    g014(.A(G78gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G71gat), .B(G78gat), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n213), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n218), .B1(new_n213), .B2(new_n217), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT90), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n211), .B1(new_n212), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(G183gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n222), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n228), .ZN(new_n231));
  XNOR2_X1  g030(.A(G127gat), .B(G155gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(G211gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n224), .A2(new_n228), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n233), .B1(new_n236), .B2(new_n229), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT92), .ZN(new_n240));
  NAND2_X1  g039(.A1(G231gat), .A2(G233gat), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n240), .B(new_n241), .Z(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n235), .A2(new_n237), .A3(new_n242), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT100), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT17), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT15), .ZN(new_n249));
  XNOR2_X1  g048(.A(G43gat), .B(G50gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT86), .B(G29gat), .ZN(new_n252));
  INV_X1    g051(.A(G36gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT87), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT85), .ZN(new_n256));
  OAI22_X1  g055(.A1(new_n256), .A2(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(KEYINPUT14), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  AOI211_X1 g058(.A(new_n249), .B(new_n251), .C1(new_n255), .C2(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n251), .A2(new_n249), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n251), .A2(new_n249), .ZN(new_n263));
  AND4_X1   g062(.A1(new_n262), .A2(new_n255), .A3(new_n263), .A4(new_n259), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n248), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n255), .A2(new_n263), .A3(new_n259), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n261), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n255), .A2(new_n262), .A3(new_n263), .A4(new_n259), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(KEYINPUT17), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G85gat), .ZN(new_n270));
  INV_X1    g069(.A(G92gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT95), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT7), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n272), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G99gat), .ZN(new_n276));
  INV_X1    g075(.A(G106gat), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT96), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT96), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(G99gat), .A3(G106gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(KEYINPUT8), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT97), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n270), .A2(new_n271), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n281), .B2(new_n283), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n275), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(G99gat), .B(G106gat), .Z(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n287), .B(new_n275), .C1(new_n284), .C2(new_n285), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(KEYINPUT98), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT98), .B1(new_n289), .B2(new_n290), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n265), .B(new_n269), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G232gat), .A2(G233gat), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n295), .B(KEYINPUT93), .Z(new_n296));
  INV_X1    g095(.A(KEYINPUT41), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n289), .A2(new_n290), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT98), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n267), .A2(new_n268), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(new_n291), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n294), .A2(new_n298), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT99), .ZN(new_n305));
  XOR2_X1   g104(.A(G190gat), .B(G218gat), .Z(new_n306));
  INV_X1    g105(.A(KEYINPUT99), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n294), .A2(new_n303), .A3(new_n307), .A4(new_n298), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n306), .B1(new_n305), .B2(new_n308), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n247), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n311), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(KEYINPUT100), .A3(new_n309), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT94), .B(G134gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(G162gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n296), .A2(new_n297), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n316), .B(new_n317), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n312), .A2(new_n314), .A3(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n313), .A2(KEYINPUT100), .A3(new_n309), .A4(new_n318), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT35), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(G169gat), .B2(G176gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT24), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(G183gat), .A3(G190gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT24), .ZN(new_n331));
  NOR2_X1   g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n327), .B(new_n329), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n326), .A2(G169gat), .A3(G176gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n333), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT25), .B1(new_n333), .B2(KEYINPUT64), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n335), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT67), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT26), .ZN(new_n343));
  INV_X1    g142(.A(G169gat), .ZN(new_n344));
  INV_X1    g143(.A(G176gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT67), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n340), .A2(new_n347), .A3(new_n335), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n342), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT65), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT66), .B1(new_n350), .B2(KEYINPUT28), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT66), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT65), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT27), .ZN(new_n356));
  INV_X1    g155(.A(G183gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n359));
  AOI21_X1  g158(.A(G190gat), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n353), .A2(KEYINPUT65), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G190gat), .ZN(new_n363));
  AND2_X1   g162(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n361), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n351), .A4(new_n354), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n349), .A2(new_n362), .A3(new_n330), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n357), .A2(new_n363), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(KEYINPUT24), .A3(new_n330), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT64), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n371), .A2(new_n372), .A3(new_n327), .A4(new_n329), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n371), .A2(new_n327), .A3(new_n329), .A4(new_n335), .ZN(new_n374));
  OAI211_X1 g173(.A(KEYINPUT25), .B(new_n373), .C1(new_n374), .C2(new_n334), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n339), .A2(new_n369), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G120gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G113gat), .ZN(new_n378));
  INV_X1    g177(.A(G113gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(G120gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT1), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G134gat), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n384), .A2(KEYINPUT68), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(KEYINPUT68), .ZN(new_n386));
  OAI21_X1  g185(.A(G127gat), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT69), .B(G127gat), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n383), .B(new_n387), .C1(new_n384), .C2(new_n388), .ZN(new_n389));
  OR2_X1    g188(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n384), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(G134gat), .A3(new_n391), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n393), .A2(new_n382), .A3(new_n381), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n376), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n339), .A2(new_n369), .A3(new_n396), .A4(new_n375), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G227gat), .ZN(new_n401));
  INV_X1    g200(.A(G233gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n325), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n403), .ZN(new_n405));
  AOI211_X1 g204(.A(KEYINPUT71), .B(new_n405), .C1(new_n398), .C2(new_n399), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT32), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT33), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n408), .B1(new_n404), .B2(new_n406), .ZN(new_n409));
  XNOR2_X1  g208(.A(G15gat), .B(G43gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(G71gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(new_n276), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n407), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n412), .ZN(new_n414));
  OAI221_X1 g213(.A(KEYINPUT32), .B1(new_n408), .B2(new_n414), .C1(new_n404), .C2(new_n406), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n398), .A2(new_n405), .A3(new_n399), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT34), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n413), .A2(new_n418), .A3(new_n415), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(G211gat), .B(G218gat), .Z(new_n423));
  XOR2_X1   g222(.A(G197gat), .B(G204gat), .Z(new_n424));
  AOI21_X1  g223(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n425));
  OR3_X1    g224(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT73), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n428), .A2(new_n427), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT29), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT3), .ZN(new_n435));
  INV_X1    g234(.A(G141gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(G148gat), .ZN(new_n437));
  INV_X1    g236(.A(G148gat), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n438), .A2(G141gat), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT75), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(G155gat), .ZN(new_n441));
  INV_X1    g240(.A(G162gat), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT2), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n438), .A2(G141gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n436), .A2(G148gat), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT75), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G155gat), .B(G162gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT76), .B1(new_n436), .B2(G148gat), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT76), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n438), .A3(G141gat), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n454), .A3(new_n445), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(new_n449), .A3(new_n443), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT77), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n455), .A2(KEYINPUT77), .A3(new_n449), .A4(new_n443), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n434), .A2(new_n435), .B1(new_n451), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n451), .A2(new_n458), .A3(new_n435), .A4(new_n459), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n462), .A2(new_n433), .B1(new_n429), .B2(new_n430), .ZN(new_n463));
  OAI211_X1 g262(.A(G228gat), .B(G233gat), .C1(new_n461), .C2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n451), .A2(new_n458), .A3(new_n459), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT29), .B1(new_n426), .B2(new_n428), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n465), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n467));
  XOR2_X1   g266(.A(new_n467), .B(KEYINPUT79), .Z(new_n468));
  AOI21_X1  g267(.A(new_n463), .B1(G228gat), .B2(G233gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G78gat), .B(G106gat), .ZN(new_n471));
  INV_X1    g270(.A(G22gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  XOR2_X1   g272(.A(KEYINPUT31), .B(G50gat), .Z(new_n474));
  XOR2_X1   g273(.A(new_n473), .B(new_n474), .Z(new_n475));
  AND3_X1   g274(.A1(new_n464), .A2(new_n470), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n464), .B2(new_n470), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G8gat), .B(G36gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(G64gat), .B(G92gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n376), .A2(new_n433), .ZN(new_n483));
  NAND2_X1  g282(.A1(G226gat), .A2(G233gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n484), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n376), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n432), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n376), .A2(new_n486), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n486), .B1(new_n376), .B2(new_n433), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n431), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n488), .A2(new_n491), .A3(KEYINPUT74), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT74), .B1(new_n488), .B2(new_n491), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n482), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n489), .A2(new_n490), .A3(new_n431), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n432), .B1(new_n485), .B2(new_n487), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n482), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n494), .A2(KEYINPUT30), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT30), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n497), .A2(new_n501), .A3(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AND4_X1   g302(.A1(new_n324), .A2(new_n422), .A3(new_n479), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(new_n397), .A3(new_n462), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n460), .A2(KEYINPUT4), .A3(new_n451), .A4(new_n396), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n396), .A2(new_n451), .A3(new_n458), .A4(new_n459), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT4), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G225gat), .A2(G233gat), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n506), .A2(new_n507), .A3(new_n510), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n397), .A2(new_n465), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n508), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n512), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n514), .A2(KEYINPUT5), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n506), .A2(new_n507), .A3(new_n510), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G1gat), .B(G29gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G85gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT0), .B(G57gat), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n523), .B(new_n524), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n518), .A2(new_n525), .A3(new_n520), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT81), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI211_X1 g331(.A(new_n528), .B(new_n525), .C1(new_n518), .C2(new_n520), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT83), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n527), .A2(KEYINPUT81), .A3(new_n529), .A4(new_n528), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n525), .B1(new_n518), .B2(new_n520), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT6), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT83), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n532), .A2(new_n535), .A3(new_n536), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n504), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n530), .A2(new_n538), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n503), .A2(KEYINPUT78), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n419), .B1(new_n416), .B2(KEYINPUT72), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT72), .ZN(new_n545));
  AOI211_X1 g344(.A(new_n545), .B(new_n418), .C1(new_n413), .C2(new_n415), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n479), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT78), .B1(new_n503), .B2(new_n542), .ZN(new_n548));
  NOR3_X1   g347(.A1(new_n543), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n541), .B1(new_n549), .B2(new_n324), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT40), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT39), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n516), .A2(new_n512), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n506), .A2(new_n507), .A3(new_n510), .ZN(new_n554));
  AOI211_X1 g353(.A(new_n552), .B(new_n553), .C1(new_n512), .C2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n552), .A3(new_n512), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n525), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n551), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n500), .A2(new_n527), .A3(new_n502), .A4(new_n558), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n555), .A2(new_n557), .A3(new_n551), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n498), .B1(new_n497), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT38), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT37), .B1(new_n488), .B2(KEYINPUT82), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n488), .A2(new_n491), .A3(KEYINPUT82), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n562), .B(new_n563), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n488), .A2(new_n491), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n482), .B1(new_n567), .B2(KEYINPUT37), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT74), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n495), .B2(new_n496), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n488), .A2(new_n491), .A3(KEYINPUT74), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n568), .B1(new_n572), .B2(KEYINPUT37), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n566), .B(new_n499), .C1(new_n573), .C2(new_n563), .ZN(new_n574));
  OAI221_X1 g373(.A(new_n479), .B1(new_n559), .B2(new_n560), .C1(new_n540), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n478), .A2(KEYINPUT80), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT80), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n577), .B1(new_n476), .B2(new_n477), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(new_n543), .B2(new_n548), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT36), .B1(new_n544), .B2(new_n546), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n581), .B1(KEYINPUT36), .B2(new_n422), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n575), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  AOI211_X1 g382(.A(new_n246), .B(new_n323), .C1(new_n550), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT101), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n286), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n288), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n286), .A2(new_n587), .A3(new_n287), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n589), .A2(new_n221), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n222), .A2(new_n289), .A3(new_n290), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT10), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n301), .A2(KEYINPUT10), .A3(new_n225), .A4(new_n291), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n586), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n585), .B1(new_n591), .B2(new_n592), .ZN(new_n597));
  XNOR2_X1  g396(.A(G120gat), .B(G148gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n596), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n265), .A2(new_n211), .A3(new_n269), .ZN(new_n602));
  INV_X1    g401(.A(new_n211), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n302), .ZN(new_n604));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT18), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n211), .A2(new_n267), .A3(new_n268), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n605), .B(KEYINPUT13), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n602), .A2(KEYINPUT18), .A3(new_n604), .A4(new_n605), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n608), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G169gat), .B(G197gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G113gat), .B(G141gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n608), .A2(new_n621), .A3(new_n613), .A4(new_n614), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n601), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n600), .B1(new_n596), .B2(new_n597), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n584), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(new_n542), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n202), .ZN(G1324gat));
  NOR2_X1   g429(.A1(new_n628), .A2(new_n503), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT16), .B(G8gat), .Z(new_n632));
  OAI211_X1 g431(.A(new_n631), .B(new_n632), .C1(KEYINPUT102), .C2(KEYINPUT42), .ZN(new_n633));
  NAND2_X1  g432(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n631), .A2(KEYINPUT102), .A3(KEYINPUT42), .A4(new_n632), .ZN(new_n636));
  INV_X1    g435(.A(G8gat), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n631), .ZN(G1325gat));
  INV_X1    g437(.A(G15gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n422), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n628), .B2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT103), .Z(new_n642));
  NOR3_X1   g441(.A1(new_n628), .A2(new_n639), .A3(new_n582), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(G1326gat));
  INV_X1    g443(.A(new_n579), .ZN(new_n645));
  OAI21_X1  g444(.A(G22gat), .B1(new_n628), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n584), .A2(new_n472), .A3(new_n627), .A4(new_n579), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(G1327gat));
  AND3_X1   g449(.A1(new_n575), .A2(new_n580), .A3(new_n582), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT78), .ZN(new_n652));
  INV_X1    g451(.A(new_n502), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n501), .B1(new_n572), .B2(new_n482), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n653), .B1(new_n654), .B2(new_n499), .ZN(new_n655));
  INV_X1    g454(.A(new_n529), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n537), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n533), .B1(new_n657), .B2(new_n528), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n652), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n545), .B1(new_n413), .B2(new_n415), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(new_n419), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n503), .A2(KEYINPUT78), .A3(new_n542), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n659), .A2(new_n661), .A3(new_n479), .A4(new_n662), .ZN(new_n663));
  AOI22_X1  g462(.A1(new_n663), .A2(KEYINPUT35), .B1(new_n504), .B2(new_n540), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n323), .B1(new_n651), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n246), .A2(new_n627), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(new_n658), .A3(new_n252), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT45), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  OAI211_X1 g470(.A(KEYINPUT44), .B(new_n323), .C1(new_n651), .C2(new_n664), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n666), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n542), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n669), .B1(new_n676), .B2(new_n252), .ZN(G1328gat));
  NAND3_X1  g476(.A1(new_n667), .A2(new_n253), .A3(new_n655), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT46), .Z(new_n679));
  OAI21_X1  g478(.A(G36gat), .B1(new_n675), .B2(new_n503), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(G1329gat));
  INV_X1    g480(.A(new_n582), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n671), .A2(new_n682), .A3(new_n672), .A4(new_n674), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(G43gat), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n322), .B1(new_n550), .B2(new_n583), .ZN(new_n685));
  INV_X1    g484(.A(G43gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n686), .A3(new_n674), .ZN(new_n687));
  OR3_X1    g486(.A1(new_n687), .A2(KEYINPUT106), .A3(new_n640), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT106), .B1(new_n687), .B2(new_n640), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n684), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n690), .A2(KEYINPUT105), .A3(KEYINPUT47), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT47), .B1(new_n690), .B2(KEYINPUT105), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(G1330gat));
  OAI21_X1  g492(.A(G50gat), .B1(new_n675), .B2(new_n479), .ZN(new_n694));
  INV_X1    g493(.A(new_n667), .ZN(new_n695));
  AOI21_X1  g494(.A(G50gat), .B1(new_n695), .B2(KEYINPUT107), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n645), .B1(new_n667), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n694), .A2(new_n699), .A3(KEYINPUT48), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n673), .A2(new_n579), .A3(new_n674), .ZN(new_n701));
  AOI22_X1  g500(.A1(new_n701), .A2(G50gat), .B1(new_n696), .B2(new_n698), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(KEYINPUT48), .B2(new_n702), .ZN(G1331gat));
  INV_X1    g502(.A(new_n601), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n626), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n623), .A2(new_n624), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n584), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n658), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g511(.A(new_n503), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT108), .ZN(new_n714));
  OR3_X1    g513(.A1(new_n709), .A2(KEYINPUT109), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT109), .B1(new_n709), .B2(new_n714), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OR2_X1    g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1333gat));
  OAI21_X1  g518(.A(new_n215), .B1(new_n709), .B2(new_n640), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n682), .A2(G71gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n709), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g522(.A1(new_n709), .A2(new_n645), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(new_n216), .ZN(G1335gat));
  NAND2_X1  g524(.A1(new_n246), .A2(new_n708), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT110), .Z(new_n727));
  NAND2_X1  g526(.A1(new_n673), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G85gat), .B1(new_n728), .B2(new_n542), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n244), .A2(new_n245), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n707), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n323), .B(new_n731), .C1(new_n651), .C2(new_n664), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT51), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n685), .A2(KEYINPUT51), .A3(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n736), .A2(KEYINPUT111), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(KEYINPUT111), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n737), .A2(new_n270), .A3(new_n705), .A4(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n729), .B1(new_n739), .B2(new_n542), .ZN(G1336gat));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n671), .A2(new_n655), .A3(new_n672), .A4(new_n727), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G92gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n503), .A2(G92gat), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n732), .A2(new_n733), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT51), .B1(new_n685), .B2(new_n731), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n705), .B(new_n744), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n741), .B1(new_n748), .B2(KEYINPUT52), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750));
  AOI211_X1 g549(.A(KEYINPUT112), .B(new_n750), .C1(new_n743), .C2(new_n747), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n706), .B1(new_n734), .B2(new_n735), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n752), .A2(new_n744), .B1(new_n742), .B2(G92gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT114), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AND4_X1   g554(.A1(KEYINPUT114), .A2(new_n743), .A3(new_n747), .A4(new_n754), .ZN(new_n756));
  OAI22_X1  g555(.A1(new_n749), .A2(new_n751), .B1(new_n755), .B2(new_n756), .ZN(G1337gat));
  OAI21_X1  g556(.A(KEYINPUT115), .B1(new_n728), .B2(new_n582), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n673), .A2(new_n759), .A3(new_n682), .A4(new_n727), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(G99gat), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n422), .A2(new_n276), .A3(new_n705), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT116), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n737), .A2(new_n738), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(G1338gat));
  OAI21_X1  g564(.A(G106gat), .B1(new_n728), .B2(new_n479), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n277), .A3(new_n478), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n671), .A2(new_n579), .A3(new_n672), .A4(new_n727), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G106gat), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n767), .B2(new_n772), .ZN(G1339gat));
  NOR2_X1   g572(.A1(new_n610), .A2(new_n612), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n605), .B1(new_n602), .B2(new_n604), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n620), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n624), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n594), .A2(new_n595), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n585), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n594), .A2(new_n595), .A3(new_n586), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(KEYINPUT54), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n600), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n596), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n781), .A2(KEYINPUT55), .A3(new_n784), .ZN(new_n788));
  AND4_X1   g587(.A1(new_n704), .A2(new_n777), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n320), .A2(new_n789), .A3(new_n321), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n707), .A2(new_n787), .A3(new_n704), .A4(new_n788), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n777), .A2(new_n705), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n320), .A2(new_n321), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n246), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n707), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n322), .A2(new_n730), .A3(new_n795), .A4(new_n706), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n547), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n655), .A2(new_n542), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n799), .A2(new_n379), .A3(new_n707), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n579), .B1(new_n794), .B2(new_n796), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n801), .A2(new_n422), .A3(new_n798), .ZN(new_n802));
  OAI21_X1  g601(.A(G113gat), .B1(new_n802), .B2(new_n795), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT117), .Z(G1340gat));
  NAND3_X1  g604(.A1(new_n799), .A2(new_n377), .A3(new_n705), .ZN(new_n806));
  OAI21_X1  g605(.A(G120gat), .B1(new_n802), .B2(new_n706), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(G1341gat));
  AOI21_X1  g607(.A(new_n388), .B1(new_n799), .B2(new_n730), .ZN(new_n809));
  INV_X1    g608(.A(new_n388), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n802), .A2(new_n810), .A3(new_n246), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n809), .A2(new_n811), .ZN(G1342gat));
  OAI211_X1 g611(.A(new_n799), .B(new_n323), .C1(new_n385), .C2(new_n386), .ZN(new_n813));
  OR2_X1    g612(.A1(new_n813), .A2(KEYINPUT56), .ZN(new_n814));
  OAI21_X1  g613(.A(G134gat), .B1(new_n802), .B2(new_n322), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(KEYINPUT56), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(G1343gat));
  AOI21_X1  g616(.A(new_n479), .B1(new_n794), .B2(new_n796), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n582), .A2(new_n798), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n777), .A2(KEYINPUT118), .A3(new_n705), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT118), .B1(new_n777), .B2(new_n705), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT119), .B1(new_n781), .B2(new_n784), .ZN(new_n825));
  OAI221_X1 g624(.A(new_n625), .B1(new_n825), .B2(new_n786), .C1(KEYINPUT119), .C2(new_n787), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n824), .A2(new_n826), .B1(new_n321), .B2(new_n320), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n246), .B1(new_n827), .B2(new_n790), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n645), .B1(new_n828), .B2(new_n796), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n820), .B(new_n821), .C1(new_n819), .C2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(G141gat), .B1(new_n830), .B2(new_n795), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n818), .A2(new_n821), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(new_n436), .A3(new_n707), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT58), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n831), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(G1344gat));
  NAND3_X1  g637(.A1(new_n832), .A2(new_n438), .A3(new_n705), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n791), .A2(new_n792), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n322), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n320), .A2(new_n789), .A3(new_n321), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n730), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n796), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n478), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT57), .ZN(new_n847));
  INV_X1    g646(.A(new_n823), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n777), .A2(KEYINPUT118), .A3(new_n705), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n625), .B1(new_n786), .B2(new_n825), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n787), .A2(KEYINPUT119), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n848), .B(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n322), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n730), .B1(new_n853), .B2(new_n843), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n819), .B(new_n579), .C1(new_n854), .C2(new_n845), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n847), .A2(new_n855), .A3(new_n705), .A4(new_n821), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n438), .B1(new_n856), .B2(KEYINPUT120), .ZN(new_n857));
  AOI211_X1 g656(.A(KEYINPUT57), .B(new_n645), .C1(new_n828), .C2(new_n796), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n794), .A2(new_n796), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n819), .B1(new_n859), .B2(new_n478), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n861), .A2(new_n862), .A3(new_n705), .A4(new_n821), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n840), .B1(new_n857), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n840), .B(G148gat), .C1(new_n830), .C2(new_n706), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n839), .B1(new_n864), .B2(new_n866), .ZN(G1345gat));
  NAND2_X1  g666(.A1(new_n832), .A2(new_n730), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n441), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n730), .A2(G155gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n830), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n869), .B(KEYINPUT121), .C1(new_n830), .C2(new_n870), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1346gat));
  NOR3_X1   g674(.A1(new_n830), .A2(new_n442), .A3(new_n322), .ZN(new_n876));
  AOI21_X1  g675(.A(G162gat), .B1(new_n832), .B2(new_n323), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(G1347gat));
  NOR2_X1   g677(.A1(new_n658), .A2(new_n503), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n797), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n344), .A3(new_n707), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n801), .A2(new_n422), .A3(new_n879), .ZN(new_n882));
  OAI21_X1  g681(.A(G169gat), .B1(new_n882), .B2(new_n795), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1348gat));
  NAND3_X1  g683(.A1(new_n880), .A2(new_n345), .A3(new_n705), .ZN(new_n885));
  OAI21_X1  g684(.A(G176gat), .B1(new_n882), .B2(new_n706), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT122), .ZN(G1349gat));
  OAI211_X1 g687(.A(new_n880), .B(new_n730), .C1(new_n365), .C2(new_n364), .ZN(new_n889));
  OAI21_X1  g688(.A(G183gat), .B1(new_n882), .B2(new_n246), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g690(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n891), .B(new_n893), .ZN(G1350gat));
  NAND3_X1  g693(.A1(new_n880), .A2(new_n363), .A3(new_n323), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n882), .A2(new_n322), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n896), .A2(new_n897), .A3(G190gat), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n896), .B2(G190gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(G1351gat));
  XOR2_X1   g699(.A(KEYINPUT124), .B(G197gat), .Z(new_n901));
  NAND2_X1  g700(.A1(new_n582), .A2(new_n879), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n861), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n901), .B1(new_n904), .B2(new_n795), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n846), .A2(new_n902), .ZN(new_n906));
  INV_X1    g705(.A(new_n901), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n707), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n905), .A2(new_n908), .ZN(G1352gat));
  INV_X1    g708(.A(G204gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n906), .A2(new_n910), .A3(new_n705), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(KEYINPUT62), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(KEYINPUT62), .ZN(new_n913));
  NOR4_X1   g712(.A1(new_n858), .A2(new_n860), .A3(new_n706), .A4(new_n902), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n912), .B(new_n913), .C1(new_n910), .C2(new_n914), .ZN(G1353gat));
  NOR4_X1   g714(.A1(new_n846), .A2(G211gat), .A3(new_n246), .A4(new_n902), .ZN(new_n916));
  XOR2_X1   g715(.A(new_n916), .B(KEYINPUT125), .Z(new_n917));
  NAND4_X1  g716(.A1(new_n847), .A2(new_n855), .A3(new_n730), .A4(new_n903), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT63), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n918), .A2(new_n919), .A3(new_n920), .A4(G211gat), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n918), .A2(G211gat), .ZN(new_n922));
  NAND2_X1  g721(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n919), .A2(new_n920), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n917), .A2(new_n921), .A3(new_n925), .ZN(G1354gat));
  OAI21_X1  g725(.A(G218gat), .B1(new_n904), .B2(new_n322), .ZN(new_n927));
  INV_X1    g726(.A(G218gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n906), .A2(new_n928), .A3(new_n323), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1355gat));
endmodule


