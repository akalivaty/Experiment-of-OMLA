//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G116), .A2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n212), .B(new_n218), .C1(G107), .C2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT64), .B(G238), .Z(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G68), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n208), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(G13), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n208), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT0), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n231), .B(new_n236), .C1(new_n223), .C2(new_n224), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n226), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n215), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT2), .B(G226), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G58), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n256), .A2(new_n258), .A3(G226), .A4(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n256), .A2(new_n258), .A3(G223), .A4(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G87), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT76), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n259), .A2(new_n261), .A3(KEYINPUT76), .A4(new_n262), .ZN(new_n266));
  AND2_X1   g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n229), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G179), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n206), .A2(G274), .ZN(new_n271));
  OR2_X1    g0071(.A1(KEYINPUT66), .A2(G41), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT66), .A2(G41), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT67), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n206), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n268), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n277), .B1(new_n282), .B2(G232), .ZN(new_n283));
  AND3_X1   g0083(.A1(new_n269), .A2(new_n270), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(G169), .B1(new_n269), .B2(new_n283), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n287), .A2(new_n229), .ZN(new_n288));
  XNOR2_X1  g0088(.A(G58), .B(G68), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT74), .B1(new_n289), .B2(G20), .ZN(new_n290));
  AND2_X1   g0090(.A1(G58), .A2(G68), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G58), .A2(G68), .ZN(new_n292));
  OAI211_X1 g0092(.A(KEYINPUT74), .B(G20), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G159), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n207), .A2(new_n255), .A3(KEYINPUT68), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT68), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(G20), .B2(G33), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n290), .A2(new_n294), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G68), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT7), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT3), .B(G33), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(G20), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n256), .A2(new_n258), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n301), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT75), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT16), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(KEYINPUT7), .B1(new_n305), .B2(new_n207), .ZN(new_n311));
  AOI211_X1 g0111(.A(new_n302), .B(G20), .C1(new_n256), .C2(new_n258), .ZN(new_n312));
  OAI21_X1  g0112(.A(G68), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(G20), .B1(new_n291), .B2(new_n292), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT74), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n296), .A2(new_n298), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n316), .A2(new_n293), .B1(G159), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(KEYINPUT75), .A3(KEYINPUT16), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n288), .B1(new_n310), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT8), .B(G58), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n287), .A2(new_n229), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT70), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n206), .A2(G20), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT70), .B1(new_n324), .B2(new_n326), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n325), .B1(new_n332), .B2(new_n322), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n286), .B(KEYINPUT18), .C1(new_n321), .C2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT77), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n286), .B1(new_n321), .B2(new_n333), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT18), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(new_n335), .A3(new_n338), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT16), .B1(new_n319), .B2(KEYINPUT75), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT75), .ZN(new_n344));
  AOI211_X1 g0144(.A(new_n344), .B(new_n309), .C1(new_n313), .C2(new_n318), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n326), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n333), .ZN(new_n347));
  INV_X1    g0147(.A(G190), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n269), .A2(new_n283), .A3(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n206), .B(G274), .C1(new_n274), .C2(G45), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n280), .A2(new_n281), .ZN(new_n351));
  INV_X1    g0151(.A(new_n229), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G33), .A2(G41), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n350), .B1(new_n355), .B2(new_n215), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n354), .B1(new_n263), .B2(new_n264), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n356), .B1(new_n266), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n349), .B1(new_n358), .B2(G200), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n346), .A2(new_n347), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT17), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n346), .A2(new_n359), .A3(KEYINPUT17), .A4(new_n347), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n342), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n303), .A2(G1698), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(G223), .B1(G77), .B2(new_n305), .ZN(new_n368));
  INV_X1    g0168(.A(G222), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n303), .A2(new_n260), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n268), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n277), .B1(new_n282), .B2(G226), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n374), .A2(G169), .ZN(new_n375));
  INV_X1    g0175(.A(G50), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n324), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n322), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n255), .A2(G20), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n207), .B1(new_n292), .B2(new_n376), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n381), .A2(KEYINPUT69), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n317), .A2(G150), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(KEYINPUT69), .ZN(new_n384));
  AND4_X1   g0184(.A1(new_n380), .A2(new_n382), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n377), .B1(new_n332), .B2(new_n376), .C1(new_n385), .C2(new_n288), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n374), .A2(new_n270), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n375), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n386), .B(KEYINPUT9), .ZN(new_n389));
  INV_X1    g0189(.A(G200), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n372), .B2(new_n373), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(G190), .B2(new_n374), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT10), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n393), .B1(new_n389), .B2(new_n392), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n388), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n379), .A2(G77), .B1(G20), .B2(new_n301), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n299), .A2(KEYINPUT72), .A3(new_n376), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT72), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n317), .B2(G50), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n398), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT73), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n326), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n403), .B1(new_n402), .B2(new_n326), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT11), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n406), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT11), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(new_n404), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n327), .A2(G68), .A3(new_n330), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT12), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n324), .B2(new_n301), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n323), .A2(KEYINPUT12), .A3(G68), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n407), .A2(new_n410), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT14), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n215), .A2(G1698), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n303), .B(new_n419), .C1(G226), .C2(G1698), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G97), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n354), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n277), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT13), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n282), .A2(G238), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n423), .B2(new_n425), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n418), .B(G169), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n428), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n426), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n429), .B1(new_n270), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n418), .B1(new_n431), .B2(G169), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n417), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n407), .A2(new_n416), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n430), .A2(G190), .A3(new_n426), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(G200), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n435), .A2(new_n410), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G169), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT71), .B1(new_n370), .B2(new_n215), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT71), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n303), .A2(new_n441), .A3(G232), .A4(new_n260), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n366), .A2(new_n220), .B1(new_n203), .B2(new_n303), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n354), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n277), .B1(new_n282), .B2(G244), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n439), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n444), .B1(new_n442), .B2(new_n440), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n270), .B(new_n447), .C1(new_n450), .C2(new_n354), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT15), .B(G87), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n453), .A2(new_n379), .B1(G20), .B2(G77), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n299), .B2(new_n322), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n326), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n216), .B1(new_n206), .B2(G20), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n327), .A2(new_n457), .B1(new_n216), .B2(new_n324), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n449), .A2(new_n451), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n447), .B1(new_n450), .B2(new_n354), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n459), .B1(new_n461), .B2(G200), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(new_n348), .B2(new_n461), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n434), .A2(new_n438), .A3(new_n460), .A4(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n365), .A2(new_n397), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT5), .B1(new_n272), .B2(new_n273), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT5), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n206), .B(G45), .C1(new_n467), .C2(G41), .ZN(new_n468));
  OAI211_X1 g0268(.A(G270), .B(new_n354), .C1(new_n466), .C2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT85), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n273), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT66), .A2(G41), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n468), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n476), .A2(KEYINPUT85), .A3(G270), .A4(new_n354), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n466), .A2(new_n468), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT80), .ZN(new_n480));
  INV_X1    g0280(.A(G274), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n352), .B2(new_n353), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(G274), .B1(new_n267), .B2(new_n229), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT80), .B1(new_n476), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n256), .A2(new_n258), .A3(G264), .A4(G1698), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT86), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT86), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n303), .A2(new_n489), .A3(G264), .A4(G1698), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n305), .A2(G303), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n303), .A2(G257), .A3(new_n260), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n488), .A2(new_n490), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n268), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n478), .A2(new_n486), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G116), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n323), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n206), .A2(G33), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n288), .A2(new_n323), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n497), .B1(new_n500), .B2(new_n496), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n288), .B1(G20), .B2(new_n496), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G283), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n503), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT87), .ZN(new_n505));
  AOI21_X1  g0305(.A(G20), .B1(new_n255), .B2(G97), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT87), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(new_n507), .A3(new_n503), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n502), .A2(new_n509), .A3(KEYINPUT20), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT20), .B1(new_n502), .B2(new_n509), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n501), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n495), .A2(new_n512), .A3(G169), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT21), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT88), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n513), .A2(KEYINPUT88), .A3(new_n514), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n495), .A2(new_n512), .A3(KEYINPUT21), .A4(G169), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n483), .A2(new_n485), .B1(new_n493), .B2(new_n268), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n512), .A2(new_n521), .A3(G179), .A4(new_n478), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n512), .B1(new_n495), .B2(G200), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n348), .B2(new_n495), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n519), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n256), .A2(new_n258), .A3(G244), .A4(new_n260), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT4), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT78), .ZN(new_n531));
  OR2_X1    g0331(.A1(new_n528), .A2(new_n529), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT78), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n528), .A2(new_n533), .A3(new_n529), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n256), .A2(new_n258), .A3(G250), .A4(G1698), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n535), .A2(new_n503), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n531), .A2(new_n532), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n268), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n268), .B1(new_n474), .B2(new_n475), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n483), .A2(new_n485), .B1(G257), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G190), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT6), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n543), .A2(new_n202), .A3(G107), .ZN(new_n544));
  XNOR2_X1  g0344(.A(G97), .B(G107), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n546), .A2(new_n207), .B1(new_n216), .B2(new_n299), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n203), .B1(new_n304), .B2(new_n306), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n326), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n323), .A2(G97), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n500), .B2(G97), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n539), .A2(G257), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n480), .B1(new_n479), .B2(new_n482), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n476), .A2(KEYINPUT80), .A3(new_n484), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n538), .A2(KEYINPUT79), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT79), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n537), .A2(new_n558), .A3(new_n268), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n556), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n542), .B(new_n552), .C1(new_n560), .C2(new_n390), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n549), .A2(new_n551), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT81), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n549), .A2(KEYINPUT81), .A3(new_n551), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n537), .A2(new_n558), .A3(new_n268), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n558), .B1(new_n537), .B2(new_n268), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n270), .B(new_n540), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n538), .A2(new_n540), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n439), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n566), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n561), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n276), .A2(G1), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n268), .A2(new_n211), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT82), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n482), .A2(new_n576), .A3(new_n574), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n206), .A2(G45), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT82), .B1(new_n484), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n575), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n256), .A2(new_n258), .A3(G238), .A4(new_n260), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n256), .A2(new_n258), .A3(G244), .A4(G1698), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n581), .B(new_n582), .C1(new_n255), .C2(new_n496), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n268), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(new_n348), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT84), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n499), .B2(new_n210), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n327), .A2(KEYINPUT84), .A3(G87), .A4(new_n498), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n303), .A2(new_n207), .A3(G68), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n207), .B1(new_n421), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(G87), .B2(new_n204), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n596), .A2(KEYINPUT83), .A3(new_n592), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT83), .B1(new_n596), .B2(new_n592), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n326), .B1(new_n595), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n452), .A2(new_n324), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n590), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n390), .B1(new_n580), .B2(new_n584), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n586), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n580), .A2(new_n584), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n270), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n500), .A2(new_n453), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n600), .A2(new_n601), .A3(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n585), .A2(new_n439), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n604), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n303), .A2(new_n207), .A3(G87), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT22), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT22), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n303), .A2(new_n614), .A3(new_n207), .A4(G87), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT24), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT23), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(new_n203), .A3(G20), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT89), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n618), .B2(new_n203), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n622));
  OAI22_X1  g0422(.A1(new_n619), .A2(KEYINPUT89), .B1(new_n622), .B2(G20), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n616), .A2(new_n617), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n617), .B1(new_n616), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n326), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT25), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n323), .B2(G107), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n323), .A2(new_n628), .A3(G107), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n203), .A2(new_n499), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(G264), .B(new_n354), .C1(new_n466), .C2(new_n468), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n303), .A2(G257), .A3(G1698), .ZN(new_n636));
  NAND2_X1  g0436(.A1(G33), .A2(G294), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n636), .B(new_n637), .C1(new_n370), .C2(new_n211), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n268), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n486), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G169), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n485), .A2(new_n483), .B1(new_n638), .B2(new_n268), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n539), .A2(KEYINPUT90), .A3(G264), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT90), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n635), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n642), .A2(G179), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n634), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n640), .A2(G190), .ZN(new_n650));
  AOI21_X1  g0450(.A(G200), .B1(new_n642), .B2(new_n646), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n627), .B(new_n633), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n611), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n527), .A2(new_n573), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n465), .A2(new_n654), .ZN(G372));
  INV_X1    g0455(.A(new_n388), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n339), .A2(new_n334), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT92), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n460), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n449), .A2(KEYINPUT92), .A3(new_n451), .A4(new_n459), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n438), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n663), .A2(new_n434), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n362), .A2(new_n363), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n657), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n395), .A2(new_n396), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n656), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT91), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n610), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n585), .A2(KEYINPUT91), .A3(new_n439), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n609), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n602), .ZN(new_n675));
  INV_X1    g0475(.A(new_n603), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n675), .B(new_n676), .C1(new_n348), .C2(new_n585), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(new_n562), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n569), .A2(new_n571), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n669), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n569), .A2(new_n571), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n681), .A2(new_n611), .A3(KEYINPUT26), .A4(new_n566), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n561), .A2(new_n572), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n513), .A2(KEYINPUT88), .A3(new_n514), .ZN(new_n685));
  AOI21_X1  g0485(.A(KEYINPUT88), .B1(new_n513), .B2(new_n514), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n524), .B(new_n649), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n642), .A2(new_n646), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n688), .A2(G200), .B1(G190), .B2(new_n640), .ZN(new_n689));
  INV_X1    g0489(.A(new_n626), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n616), .A2(new_n617), .A3(new_n624), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n632), .B1(new_n692), .B2(new_n326), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n604), .B1(new_n689), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n684), .A2(new_n687), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n683), .A2(new_n695), .A3(new_n674), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n465), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n668), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT93), .ZN(G369));
  NAND3_X1  g0499(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  XOR2_X1   g0501(.A(new_n701), .B(KEYINPUT94), .Z(new_n702));
  OAI21_X1  g0502(.A(G213), .B1(new_n700), .B2(KEYINPUT27), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G343), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n512), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n527), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n524), .B1(new_n685), .B2(new_n686), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n708), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(G330), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n649), .A2(new_n652), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n693), .B2(new_n705), .ZN(new_n716));
  INV_X1    g0516(.A(new_n649), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n706), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n649), .A2(new_n706), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n706), .B1(new_n519), .B2(new_n524), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(new_n715), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n720), .A2(new_n723), .ZN(G399));
  NOR2_X1   g0524(.A1(new_n233), .A2(new_n274), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(G1), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n227), .B2(new_n726), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT95), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n646), .A2(new_n639), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n731), .B1(new_n732), .B2(new_n585), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n478), .A2(new_n486), .A3(new_n494), .A4(G179), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n605), .A2(KEYINPUT95), .A3(new_n639), .A4(new_n646), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n733), .A2(new_n541), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT30), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n570), .A2(new_n734), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n739), .A2(new_n740), .A3(new_n736), .A4(new_n733), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n642), .A2(new_n646), .ZN(new_n743));
  AOI21_X1  g0543(.A(G179), .B1(new_n580), .B2(new_n584), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(new_n495), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n560), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT96), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n742), .A2(KEYINPUT96), .A3(new_n747), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(new_n706), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT31), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n705), .A2(new_n753), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n654), .A2(new_n705), .B1(new_n748), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n696), .A2(new_n705), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT29), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n606), .A2(new_n608), .A3(new_n610), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n677), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n669), .B1(new_n572), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n604), .B1(new_n609), .B2(new_n673), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n681), .A2(new_n764), .A3(new_n562), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n763), .B1(new_n765), .B2(new_n669), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n695), .A2(new_n766), .A3(new_n674), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(KEYINPUT29), .A3(new_n705), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G330), .A2(new_n757), .B1(new_n760), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n730), .B1(new_n769), .B2(G1), .ZN(G364));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT97), .Z(new_n774));
  NOR3_X1   g0574(.A1(new_n709), .A2(new_n712), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n229), .B1(G20), .B2(new_n439), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n348), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n207), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n202), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n207), .A2(new_n270), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n348), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n207), .A2(G179), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(new_n348), .A3(G200), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n784), .A2(new_n376), .B1(new_n786), .B2(new_n203), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n782), .A2(G190), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n780), .B(new_n787), .C1(G68), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G190), .A2(G200), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G159), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT32), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n793), .A2(KEYINPUT32), .B1(new_n796), .B2(G87), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n781), .A2(new_n790), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n303), .B1(new_n798), .B2(new_n216), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n781), .A2(G190), .A3(new_n390), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n799), .B1(G58), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n789), .A2(new_n794), .A3(new_n797), .A4(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n801), .A2(G322), .B1(new_n792), .B2(G329), .ZN(new_n804));
  INV_X1    g0604(.A(new_n798), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n303), .B1(new_n805), .B2(G311), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n783), .A2(G326), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT33), .B(G317), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n788), .A2(new_n809), .B1(new_n796), .B2(G303), .ZN(new_n810));
  INV_X1    g0610(.A(new_n779), .ZN(new_n811));
  INV_X1    g0611(.A(new_n786), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n811), .A2(G294), .B1(new_n812), .B2(G283), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n807), .A2(new_n808), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n777), .B1(new_n803), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n232), .A2(G20), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n206), .B1(new_n816), .B2(G45), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n725), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n234), .A2(new_n303), .ZN(new_n820));
  INV_X1    g0620(.A(G355), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n820), .A2(new_n821), .B1(G116), .B2(new_n234), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n250), .A2(G45), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n233), .A2(new_n303), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n276), .B2(new_n228), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n822), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n773), .A2(new_n776), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n819), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  OR3_X1    g0630(.A1(new_n775), .A2(new_n815), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G330), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n711), .B(new_n832), .C1(new_n527), .C2(new_n708), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n833), .B(new_n713), .C1(new_n725), .C2(new_n818), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G396));
  NOR2_X1   g0636(.A1(new_n776), .A2(new_n771), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT98), .Z(new_n838));
  OAI21_X1  g0638(.A(new_n819), .B1(new_n838), .B2(G77), .ZN(new_n839));
  INV_X1    g0639(.A(G294), .ZN(new_n840));
  INV_X1    g0640(.A(G311), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n800), .A2(new_n840), .B1(new_n791), .B2(new_n841), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n303), .B(new_n842), .C1(G116), .C2(new_n805), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n796), .A2(G107), .ZN(new_n844));
  AOI22_X1  g0644(.A1(G283), .A2(new_n788), .B1(new_n783), .B2(G303), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n780), .B1(G87), .B2(new_n812), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n801), .A2(G143), .B1(new_n805), .B2(G159), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  INV_X1    g0649(.A(G150), .ZN(new_n850));
  INV_X1    g0650(.A(new_n788), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n848), .B1(new_n784), .B2(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT34), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(G132), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n303), .B1(new_n791), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(G68), .B2(new_n812), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n811), .A2(G58), .B1(new_n796), .B2(G50), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n854), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n852), .A2(new_n853), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n847), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n839), .B1(new_n861), .B2(new_n776), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n706), .A2(new_n459), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n661), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n463), .A2(new_n460), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n863), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT99), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n863), .B1(new_n659), .B2(new_n660), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n864), .B1(new_n463), .B2(new_n460), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT99), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n862), .B1(new_n873), .B2(new_n772), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT100), .Z(new_n875));
  NAND2_X1  g0675(.A1(new_n757), .A2(G330), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n706), .B1(new_n869), .B2(new_n872), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n696), .ZN(new_n878));
  INV_X1    g0678(.A(new_n674), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n694), .A2(new_n561), .A3(new_n572), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n879), .B1(new_n880), .B2(new_n687), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n706), .B1(new_n881), .B2(new_n683), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n878), .B1(new_n882), .B2(new_n873), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n876), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n819), .B1(new_n876), .B2(new_n883), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n875), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(G384));
  NOR2_X1   g0688(.A1(new_n816), .A2(new_n206), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n434), .A2(new_n706), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n704), .B1(new_n321), .B2(new_n333), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n337), .A2(new_n891), .A3(new_n360), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n337), .A2(new_n891), .A3(new_n360), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n665), .B1(new_n340), .B2(new_n341), .ZN(new_n897));
  OAI211_X1 g0697(.A(KEYINPUT38), .B(new_n896), .C1(new_n897), .C2(new_n891), .ZN(new_n898));
  XOR2_X1   g0698(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n899));
  NAND2_X1  g0699(.A1(new_n346), .A2(new_n347), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT18), .B1(new_n900), .B2(new_n286), .ZN(new_n901));
  INV_X1    g0701(.A(new_n334), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n362), .B(new_n363), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n891), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n896), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT103), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n903), .A2(new_n904), .B1(new_n893), .B2(new_n895), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT103), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n898), .B(new_n899), .C1(new_n908), .C2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n896), .B1(new_n897), .B2(new_n891), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n907), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n898), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT39), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n890), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n417), .A2(new_n706), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT102), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT102), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n417), .A2(new_n920), .A3(new_n706), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n919), .A2(new_n434), .A3(new_n438), .A4(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n417), .B(new_n706), .C1(new_n432), .C2(new_n433), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n460), .A2(new_n706), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n924), .B1(new_n878), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n915), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n657), .A2(new_n704), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n917), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT105), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n768), .B(new_n465), .C1(KEYINPUT29), .C2(new_n882), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n668), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT96), .B1(new_n742), .B2(new_n747), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n749), .B(new_n746), .C1(new_n738), .C2(new_n741), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n939), .A2(new_n755), .B1(new_n654), .B2(new_n705), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n754), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n922), .A2(new_n923), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n942), .A2(new_n873), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n910), .B1(new_n909), .B2(KEYINPUT38), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n893), .A2(new_n895), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n891), .B1(new_n364), .B2(new_n657), .ZN(new_n947));
  OAI211_X1 g0747(.A(KEYINPUT103), .B(new_n907), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n946), .B1(new_n365), .B2(new_n904), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n945), .A2(new_n948), .B1(new_n949), .B2(KEYINPUT38), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT40), .B1(new_n944), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT40), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n915), .A2(new_n941), .A3(new_n952), .A4(new_n943), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(new_n465), .A3(new_n941), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n941), .A2(new_n465), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n951), .A2(new_n956), .A3(new_n953), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n955), .A2(G330), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n889), .B1(new_n936), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n958), .B2(new_n936), .ZN(new_n960));
  INV_X1    g0760(.A(new_n546), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT35), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(KEYINPUT35), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n962), .A2(G116), .A3(new_n230), .A4(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT36), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n227), .A2(new_n291), .A3(new_n216), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT101), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n966), .A2(new_n967), .B1(new_n376), .B2(G68), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n967), .B2(new_n966), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(G1), .A3(new_n232), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n960), .A2(new_n965), .A3(new_n970), .ZN(G367));
  OAI221_X1 g0771(.A(new_n828), .B1(new_n234), .B2(new_n452), .C1(new_n245), .C2(new_n825), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(new_n819), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n706), .A2(new_n602), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n764), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n674), .B2(new_n974), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n851), .A2(new_n295), .B1(new_n795), .B2(new_n214), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G68), .B2(new_n811), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n800), .A2(new_n850), .B1(new_n791), .B2(new_n849), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n305), .B(new_n979), .C1(G50), .C2(new_n805), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n783), .A2(G143), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n812), .A2(G77), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n978), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n795), .A2(new_n496), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT46), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G107), .A2(new_n811), .B1(new_n783), .B2(G311), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n303), .B1(new_n801), .B2(G303), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G283), .A2(new_n805), .B1(new_n792), .B2(G317), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n788), .A2(G294), .B1(new_n812), .B2(G97), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n986), .A2(new_n987), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n983), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT47), .Z(new_n992));
  OAI221_X1 g0792(.A(new_n973), .B1(new_n976), .B2(new_n774), .C1(new_n777), .C2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n710), .A2(new_n715), .A3(new_n705), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n719), .B2(new_n722), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n714), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n713), .B(new_n994), .C1(new_n719), .C2(new_n722), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n760), .A2(new_n768), .ZN(new_n999));
  AND3_X1   g0799(.A1(new_n876), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT109), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n552), .A2(new_n705), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n681), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n573), .B2(new_n1003), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT108), .B1(new_n723), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n721), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n994), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n573), .A2(new_n1003), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1004), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT108), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1008), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1006), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT44), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n723), .A2(new_n1005), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1016), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1014), .A2(new_n1015), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1006), .A2(KEYINPUT44), .A3(new_n1013), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1001), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AND3_X1   g0822(.A1(new_n1008), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1012), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1015), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1025), .A2(new_n1021), .A3(new_n1001), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n720), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1000), .B1(new_n1022), .B2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1025), .A2(new_n720), .A3(new_n1021), .A4(new_n1026), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT110), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n769), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n725), .B(KEYINPUT41), .Z(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n818), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n720), .A2(new_n1011), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1011), .A2(new_n994), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT42), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n572), .B1(new_n1011), .B2(new_n649), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n705), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(KEYINPUT106), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT106), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1039), .A2(new_n1045), .A3(new_n1041), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n976), .B(KEYINPUT43), .Z(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1037), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1037), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1052), .B(new_n1047), .C1(new_n1053), .C2(new_n1049), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n993), .B1(new_n1036), .B2(new_n1055), .ZN(G387));
  NAND2_X1  g0856(.A1(new_n876), .A2(new_n999), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1057), .A2(KEYINPUT114), .A3(new_n996), .A4(new_n997), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT114), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n769), .B2(new_n998), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n726), .B1(new_n769), .B2(new_n998), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n719), .A2(new_n774), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n801), .A2(G317), .B1(new_n805), .B2(G303), .ZN(new_n1064));
  XOR2_X1   g0864(.A(KEYINPUT113), .B(G322), .Z(new_n1065));
  OAI221_X1 g0865(.A(new_n1064), .B1(new_n784), .B2(new_n1065), .C1(new_n841), .C2(new_n851), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT48), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n811), .A2(G283), .B1(new_n796), .B2(G294), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT49), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n786), .A2(new_n496), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n303), .B(new_n1075), .C1(G326), .C2(new_n792), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n798), .A2(new_n301), .B1(new_n791), .B2(new_n850), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n305), .B(new_n1078), .C1(G50), .C2(new_n801), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n795), .A2(new_n216), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n453), .A2(new_n811), .B1(new_n788), .B2(new_n378), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n783), .A2(G159), .B1(new_n812), .B2(G97), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n777), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n820), .A2(new_n727), .B1(G107), .B2(new_n234), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n242), .A2(new_n276), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n727), .B(new_n276), .C1(new_n301), .C2(new_n216), .ZN(new_n1088));
  XOR2_X1   g0888(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1089));
  NOR3_X1   g0889(.A1(new_n1089), .A2(G50), .A3(new_n322), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1089), .B1(G50), .B2(new_n322), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n825), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1086), .B1(new_n1087), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n819), .B1(new_n1094), .B2(new_n829), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT112), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1063), .A2(new_n1085), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n998), .B2(new_n818), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1062), .A2(new_n1098), .ZN(G393));
  NAND2_X1  g0899(.A1(new_n1011), .A2(new_n773), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n784), .A2(new_n850), .B1(new_n295), .B2(new_n800), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT51), .Z(new_n1102));
  AOI21_X1  g0902(.A(new_n305), .B1(new_n792), .B2(G143), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n322), .B2(new_n798), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n301), .A2(new_n795), .B1(new_n786), .B2(new_n210), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n851), .A2(new_n376), .B1(new_n216), .B2(new_n779), .ZN(new_n1106));
  OR4_X1    g0906(.A1(new_n1102), .A2(new_n1104), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G317), .A2(new_n783), .B1(new_n801), .B2(G311), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT116), .ZN(new_n1109));
  XOR2_X1   g0909(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1110));
  XNOR2_X1  g0910(.A(new_n1109), .B(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n788), .A2(G303), .B1(new_n812), .B2(G107), .ZN(new_n1112));
  INV_X1    g0912(.A(G283), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1112), .B1(new_n496), .B2(new_n779), .C1(new_n1113), .C2(new_n795), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n305), .B1(new_n798), .B2(new_n840), .C1(new_n791), .C2(new_n1065), .ZN(new_n1115));
  OR2_X1    g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1107), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n776), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n253), .A2(new_n824), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1119), .B(new_n828), .C1(new_n202), .C2(new_n234), .ZN(new_n1120));
  AND4_X1   g0920(.A1(new_n819), .A2(new_n1100), .A3(new_n1118), .A4(new_n1120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1020), .A2(KEYINPUT110), .A3(new_n720), .A4(new_n1021), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT110), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1031), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1122), .A2(new_n1124), .B1(new_n1125), .B2(new_n1028), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1121), .B1(new_n1126), .B2(new_n818), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n725), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1126), .A2(new_n1000), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(G390));
  AOI21_X1  g0930(.A(new_n925), .B1(new_n877), .B2(new_n696), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n890), .B1(new_n1131), .B2(new_n924), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n912), .A2(new_n916), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n898), .B1(new_n908), .B2(new_n911), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n767), .A2(new_n705), .A3(new_n873), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n926), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n942), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1134), .A2(new_n1137), .A3(new_n890), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n873), .A2(G330), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n924), .B(new_n1140), .C1(new_n940), .C2(new_n754), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT117), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT117), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n832), .B1(new_n869), .B2(new_n872), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT31), .B1(new_n939), .B2(new_n706), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n750), .A2(new_n751), .A3(new_n755), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n527), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n653), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1149), .A2(new_n684), .A3(new_n1150), .A4(new_n705), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1145), .B(new_n1146), .C1(new_n1147), .C2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1153), .A2(new_n757), .A3(new_n942), .A4(new_n1146), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1133), .A2(new_n1154), .A3(new_n1138), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1144), .A2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g0956(.A(G330), .B(new_n465), .C1(new_n1147), .C2(new_n1152), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT118), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT118), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n941), .A2(new_n1159), .A3(G330), .A4(new_n465), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n935), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n748), .A2(new_n755), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1151), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1147), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n924), .B1(new_n1164), .B2(new_n1140), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1140), .B1(new_n940), .B2(new_n754), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n942), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1131), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n942), .B(new_n1146), .C1(new_n1147), .C2(new_n1163), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1135), .A2(new_n926), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n942), .B1(new_n941), .B2(new_n1146), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1161), .B1(new_n1168), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1156), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1131), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n942), .B1(new_n757), .B2(new_n1146), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1176), .B1(new_n1141), .B2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1169), .B(new_n1170), .C1(new_n1166), .C2(new_n942), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1144), .A2(new_n1155), .A3(new_n1161), .A4(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1175), .A2(new_n1181), .A3(new_n725), .ZN(new_n1182));
  INV_X1    g0982(.A(G128), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n784), .A2(new_n1183), .B1(new_n786), .B2(new_n376), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n851), .A2(new_n849), .B1(new_n295), .B2(new_n779), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(G125), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n800), .A2(new_n855), .B1(new_n791), .B2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT54), .B(G143), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n305), .B(new_n1188), .C1(new_n805), .C2(new_n1190), .ZN(new_n1191));
  OR3_X1    g0991(.A1(new_n795), .A2(KEYINPUT53), .A3(new_n850), .ZN(new_n1192));
  OAI21_X1  g0992(.A(KEYINPUT53), .B1(new_n795), .B2(new_n850), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1186), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n779), .A2(new_n216), .B1(new_n800), .B2(new_n496), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT120), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n305), .B1(new_n798), .B2(new_n202), .C1(new_n210), .C2(new_n795), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n203), .A2(new_n851), .B1(new_n784), .B2(new_n1113), .ZN(new_n1198));
  OR3_X1    g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n786), .A2(new_n301), .B1(new_n791), .B2(new_n840), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT119), .Z(new_n1201));
  OAI21_X1  g1001(.A(new_n1194), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n777), .B1(new_n1202), .B2(KEYINPUT121), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(KEYINPUT121), .B2(new_n1202), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1204), .B(new_n819), .C1(new_n378), .C2(new_n838), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n950), .A2(new_n899), .B1(new_n915), .B2(KEYINPUT39), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1205), .B1(new_n1206), .B2(new_n771), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1156), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n1208), .B2(new_n818), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1182), .A2(new_n1209), .ZN(G378));
  AOI21_X1  g1010(.A(new_n832), .B1(new_n951), .B2(new_n953), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n386), .A2(new_n704), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n397), .A2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n397), .A2(new_n1214), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  OR3_X1    g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1218), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n912), .A2(new_n916), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n890), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n929), .B1(new_n927), .B2(new_n915), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1221), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1221), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n917), .A2(new_n931), .A3(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1212), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1227), .B1(new_n917), .B2(new_n931), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1225), .B(new_n1221), .C1(new_n1206), .C2(new_n890), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1211), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n818), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1227), .A2(new_n771), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n837), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n819), .B1(G50), .B2(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n274), .A2(new_n303), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n376), .B1(G33), .B2(G41), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G68), .A2(new_n811), .B1(new_n783), .B2(G116), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT122), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1238), .B1(new_n203), .B2(new_n800), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n798), .A2(new_n452), .B1(new_n791), .B2(new_n1113), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1081), .B1(new_n214), .B2(new_n786), .C1(new_n851), .C2(new_n202), .ZN(new_n1245));
  OR4_X1    g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT58), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1240), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  AOI211_X1 g1048(.A(G33), .B(G41), .C1(new_n792), .C2(G124), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n800), .A2(new_n1183), .B1(new_n795), .B2(new_n1189), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT123), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n784), .A2(new_n1187), .B1(new_n798), .B2(new_n849), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n851), .A2(new_n855), .B1(new_n850), .B2(new_n779), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT59), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1249), .B1(new_n295), .B2(new_n786), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1248), .B1(new_n1247), .B2(new_n1246), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1237), .B1(new_n1258), .B2(new_n776), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1235), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1234), .A2(new_n1260), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1133), .A2(new_n1138), .A3(new_n1154), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1142), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1174), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1161), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1230), .A2(new_n1211), .A3(new_n1231), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1211), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n1264), .A2(new_n1265), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT57), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n726), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1232), .A2(new_n1229), .B1(new_n1181), .B2(new_n1161), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(KEYINPUT57), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1261), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(G375));
  NOR2_X1   g1074(.A1(new_n1180), .A2(new_n1161), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1035), .A3(new_n1174), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n496), .A2(new_n851), .B1(new_n784), .B2(new_n840), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(G97), .B2(new_n796), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n811), .A2(new_n453), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n800), .A2(new_n1113), .B1(new_n798), .B2(new_n203), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n303), .B(new_n1281), .C1(G303), .C2(new_n792), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1279), .A2(new_n982), .A3(new_n1280), .A4(new_n1282), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n779), .A2(new_n376), .B1(new_n795), .B2(new_n295), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(G132), .B2(new_n783), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n305), .B1(new_n792), .B2(G128), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n801), .A2(G137), .B1(new_n805), .B2(G150), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n788), .A2(new_n1190), .B1(new_n812), .B2(G58), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n777), .B1(new_n1283), .B2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n819), .B1(new_n838), .B2(G68), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n1290), .B(new_n1291), .C1(new_n924), .C2(new_n771), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n1180), .B2(new_n818), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1277), .A2(new_n1293), .ZN(G381));
  NAND3_X1  g1094(.A1(new_n1277), .A2(new_n887), .A3(new_n1293), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1062), .A2(new_n835), .A3(new_n1098), .ZN(new_n1296));
  NOR4_X1   g1096(.A1(G378), .A2(G390), .A3(new_n1295), .A4(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(G387), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n1273), .ZN(G407));
  INV_X1    g1099(.A(G378), .ZN(new_n1300));
  INV_X1    g1100(.A(G213), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1301), .A2(G343), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1273), .A2(new_n1300), .A3(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(G407), .A2(new_n1303), .A3(G213), .ZN(G409));
  OAI211_X1 g1104(.A(new_n993), .B(G390), .C1(new_n1036), .C2(new_n1055), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(KEYINPUT126), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G393), .A2(G396), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT125), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1307), .A2(new_n1308), .A3(new_n1296), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1307), .B2(new_n1296), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1306), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(G390), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G387), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1305), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1312), .A2(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1306), .A2(new_n1314), .A3(new_n1311), .A4(new_n1305), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1275), .B1(KEYINPUT60), .B2(new_n1174), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1265), .A2(KEYINPUT60), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n725), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1293), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n887), .ZN(new_n1323));
  OAI211_X1 g1123(.A(G384), .B(new_n1293), .C1(new_n1319), .C2(new_n1321), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1302), .A2(G2897), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1323), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1325), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1271), .A2(new_n1035), .ZN(new_n1329));
  AOI22_X1  g1129(.A1(new_n1233), .A2(new_n818), .B1(new_n1235), .B2(new_n1259), .ZN(new_n1330));
  AOI21_X1  g1130(.A(G378), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1331), .B1(new_n1273), .B2(G378), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1328), .B1(new_n1332), .B2(new_n1302), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n725), .B1(new_n1271), .B2(KEYINPUT57), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1335));
  OAI211_X1 g1135(.A(G378), .B(new_n1330), .C1(new_n1334), .C2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1300), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1336), .A2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT62), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1302), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1339), .A2(new_n1340), .A3(new_n1341), .A4(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT61), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1333), .A2(new_n1344), .A3(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1302), .B1(new_n1336), .B2(new_n1338), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1340), .B1(new_n1347), .B2(new_n1343), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1318), .B1(new_n1346), .B2(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1316), .A2(new_n1345), .A3(new_n1317), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1339), .A2(new_n1341), .A3(new_n1343), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT63), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1350), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT124), .ZN(new_n1354));
  OAI211_X1 g1154(.A(new_n1328), .B(new_n1354), .C1(new_n1332), .C2(new_n1302), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1347), .A2(KEYINPUT63), .A3(new_n1343), .ZN(new_n1356));
  OR2_X1    g1156(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1357));
  OAI21_X1  g1157(.A(KEYINPUT124), .B1(new_n1357), .B2(new_n1347), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1353), .A2(new_n1355), .A3(new_n1356), .A4(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1349), .A2(new_n1359), .ZN(G405));
  NOR2_X1   g1160(.A1(new_n1273), .A2(G378), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1361), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1362), .A2(new_n1336), .A3(new_n1342), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1336), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1343), .B1(new_n1361), .B2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1363), .A2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT127), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1366), .A2(new_n1367), .A3(new_n1318), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1318), .A2(new_n1367), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1316), .A2(KEYINPUT127), .A3(new_n1317), .ZN(new_n1370));
  NAND4_X1  g1170(.A1(new_n1363), .A2(new_n1369), .A3(new_n1370), .A4(new_n1365), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1368), .A2(new_n1371), .ZN(G402));
endmodule


