//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n558, new_n559, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT67), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n461), .A2(new_n463), .A3(new_n466), .A4(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(new_n462), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(KEYINPUT3), .A3(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  AND3_X1   g049(.A1(new_n473), .A2(new_n474), .A3(new_n461), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n469), .A2(G2105), .B1(new_n475), .B2(G137), .ZN(new_n476));
  INV_X1    g051(.A(G101), .ZN(new_n477));
  AND2_X1   g052(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n474), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(KEYINPUT69), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(new_n474), .C1(new_n478), .C2(new_n479), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n477), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI211_X1 g061(.A(KEYINPUT70), .B(new_n477), .C1(new_n481), .C2(new_n483), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n476), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT71), .ZN(G160));
  AND3_X1   g064(.A1(new_n473), .A2(G2105), .A3(new_n461), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT72), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n494));
  XNOR2_X1  g069(.A(new_n494), .B(KEYINPUT73), .ZN(new_n495));
  INV_X1    g070(.A(G136), .ZN(new_n496));
  INV_X1    g071(.A(new_n475), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n492), .A2(new_n498), .ZN(G162));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n473), .A2(new_n461), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n461), .A2(new_n463), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n500), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n473), .A2(G126), .A3(G2105), .A4(new_n461), .ZN(new_n508));
  OR2_X1    g083(.A1(G102), .A2(G2105), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n509), .B(G2104), .C1(G114), .C2(new_n474), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  XOR2_X1   g089(.A(KEYINPUT5), .B(G543), .Z(new_n515));
  INV_X1    g090(.A(G62), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n517), .A2(G651), .B1(new_n520), .B2(G50), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT5), .B(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT74), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n518), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n521), .B1(new_n522), .B2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND3_X1  g105(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT75), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n520), .A2(G51), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n532), .B(new_n536), .C1(new_n537), .C2(new_n528), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  AND2_X1   g114(.A1(new_n525), .A2(new_n527), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT76), .B(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n515), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n545), .A2(G651), .B1(new_n520), .B2(G52), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  NAND2_X1  g123(.A1(new_n540), .A2(G81), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n515), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n552), .A2(G651), .B1(new_n520), .B2(G43), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n540), .A2(G91), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OR3_X1    g137(.A1(new_n519), .A2(KEYINPUT9), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n519), .B2(new_n562), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n523), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G651), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n561), .A2(new_n565), .A3(new_n568), .ZN(G299));
  NAND2_X1  g144(.A1(new_n540), .A2(G87), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n523), .A2(G74), .ZN(new_n571));
  AOI22_X1  g146(.A1(G49), .A2(new_n520), .B1(new_n571), .B2(G651), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n515), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G651), .ZN(new_n577));
  INV_X1    g152(.A(G48), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n519), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n525), .A2(G86), .A3(new_n527), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT77), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n525), .A2(new_n582), .A3(G86), .A4(new_n527), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  XOR2_X1   g160(.A(KEYINPUT78), .B(G47), .Z(new_n586));
  NAND2_X1  g161(.A1(new_n520), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  OAI221_X1 g164(.A(new_n587), .B1(new_n567), .B2(new_n588), .C1(new_n528), .C2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n540), .A2(G92), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n515), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(new_n520), .B2(G54), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n591), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n591), .B1(new_n600), .B2(G868), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G280));
  XOR2_X1   g181(.A(KEYINPUT79), .B(G559), .Z(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(G860), .B2(new_n607), .ZN(G148));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n554), .A2(new_n609), .ZN(new_n610));
  AND3_X1   g185(.A1(new_n594), .A2(new_n598), .A3(new_n607), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(new_n609), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n475), .A2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n490), .A2(G123), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n474), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT81), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n481), .A2(new_n483), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(new_n504), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT80), .B(G2100), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n623), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n620), .A2(new_n626), .ZN(G156));
  INV_X1    g202(.A(KEYINPUT14), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(new_n630), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n633), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(new_n641), .A3(G14), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT82), .Z(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT83), .Z(G401));
  INV_X1    g219(.A(KEYINPUT18), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT17), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n645), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2100), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n648), .B2(KEYINPUT18), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2096), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  AND2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT20), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n658), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n658), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n667), .B(new_n668), .Z(new_n669));
  XOR2_X1   g244(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT84), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G229));
  INV_X1    g250(.A(G29), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G33), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT25), .Z(new_n679));
  INV_X1    g254(.A(G139), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n497), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT91), .ZN(new_n682));
  AOI22_X1  g257(.A1(new_n504), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(new_n474), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n677), .B1(new_n685), .B2(new_n676), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n686), .A2(KEYINPUT92), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(KEYINPUT92), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G2072), .ZN(new_n690));
  NAND2_X1  g265(.A1(G162), .A2(G29), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G29), .B2(G35), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G2090), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n692), .A2(new_n694), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI22_X1  g273(.A1(new_n689), .A2(new_n690), .B1(new_n698), .B2(KEYINPUT98), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n555), .A2(G16), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G16), .B2(G19), .ZN(new_n701));
  INV_X1    g276(.A(G1341), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G5), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G171), .B2(new_n705), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n703), .B(new_n704), .C1(G1961), .C2(new_n707), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n490), .A2(G129), .B1(new_n475), .B2(G141), .ZN(new_n709));
  NAND3_X1  g284(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT26), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n621), .B2(G105), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(new_n676), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n676), .B2(G32), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT27), .B(G1996), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(G27), .A2(G29), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G164), .B2(G29), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n718), .B1(G2078), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(G2078), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n716), .B2(new_n717), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT99), .B(KEYINPUT23), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n705), .A2(G20), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G299), .B2(G16), .ZN(new_n727));
  INV_X1    g302(.A(G1956), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR4_X1   g304(.A1(new_n708), .A2(new_n721), .A3(new_n723), .A4(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n698), .A2(KEYINPUT98), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n705), .A2(G4), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n600), .B2(new_n705), .ZN(new_n733));
  INV_X1    g308(.A(G1348), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n699), .A2(new_n730), .A3(new_n731), .A4(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n687), .A2(G2072), .A3(new_n688), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT94), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT89), .B(KEYINPUT36), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n705), .A2(G23), .ZN(new_n742));
  INV_X1    g317(.A(G288), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(new_n705), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT33), .B(G1976), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT88), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT87), .B(KEYINPUT34), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n705), .A2(G22), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G166), .B2(new_n705), .ZN(new_n751));
  INV_X1    g326(.A(G1971), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n705), .A2(G6), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n584), .B2(new_n705), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT32), .B(G1981), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  AND3_X1   g333(.A1(new_n753), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n748), .A2(new_n749), .A3(new_n759), .ZN(new_n760));
  MUX2_X1   g335(.A(G24), .B(G290), .S(G16), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT86), .ZN(new_n762));
  INV_X1    g337(.A(G1986), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n676), .A2(G25), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n475), .A2(G131), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n490), .A2(G119), .ZN(new_n768));
  OR2_X1    g343(.A1(G95), .A2(G2105), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G2104), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n474), .A2(G107), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n767), .A2(new_n768), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n766), .B1(new_n774), .B2(new_n676), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT35), .B(G1991), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(KEYINPUT85), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n777), .A2(KEYINPUT85), .ZN(new_n779));
  NOR4_X1   g354(.A1(new_n764), .A2(new_n765), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n760), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n749), .B1(new_n748), .B2(new_n759), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n741), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n619), .A2(new_n676), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(KEYINPUT95), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(KEYINPUT95), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n705), .A2(G21), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G286), .B2(G16), .ZN(new_n788));
  INV_X1    g363(.A(G1966), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n791), .A2(G28), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n676), .B1(new_n791), .B2(G28), .ZN(new_n793));
  AND2_X1   g368(.A1(KEYINPUT31), .A2(G11), .ZN(new_n794));
  NOR2_X1   g369(.A1(KEYINPUT31), .A2(G11), .ZN(new_n795));
  OAI22_X1  g370(.A1(new_n792), .A2(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n707), .A2(G1961), .B1(new_n789), .B2(new_n788), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n785), .A2(new_n786), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT96), .ZN(new_n800));
  INV_X1    g375(.A(G34), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT24), .ZN(new_n802));
  AOI21_X1  g377(.A(G29), .B1(new_n801), .B2(KEYINPUT24), .ZN(new_n803));
  AOI22_X1  g378(.A1(G160), .A2(G29), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G2084), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT93), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n696), .B1(new_n695), .B2(new_n697), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n804), .A2(G2084), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n475), .A2(G140), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n490), .A2(G128), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n474), .A2(G116), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n809), .B(new_n810), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G29), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT90), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n676), .A2(G26), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT28), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G2067), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n807), .A2(new_n808), .A3(new_n819), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n800), .A2(new_n806), .A3(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n782), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n823), .A2(KEYINPUT89), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n822), .A2(new_n824), .A3(new_n760), .A4(new_n780), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n740), .A2(new_n783), .A3(new_n821), .A4(new_n825), .ZN(G150));
  INV_X1    g401(.A(KEYINPUT100), .ZN(new_n827));
  XNOR2_X1  g402(.A(G150), .B(new_n827), .ZN(G311));
  AOI22_X1  g403(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n829), .A2(new_n567), .B1(new_n830), .B2(new_n519), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n540), .B2(G93), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT101), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(new_n555), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT101), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n832), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(new_n554), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n600), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n842));
  AOI21_X1  g417(.A(G860), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n842), .B2(new_n841), .ZN(new_n844));
  INV_X1    g419(.A(new_n832), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n847), .ZN(G145));
  NAND2_X1  g423(.A1(new_n475), .A2(G142), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n490), .A2(G130), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n474), .A2(G118), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n623), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n774), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n813), .B(new_n512), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n685), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n857), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n682), .A2(new_n684), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n858), .A2(new_n714), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n714), .B1(new_n858), .B2(new_n861), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n856), .B(KEYINPUT104), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n864), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n866), .B(new_n862), .C1(new_n867), .C2(new_n855), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(G160), .B(KEYINPUT102), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(new_n619), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n619), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G162), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n871), .A2(G162), .A3(new_n872), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n869), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT105), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n869), .A2(new_n875), .A3(KEYINPUT105), .A4(new_n876), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n863), .A2(new_n864), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(KEYINPUT103), .A3(new_n856), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n866), .A2(KEYINPUT103), .A3(new_n862), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n855), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n883), .B(new_n885), .C1(KEYINPUT103), .C2(new_n882), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n875), .A2(new_n876), .ZN(new_n887));
  AOI21_X1  g462(.A(G37), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g465(.A(new_n584), .B(G290), .Z(new_n891));
  XNOR2_X1  g466(.A(G166), .B(G288), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(KEYINPUT42), .Z(new_n894));
  XNOR2_X1  g469(.A(new_n838), .B(new_n611), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n604), .B1(new_n594), .B2(new_n598), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n594), .A2(new_n604), .A3(new_n598), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  INV_X1    g476(.A(new_n898), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n901), .B1(new_n902), .B2(new_n896), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n897), .A2(KEYINPUT41), .A3(new_n898), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n900), .B1(new_n895), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n894), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  OAI21_X1  g486(.A(G868), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(G868), .B2(new_n832), .ZN(G295));
  OAI21_X1  g488(.A(new_n912), .B1(G868), .B2(new_n832), .ZN(G331));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n916));
  NAND2_X1  g491(.A1(G286), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(G286), .A2(new_n916), .ZN(new_n919));
  OAI21_X1  g494(.A(G171), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n919), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n921), .A2(new_n917), .A3(G301), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n838), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n920), .A2(new_n834), .A3(new_n837), .A4(new_n922), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n905), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n924), .A2(new_n897), .A3(new_n898), .A4(new_n925), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(G37), .B1(new_n929), .B2(new_n893), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n893), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n905), .A2(KEYINPUT108), .A3(new_n926), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n928), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n928), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT108), .B1(new_n905), .B2(new_n926), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n893), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  INV_X1    g516(.A(G37), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n940), .A2(new_n935), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n915), .B1(new_n937), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n935), .A2(new_n941), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n940), .A2(new_n942), .A3(new_n935), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n930), .A2(new_n945), .B1(new_n946), .B2(KEYINPUT43), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n944), .B1(new_n915), .B2(new_n947), .ZN(G397));
  OAI211_X1 g523(.A(new_n476), .B(G40), .C1(new_n486), .C2(new_n487), .ZN(new_n949));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n502), .A2(KEYINPUT4), .B1(new_n504), .B2(new_n505), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n508), .A2(new_n510), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G1996), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n957), .A3(new_n714), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT109), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n956), .B(KEYINPUT110), .Z(new_n960));
  INV_X1    g535(.A(G2067), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n813), .B(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n957), .B2(new_n714), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n959), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT111), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n774), .A2(new_n776), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n774), .A2(new_n776), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n960), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(G290), .B(G1986), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n956), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(G303), .A2(G8), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n973));
  OR3_X1    g548(.A1(new_n972), .A2(KEYINPUT113), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT113), .B1(new_n972), .B2(new_n973), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n973), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n949), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n980), .B(new_n950), .C1(new_n951), .C2(new_n952), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n953), .A2(KEYINPUT50), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n979), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT119), .ZN(new_n984));
  AOI21_X1  g559(.A(G2090), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n979), .A2(KEYINPUT119), .A3(new_n981), .A4(new_n982), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT45), .B1(new_n512), .B2(new_n950), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(new_n949), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT45), .B(new_n950), .C1(new_n951), .C2(new_n952), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n985), .A2(new_n986), .B1(new_n752), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G8), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n978), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n990), .A2(new_n994), .A3(new_n752), .ZN(new_n995));
  INV_X1    g570(.A(new_n989), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n987), .A2(new_n949), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT112), .B1(new_n997), .B2(G1971), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n484), .B(new_n485), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n982), .A2(new_n999), .A3(G40), .A4(new_n476), .ZN(new_n1000));
  INV_X1    g575(.A(new_n981), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n696), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n995), .A2(new_n998), .A3(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(G8), .A3(new_n977), .ZN(new_n1005));
  OAI21_X1  g580(.A(G8), .B1(new_n949), .B2(new_n953), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G87), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n572), .B(G1976), .C1(new_n1008), .C2(new_n528), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n570), .A2(KEYINPUT114), .A3(G1976), .A4(new_n572), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1976), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(G288), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1007), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT52), .B1(new_n1017), .B2(new_n1006), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n581), .A2(new_n583), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n576), .A2(G651), .B1(new_n520), .B2(G48), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT115), .B(G1981), .Z(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1981), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n1021), .B2(new_n580), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT49), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT116), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1026), .B1(new_n584), .B2(new_n1023), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n1032), .A3(KEYINPUT49), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1006), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1019), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n982), .ZN(new_n1037));
  NOR4_X1   g612(.A1(new_n1037), .A2(new_n949), .A3(new_n1001), .A4(G2084), .ZN(new_n1038));
  INV_X1    g613(.A(new_n488), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1039), .A2(KEYINPUT120), .A3(G40), .A4(new_n955), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n987), .B2(new_n949), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1040), .A2(new_n1042), .A3(new_n989), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1038), .B1(new_n1043), .B2(new_n789), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G168), .A2(G8), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n993), .A2(new_n1005), .A3(new_n1036), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT63), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT121), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT121), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1047), .A2(new_n1051), .A3(new_n1048), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n949), .A2(new_n953), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1054), .B(G8), .C1(new_n1031), .C2(KEYINPUT49), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1053), .B1(new_n1056), .B2(new_n1019), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1019), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1028), .A2(KEYINPUT116), .A3(new_n1029), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1032), .B1(new_n1031), .B2(KEYINPUT49), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1035), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1061), .A3(KEYINPUT117), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1057), .A2(new_n1062), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1044), .A2(new_n1048), .A3(new_n1045), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1004), .A2(G8), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n978), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1063), .A2(new_n1005), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1050), .A2(new_n1052), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1005), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1056), .A2(new_n1053), .A3(new_n1019), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT117), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1061), .A2(new_n1014), .A3(new_n743), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1006), .B1(new_n1074), .B2(new_n1024), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1069), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1005), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1078), .A2(KEYINPUT118), .A3(new_n1075), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n993), .A2(new_n1005), .A3(new_n1036), .ZN(new_n1081));
  INV_X1    g656(.A(G1961), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n983), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G2078), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT53), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT125), .B(new_n1083), .C1(new_n1043), .C2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n997), .A2(new_n1084), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1083), .B1(new_n1043), .B2(new_n1085), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(G301), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1087), .A2(new_n1088), .B1(new_n1082), .B2(new_n983), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n997), .A2(KEYINPUT53), .A3(new_n1084), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1095), .B1(new_n1098), .B2(G171), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1081), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(G301), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1089), .A2(G301), .A3(new_n1083), .A4(new_n1097), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT126), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT126), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1096), .A2(new_n1104), .A3(G301), .A4(new_n1097), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1095), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT51), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n992), .B1(new_n1044), .B2(G168), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n996), .B1(new_n988), .B2(KEYINPUT120), .ZN(new_n1110));
  AOI21_X1  g685(.A(G1966), .B1(new_n1110), .B2(new_n1042), .ZN(new_n1111));
  OAI21_X1  g686(.A(G286), .B1(new_n1111), .B2(new_n1038), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1108), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g688(.A(KEYINPUT51), .B(new_n992), .C1(new_n1044), .C2(G168), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT124), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1043), .A2(new_n789), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1038), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(G168), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(G8), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1044), .A2(G168), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT51), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1114), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1100), .A2(new_n1107), .A3(new_n1115), .A4(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n728), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT56), .B(G2072), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n979), .A2(new_n955), .A3(new_n989), .A4(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT122), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT57), .ZN(new_n1130));
  XNOR2_X1  g705(.A(G299), .B(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1126), .A2(KEYINPUT122), .A3(new_n1128), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n949), .A2(new_n953), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n983), .A2(new_n734), .B1(new_n961), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1126), .A2(new_n1131), .A3(new_n1128), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1138), .A2(new_n600), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1135), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n600), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1137), .A2(KEYINPUT60), .A3(new_n599), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1143), .A2(new_n1144), .B1(new_n1142), .B2(new_n1138), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1139), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1131), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NOR4_X1   g724(.A1(new_n987), .A2(new_n949), .A3(new_n996), .A4(G1996), .ZN(new_n1150));
  XOR2_X1   g725(.A(KEYINPUT58), .B(G1341), .Z(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1136), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n555), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT59), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1156), .B(new_n555), .C1(new_n1150), .C2(new_n1153), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1133), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1139), .A2(KEYINPUT61), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1149), .B(new_n1158), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1145), .B1(new_n1161), .B2(KEYINPUT123), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1135), .A2(KEYINPUT61), .A3(new_n1139), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n1149), .A4(new_n1158), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1141), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1068), .B(new_n1080), .C1(new_n1125), .C2(new_n1166), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1124), .A2(new_n1115), .A3(KEYINPUT62), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT62), .B1(new_n1124), .B2(new_n1115), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1101), .A2(new_n1005), .A3(new_n993), .A4(new_n1036), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n971), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n956), .A2(new_n957), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1173), .B(KEYINPUT46), .Z(new_n1174));
  NAND2_X1  g749(.A1(new_n962), .A2(new_n714), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1174), .B1(new_n960), .B2(new_n1175), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1176), .B(KEYINPUT47), .Z(new_n1177));
  NOR2_X1   g752(.A1(G290), .A2(G1986), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n956), .A2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT48), .Z(new_n1180));
  OAI21_X1  g755(.A(new_n1177), .B1(new_n969), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n965), .A2(new_n966), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(G2067), .B2(new_n813), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n960), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1172), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g760(.A1(G227), .A2(new_n458), .ZN(new_n1187));
  NOR2_X1   g761(.A1(new_n643), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g762(.A(new_n674), .B1(KEYINPUT127), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g763(.A(new_n1189), .B1(KEYINPUT127), .B2(new_n1188), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n1190), .A2(new_n889), .ZN(new_n1191));
  NOR2_X1   g765(.A1(new_n1191), .A2(new_n947), .ZN(G308));
  AND2_X1   g766(.A1(new_n945), .A2(new_n930), .ZN(new_n1193));
  AND2_X1   g767(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n1194));
  OAI211_X1 g768(.A(new_n889), .B(new_n1190), .C1(new_n1193), .C2(new_n1194), .ZN(G225));
endmodule


