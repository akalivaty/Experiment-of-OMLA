//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n462), .A2(G137), .B1(G101), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n460), .A2(KEYINPUT67), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n468), .A2(G125), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT68), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n468), .A2(new_n476), .A3(new_n473), .A4(G125), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n467), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n465), .B1(new_n478), .B2(new_n463), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n461), .A2(new_n463), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(G136), .B2(new_n462), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n490), .B(KEYINPUT69), .C1(new_n469), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  AOI21_X1  g068(.A(KEYINPUT69), .B1(new_n460), .B2(new_n490), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n488), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n490), .B1(new_n491), .B2(new_n469), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n498), .A2(KEYINPUT70), .A3(KEYINPUT4), .A4(new_n492), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n468), .A2(new_n473), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n489), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n495), .A2(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n504));
  OAI211_X1 g079(.A(G126), .B(G2105), .C1(new_n491), .C2(new_n469), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n502), .A2(new_n506), .ZN(G164));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  OR2_X1    g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(G651), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n518), .A2(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n522), .A2(G543), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n522), .A2(new_n511), .A3(new_n523), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n516), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT72), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n527), .A2(KEYINPUT72), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n515), .B1(new_n529), .B2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  INV_X1    g107(.A(new_n525), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G89), .ZN(new_n534));
  INV_X1    g109(.A(new_n524), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT73), .B(G51), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n540));
  AND2_X1   g115(.A1(G63), .A2(G651), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n539), .A2(new_n540), .B1(new_n511), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n534), .A2(new_n537), .A3(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND2_X1  g119(.A1(new_n533), .A2(G90), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n520), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n535), .A2(G52), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  XNOR2_X1  g125(.A(KEYINPUT74), .B(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n535), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n520), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n533), .A2(G81), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  AOI22_X1  g137(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n520), .B1(new_n563), .B2(new_n564), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n565), .A2(new_n566), .B1(new_n533), .B2(G91), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n522), .A2(G53), .A3(G543), .A4(new_n523), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT9), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(G299));
  NAND2_X1  g145(.A1(new_n535), .A2(G49), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n533), .A2(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  AOI22_X1  g149(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(new_n520), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n535), .A2(G48), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n533), .A2(G86), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G305));
  XOR2_X1   g154(.A(KEYINPUT76), .B(G85), .Z(new_n580));
  NAND2_X1  g155(.A1(new_n533), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(new_n520), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n535), .A2(G47), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(G290));
  INV_X1    g160(.A(G868), .ZN(new_n586));
  NOR2_X1   g161(.A1(G301), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n522), .A2(G92), .A3(new_n511), .A4(new_n523), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n588), .A2(KEYINPUT77), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(KEYINPUT77), .ZN(new_n590));
  AOI21_X1  g165(.A(KEYINPUT10), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G54), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n520), .A2(new_n592), .B1(new_n524), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n589), .A2(KEYINPUT10), .A3(new_n590), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT78), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n587), .B1(new_n598), .B2(new_n586), .ZN(G284));
  AOI21_X1  g174(.A(new_n587), .B1(new_n598), .B2(new_n586), .ZN(G321));
  NAND2_X1  g175(.A1(G299), .A2(new_n586), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n586), .B2(G168), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(new_n586), .B2(G168), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n598), .B1(new_n604), .B2(G860), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT79), .Z(G148));
  NOR2_X1   g181(.A1(new_n557), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n604), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT80), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n500), .A2(new_n464), .ZN(new_n612));
  XOR2_X1   g187(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G2100), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT82), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n462), .A2(G135), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n483), .A2(G123), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n463), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(G2096), .Z(new_n623));
  OAI211_X1 g198(.A(new_n617), .B(new_n623), .C1(G2100), .C2(new_n615), .ZN(G156));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT83), .B(G2438), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n625), .B(new_n626), .Z(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2430), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n631), .B(new_n635), .Z(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  AND3_X1   g214(.A1(new_n638), .A2(G14), .A3(new_n639), .ZN(G401));
  INV_X1    g215(.A(KEYINPUT18), .ZN(new_n641));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT17), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2100), .ZN(new_n648));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n644), .B2(KEYINPUT18), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2096), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(G227));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT85), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1961), .B(G1966), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT20), .Z(new_n662));
  NAND2_X1  g237(.A1(new_n655), .A2(new_n656), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n657), .A2(new_n663), .A3(new_n660), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n662), .B(new_n664), .C1(new_n660), .C2(new_n663), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1991), .B(G1996), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G229));
  NOR2_X1   g246(.A1(G6), .A2(G16), .ZN(new_n672));
  AND3_X1   g247(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n672), .B1(new_n673), .B2(G16), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT32), .ZN(new_n675));
  INV_X1    g250(.A(G1981), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G23), .ZN(new_n679));
  INV_X1    g254(.A(G288), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n678), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT33), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(G166), .A2(G16), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G16), .B2(G22), .ZN(new_n685));
  INV_X1    g260(.A(G1971), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n677), .B(new_n687), .C1(new_n686), .C2(new_n685), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G25), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n462), .A2(G131), .ZN(new_n693));
  INV_X1    g268(.A(G119), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n694), .B2(new_n484), .ZN(new_n695));
  OAI21_X1  g270(.A(KEYINPUT86), .B1(G95), .B2(G2105), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g272(.A1(KEYINPUT86), .A2(G95), .A3(G2105), .ZN(new_n698));
  OAI221_X1 g273(.A(G2104), .B1(G107), .B2(new_n463), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n692), .B1(new_n701), .B2(new_n691), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT35), .B(G1991), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G24), .ZN(new_n705));
  XOR2_X1   g280(.A(G290), .B(KEYINPUT87), .Z(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G16), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(G1986), .Z(new_n708));
  NAND4_X1  g283(.A1(new_n689), .A2(new_n690), .A3(new_n704), .A4(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT36), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n678), .A2(G4), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n598), .B2(new_n678), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT88), .Z(new_n713));
  INV_X1    g288(.A(G1348), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G29), .A2(G35), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G162), .B2(G29), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G2090), .ZN(new_n722));
  NOR2_X1   g297(.A1(G171), .A2(new_n678), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G5), .B2(new_n678), .ZN(new_n724));
  INV_X1    g299(.A(G1961), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n721), .A2(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(G168), .A2(new_n678), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n678), .B2(G21), .ZN(new_n728));
  INV_X1    g303(.A(G1966), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n726), .B(new_n730), .C1(new_n722), .C2(new_n721), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n678), .A2(G19), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n557), .B2(new_n678), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1341), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT30), .B(G28), .ZN(new_n735));
  OR2_X1    g310(.A1(KEYINPUT31), .A2(G11), .ZN(new_n736));
  NAND2_X1  g311(.A1(KEYINPUT31), .A2(G11), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n735), .A2(new_n691), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n622), .B2(new_n691), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n691), .A2(G32), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n462), .A2(G141), .B1(G105), .B2(new_n464), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n483), .A2(G129), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT26), .Z(new_n744));
  NAND3_X1  g319(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n740), .B1(new_n745), .B2(G29), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT27), .B(G1996), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n739), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n748), .B1(new_n746), .B2(new_n747), .C1(new_n724), .C2(new_n725), .ZN(new_n749));
  OR3_X1    g324(.A1(new_n731), .A2(new_n734), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n728), .A2(new_n729), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(KEYINPUT94), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(KEYINPUT94), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n691), .A2(G26), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT28), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n462), .A2(G140), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n483), .A2(G128), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n463), .A2(G116), .ZN(new_n758));
  OAI21_X1  g333(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n756), .B(new_n757), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n755), .B1(new_n762), .B2(G29), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2067), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n752), .A2(new_n753), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n500), .A2(G127), .ZN(new_n766));
  NAND2_X1  g341(.A1(G115), .A2(G2104), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n463), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT90), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT25), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n462), .B2(G139), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n770), .A2(new_n771), .A3(new_n774), .ZN(new_n775));
  MUX2_X1   g350(.A(G33), .B(new_n775), .S(G29), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2072), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n678), .A2(G20), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT23), .Z(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G299), .B2(G16), .ZN(new_n780));
  INV_X1    g355(.A(G1956), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G2084), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(G34), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(G29), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n786), .A2(KEYINPUT92), .B1(G34), .B2(new_n784), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(KEYINPUT92), .B2(new_n786), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n479), .B2(new_n691), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n782), .B1(new_n783), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(new_n783), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT93), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n691), .A2(G27), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G164), .B2(new_n691), .ZN(new_n794));
  INV_X1    g369(.A(G2078), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n790), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NOR4_X1   g372(.A1(new_n750), .A2(new_n765), .A3(new_n777), .A4(new_n797), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n717), .A2(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(KEYINPUT96), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n717), .A2(KEYINPUT96), .A3(new_n798), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n710), .B1(new_n800), .B2(new_n801), .ZN(G311));
  INV_X1    g377(.A(new_n710), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n799), .A2(KEYINPUT96), .ZN(new_n804));
  INV_X1    g379(.A(new_n801), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(G150));
  NAND2_X1  g381(.A1(new_n598), .A2(G559), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n533), .A2(G93), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(new_n520), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n535), .A2(G55), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n810), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT98), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT98), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n810), .A2(new_n812), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n815), .A2(new_n557), .A3(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n557), .B1(new_n815), .B2(new_n817), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n809), .B(new_n821), .Z(new_n822));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n823));
  AOI21_X1  g398(.A(G860), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n823), .B2(new_n822), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n814), .A2(G860), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT99), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT37), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n828), .ZN(G145));
  NOR2_X1   g404(.A1(new_n775), .A2(KEYINPUT101), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n506), .A2(KEYINPUT100), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT100), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n504), .A2(new_n505), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n495), .A2(new_n499), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n500), .A2(new_n501), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n762), .B(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n830), .B1(new_n838), .B2(new_n745), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n745), .B2(new_n838), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n775), .A2(KEYINPUT101), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n483), .A2(G130), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT102), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n462), .A2(G142), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(KEYINPUT103), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(KEYINPUT103), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(G118), .B2(new_n463), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n844), .B(new_n845), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(new_n701), .Z(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(new_n614), .Z(new_n852));
  OR2_X1    g427(.A1(new_n842), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n842), .A2(new_n852), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n479), .B(new_n622), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(G162), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G37), .ZN(new_n859));
  INV_X1    g434(.A(new_n857), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n853), .A2(new_n860), .A3(new_n854), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g438(.A1(new_n814), .A2(new_n586), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n608), .B(new_n821), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n597), .A2(new_n866), .A3(G299), .ZN(new_n867));
  NAND2_X1  g442(.A1(G299), .A2(new_n866), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n567), .A2(new_n569), .A3(KEYINPUT104), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n868), .A2(new_n595), .A3(new_n596), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n867), .A2(new_n870), .A3(KEYINPUT41), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n865), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n871), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n865), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G290), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n879), .A2(new_n680), .ZN(new_n880));
  NOR2_X1   g455(.A1(G290), .A2(G288), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n673), .B(new_n515), .C1(new_n529), .C2(new_n530), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT105), .B1(new_n880), .B2(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(G303), .A2(G305), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n884), .A2(new_n885), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  INV_X1    g464(.A(new_n885), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n883), .B(new_n882), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT42), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n878), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n864), .B1(new_n894), .B2(new_n586), .ZN(G295));
  OAI21_X1  g470(.A(new_n864), .B1(new_n894), .B2(new_n586), .ZN(G331));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n897));
  INV_X1    g472(.A(new_n892), .ZN(new_n898));
  XNOR2_X1  g473(.A(G301), .B(G286), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n820), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n901), .A3(new_n818), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n899), .B1(new_n819), .B2(new_n820), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n873), .A2(new_n904), .A3(new_n874), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(KEYINPUT106), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n907), .B(new_n899), .C1(new_n819), .C2(new_n820), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n877), .A2(new_n906), .A3(new_n902), .A4(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n898), .A2(new_n905), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n859), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n898), .B1(new_n905), .B2(new_n909), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n897), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n906), .A2(new_n902), .A3(new_n908), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(new_n874), .A3(new_n873), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n877), .A2(new_n903), .A3(new_n902), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n898), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n920), .A2(new_n859), .A3(new_n910), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT108), .B1(new_n921), .B2(KEYINPUT43), .ZN(new_n922));
  OAI211_X1 g497(.A(KEYINPUT108), .B(KEYINPUT43), .C1(new_n911), .C2(new_n919), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n915), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n920), .A2(new_n914), .A3(new_n859), .A4(new_n910), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n911), .B2(new_n912), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT107), .B1(new_n928), .B2(new_n897), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n930));
  AOI211_X1 g505(.A(new_n930), .B(KEYINPUT44), .C1(new_n926), .C2(new_n927), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n925), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n925), .B(KEYINPUT109), .C1(new_n929), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(G397));
  INV_X1    g511(.A(KEYINPUT126), .ZN(new_n937));
  INV_X1    g512(.A(G2067), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n762), .B(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G1996), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n745), .B(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n701), .A2(new_n703), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n837), .ZN(new_n946));
  XNOR2_X1  g521(.A(KEYINPUT110), .B(G1384), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT111), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT45), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g525(.A(G40), .B(new_n465), .C1(new_n478), .C2(new_n463), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n946), .A2(KEYINPUT111), .A3(new_n947), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n945), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n954), .A2(G1986), .A3(G290), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n955), .A2(G1986), .A3(G290), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n961), .A2(KEYINPUT112), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(KEYINPUT112), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n957), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT113), .B1(new_n837), .B2(G1384), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n967));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n967), .B(new_n968), .C1(new_n502), .C2(new_n834), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n951), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G8), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT117), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n673), .A2(new_n676), .ZN(new_n975));
  NAND2_X1  g550(.A1(G305), .A2(G1981), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n973), .A2(KEYINPUT117), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n977), .B1(new_n980), .B2(new_n974), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n972), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(G288), .A2(G1976), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT118), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n975), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT119), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(KEYINPUT119), .A3(new_n975), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(new_n972), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n966), .A2(new_n991), .A3(new_n969), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n835), .A2(new_n836), .ZN(new_n993));
  INV_X1    g568(.A(new_n506), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n951), .B1(new_n995), .B2(KEYINPUT45), .ZN(new_n996));
  AOI21_X1  g571(.A(G1966), .B1(new_n992), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n966), .A2(new_n999), .A3(new_n969), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n995), .A2(KEYINPUT50), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n952), .A2(new_n783), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n971), .B1(new_n998), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1976), .ZN(new_n1007));
  NOR2_X1   g582(.A1(G288), .A2(new_n1007), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n970), .A2(new_n971), .A3(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT116), .B(G1976), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(G288), .B2(new_n1010), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n1009), .A2(new_n1011), .B1(new_n972), .B2(new_n981), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1008), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n972), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT52), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1006), .A2(new_n1012), .A3(new_n1015), .A4(G168), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1002), .A2(new_n722), .A3(new_n952), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n968), .B1(new_n502), .B2(new_n506), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n991), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT45), .B(new_n947), .C1(new_n502), .C2(new_n834), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n952), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n686), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n971), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(G166), .B2(new_n971), .ZN(new_n1026));
  NAND3_X1  g601(.A1(G303), .A2(G8), .A3(new_n1024), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1023), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT63), .B1(new_n1016), .B2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g606(.A(G2090), .B(new_n951), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n951), .B1(new_n991), .B2(new_n1018), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1971), .B1(new_n1033), .B2(new_n1020), .ZN(new_n1034));
  OAI211_X1 g609(.A(G8), .B(new_n1029), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1038), .A2(KEYINPUT115), .A3(G8), .A4(new_n1029), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1003), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1040));
  OAI211_X1 g615(.A(G8), .B(G168), .C1(new_n997), .C2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(KEYINPUT63), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n966), .A2(KEYINPUT50), .A3(new_n969), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n951), .B1(new_n995), .B2(new_n999), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1022), .B1(new_n1045), .B2(G2090), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G8), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1028), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1037), .A2(new_n1039), .B1(new_n1042), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n970), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1050), .A2(G8), .A3(new_n1013), .A4(new_n1011), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1051), .B(new_n982), .C1(new_n1052), .C2(new_n1009), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n990), .B(new_n1031), .C1(new_n1049), .C2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT56), .B(G2072), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1033), .A2(new_n1020), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1956), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n567), .A2(KEYINPUT120), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n567), .A2(new_n569), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1062), .B1(new_n567), .B2(new_n569), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1061), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1065), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT57), .B1(new_n567), .B2(KEYINPUT120), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n1063), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1057), .A2(new_n1058), .A3(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(new_n597), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1002), .A2(new_n952), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n714), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n970), .A2(new_n938), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1045), .A2(new_n781), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1056), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1070), .A2(KEYINPUT122), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1066), .A2(new_n1069), .A3(new_n1080), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1072), .A2(new_n1076), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT61), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1064), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1068), .B1(new_n1067), .B2(new_n1063), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(new_n1077), .B2(new_n1056), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1084), .B1(new_n1088), .B2(new_n1071), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1079), .B(new_n1081), .C1(new_n1058), .C2(new_n1057), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1077), .A2(new_n1087), .A3(new_n1056), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(KEYINPUT61), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT123), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1019), .A2(new_n952), .A3(new_n940), .A4(new_n1020), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT58), .B(G1341), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1095), .B1(new_n970), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1094), .B1(new_n1097), .B2(new_n557), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1097), .A2(new_n557), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1089), .A2(new_n1092), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n951), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1103));
  OAI211_X1 g678(.A(KEYINPUT60), .B(new_n1075), .C1(new_n1103), .C2(G1348), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1104), .A2(new_n596), .A3(new_n595), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1074), .A2(KEYINPUT60), .A3(new_n597), .A4(new_n1075), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT60), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1105), .A2(new_n1106), .B1(new_n1107), .B2(new_n1076), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1083), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G168), .A2(new_n971), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n998), .A2(new_n1005), .A3(KEYINPUT124), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n997), .B2(new_n1040), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1111), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1114), .A3(G168), .ZN(new_n1116));
  AND2_X1   g691(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1006), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1110), .A2(KEYINPUT51), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1115), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1029), .B1(new_n1046), .B2(G8), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1053), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1033), .A2(new_n795), .A3(new_n1020), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1073), .A2(new_n725), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(G301), .B(KEYINPUT54), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n950), .A2(new_n953), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n795), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n478), .A2(KEYINPUT125), .ZN(new_n1131));
  OAI21_X1  g706(.A(G2105), .B1(new_n478), .B2(KEYINPUT125), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n465), .B(new_n1130), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1020), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1128), .B1(new_n1129), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1125), .B1(new_n1021), .B2(G2078), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n992), .A2(new_n996), .A3(KEYINPUT53), .A4(new_n795), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1137), .B(new_n1138), .C1(new_n1103), .C2(G1961), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1127), .A2(new_n1136), .B1(new_n1139), .B2(new_n1128), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT115), .B1(new_n1023), .B2(new_n1029), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1034), .B1(new_n1103), .B2(new_n722), .ZN(new_n1142));
  NOR4_X1   g717(.A1(new_n1142), .A2(new_n1036), .A3(new_n971), .A4(new_n1028), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1124), .B(new_n1140), .C1(new_n1141), .C2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1122), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1054), .B1(new_n1109), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1139), .A2(G171), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1147), .A2(new_n1124), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1122), .A2(KEYINPUT62), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1116), .A2(new_n1117), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1152), .A2(new_n1153), .A3(new_n1115), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1150), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n965), .B1(new_n1146), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n955), .A2(new_n940), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT46), .ZN(new_n1158));
  INV_X1    g733(.A(new_n939), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n955), .B1(new_n745), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT47), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT48), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n957), .B1(new_n959), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(new_n1163), .B2(new_n959), .ZN(new_n1165));
  INV_X1    g740(.A(new_n942), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1166), .A2(new_n943), .B1(G2067), .B2(new_n762), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n955), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1162), .A2(new_n1165), .A3(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n937), .B1(new_n1156), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1144), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1115), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1109), .A2(new_n1171), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1031), .A2(new_n990), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1042), .A2(new_n1048), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1053), .B1(new_n1147), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1175), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1122), .A2(KEYINPUT62), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1153), .B1(new_n1152), .B2(new_n1115), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1149), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n964), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1162), .A2(new_n1165), .A3(new_n1168), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1184), .A2(KEYINPUT126), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1170), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g762(.A1(G401), .A2(new_n458), .A3(G227), .ZN(new_n1189));
  XNOR2_X1  g763(.A(new_n1189), .B(KEYINPUT127), .ZN(new_n1190));
  NOR2_X1   g764(.A1(G229), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g765(.A1(new_n862), .A2(new_n1191), .A3(new_n928), .ZN(G225));
  INV_X1    g766(.A(G225), .ZN(G308));
endmodule


