//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT64), .Z(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XNOR2_X1  g032(.A(KEYINPUT3), .B(G2104), .ZN(new_n458));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n458), .A2(G137), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT65), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n459), .A2(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n467), .A2(G2105), .B1(G101), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n461), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  NOR2_X1   g046(.A1(new_n465), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G136), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n465), .A2(new_n459), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  INV_X1    g050(.A(G100), .ZN(new_n476));
  AND3_X1   g051(.A1(new_n476), .A2(new_n459), .A3(KEYINPUT66), .ZN(new_n477));
  AOI21_X1  g052(.A(KEYINPUT66), .B1(new_n476), .B2(new_n459), .ZN(new_n478));
  OAI221_X1 g053(.A(G2104), .B1(G112), .B2(new_n459), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n473), .A2(new_n475), .A3(new_n479), .ZN(G162));
  NAND2_X1  g055(.A1(new_n474), .A2(G126), .ZN(new_n481));
  OAI211_X1 g056(.A(G138), .B(new_n459), .C1(new_n463), .C2(new_n464), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n482), .A2(KEYINPUT68), .A3(new_n483), .ZN(new_n484));
  AND2_X1   g059(.A1(KEYINPUT67), .A2(G114), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT67), .A2(G114), .ZN(new_n486));
  OAI21_X1  g061(.A(G2105), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n481), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n482), .A2(KEYINPUT68), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n458), .A2(new_n491), .A3(G138), .A4(new_n459), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n490), .A2(new_n492), .A3(KEYINPUT4), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n489), .A2(new_n493), .ZN(G164));
  INV_X1    g069(.A(G50), .ZN(new_n495));
  INV_X1    g070(.A(G651), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT69), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G651), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT6), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT70), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n502), .A2(new_n504), .A3(G651), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(KEYINPUT5), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n508), .A2(KEYINPUT71), .A3(G543), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT72), .B(G88), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n495), .A2(new_n507), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n497), .A2(new_n499), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n517), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n500), .A2(new_n505), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(new_n511), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n531));
  AND3_X1   g106(.A1(new_n508), .A2(KEYINPUT71), .A3(G543), .ZN(new_n532));
  AOI21_X1  g107(.A(KEYINPUT71), .B1(new_n508), .B2(G543), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n526), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G89), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n525), .A2(new_n528), .A3(new_n530), .A4(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  INV_X1    g113(.A(KEYINPUT75), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT74), .B(G90), .Z(new_n540));
  NAND4_X1  g115(.A1(new_n514), .A2(new_n500), .A3(new_n505), .A4(new_n540), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n500), .A2(new_n505), .A3(G52), .A4(G543), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g118(.A(G64), .B(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(new_n519), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n539), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n541), .A2(new_n542), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n520), .B1(new_n544), .B2(new_n545), .ZN(new_n550));
  NOR3_X1   g125(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT75), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND4_X1  g128(.A1(new_n500), .A2(new_n505), .A3(G43), .A4(G543), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n514), .A2(G81), .A3(new_n500), .A4(new_n505), .ZN(new_n555));
  INV_X1    g130(.A(G68), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n511), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n557), .B1(new_n514), .B2(G56), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n554), .B(new_n555), .C1(new_n558), .C2(new_n520), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n534), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(G651), .A2(new_n568), .B1(new_n535), .B2(G91), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n500), .A2(new_n505), .A3(G53), .A4(G543), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(G299));
  OR2_X1    g147(.A1(new_n517), .A2(new_n521), .ZN(G303));
  NAND2_X1  g148(.A1(new_n535), .A2(G87), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n527), .A2(G49), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(new_n514), .A2(G61), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT76), .Z(new_n581));
  AOI21_X1  g156(.A(new_n520), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(KEYINPUT77), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n506), .A2(G86), .A3(new_n514), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n506), .A2(G48), .A3(G543), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(KEYINPUT77), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(new_n535), .A2(G85), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  OAI221_X1 g166(.A(new_n589), .B1(new_n520), .B2(new_n590), .C1(new_n591), .C2(new_n507), .ZN(G290));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n534), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(G651), .A2(new_n595), .B1(new_n527), .B2(G54), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n506), .A2(KEYINPUT10), .A3(G92), .A4(new_n514), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n514), .A2(G92), .A3(new_n500), .A4(new_n505), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g179(.A(new_n603), .B1(G171), .B2(G868), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT9), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n570), .B(new_n607), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n514), .A2(G91), .A3(new_n500), .A4(new_n505), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n496), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n606), .B1(G868), .B2(new_n612), .ZN(G297));
  OAI21_X1  g188(.A(new_n606), .B1(G868), .B2(new_n612), .ZN(G280));
  AND2_X1   g189(.A1(new_n596), .A2(new_n601), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n560), .ZN(G323));
  XOR2_X1   g195(.A(KEYINPUT78), .B(KEYINPUT11), .Z(new_n621));
  XNOR2_X1  g196(.A(G323), .B(new_n621), .ZN(G282));
  NAND2_X1  g197(.A1(new_n458), .A2(new_n468), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n472), .A2(G135), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n459), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  AND3_X1   g204(.A1(new_n474), .A2(KEYINPUT79), .A3(G123), .ZN(new_n630));
  AOI21_X1  g205(.A(KEYINPUT79), .B1(new_n474), .B2(G123), .ZN(new_n631));
  OAI221_X1 g206(.A(new_n627), .B1(new_n628), .B2(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n626), .A2(G2100), .B1(G2096), .B2(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(G2096), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n633), .B(new_n634), .C1(G2100), .C2(new_n626), .ZN(G156));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2430), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AND3_X1   g214(.A1(new_n639), .A2(KEYINPUT80), .A3(KEYINPUT14), .ZN(new_n640));
  AOI21_X1  g215(.A(KEYINPUT80), .B1(new_n639), .B2(KEYINPUT14), .ZN(new_n641));
  OAI22_X1  g216(.A1(new_n640), .A2(new_n641), .B1(new_n637), .B2(new_n638), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n644), .B(new_n645), .Z(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT81), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n646), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT82), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n654));
  NAND4_X1  g229(.A1(new_n650), .A2(new_n654), .A3(G14), .A4(new_n651), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT83), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT17), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2084), .B(G2090), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n662), .B1(new_n659), .B2(new_n661), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n660), .B2(new_n661), .ZN(new_n665));
  INV_X1    g240(.A(new_n661), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n666), .A2(new_n662), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n659), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n663), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2096), .B(G2100), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n674), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n674), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT85), .Z(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT86), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XOR2_X1   g265(.A(new_n689), .B(new_n690), .Z(new_n691));
  OR2_X1    g266(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n691), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(G229));
  NAND2_X1  g269(.A1(new_n472), .A2(G141), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n474), .A2(G129), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n468), .A2(G105), .ZN(new_n697));
  NAND3_X1  g272(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT26), .Z(new_n699));
  NAND4_X1  g274(.A1(new_n695), .A2(new_n696), .A3(new_n697), .A4(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n702), .B2(G32), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT27), .B(G1996), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT30), .B(G28), .ZN(new_n708));
  OR2_X1    g283(.A1(KEYINPUT31), .A2(G11), .ZN(new_n709));
  NAND2_X1  g284(.A1(KEYINPUT31), .A2(G11), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n708), .A2(new_n702), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n632), .B2(new_n702), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n706), .A2(new_n707), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n702), .A2(G35), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G162), .B2(new_n702), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT29), .B(G2090), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G2084), .ZN(new_n718));
  INV_X1    g293(.A(G34), .ZN(new_n719));
  AOI21_X1  g294(.A(G29), .B1(new_n719), .B2(KEYINPUT24), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(KEYINPUT24), .B2(new_n719), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n470), .B2(new_n702), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n717), .B1(new_n718), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n702), .A2(G26), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT94), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n474), .A2(G128), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT93), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n730));
  INV_X1    g305(.A(G116), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G2105), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n472), .B2(G140), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n726), .B1(new_n734), .B2(G29), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G2067), .ZN(new_n736));
  NAND2_X1  g311(.A1(G115), .A2(G2104), .ZN(new_n737));
  INV_X1    g312(.A(G127), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n465), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n459), .B1(new_n739), .B2(KEYINPUT95), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(KEYINPUT95), .B2(new_n739), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT25), .ZN(new_n742));
  NAND2_X1  g317(.A1(G103), .A2(G2104), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(G2105), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n459), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n472), .A2(G139), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  MUX2_X1   g322(.A(G33), .B(new_n747), .S(G29), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G2072), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n713), .A2(new_n723), .A3(new_n736), .A4(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n722), .A2(new_n718), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT96), .Z(new_n752));
  NOR2_X1   g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G16), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G4), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n615), .B2(new_n754), .ZN(new_n756));
  INV_X1    g331(.A(G1348), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n754), .A2(G19), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n560), .B2(new_n754), .ZN(new_n760));
  OAI22_X1  g335(.A1(new_n748), .A2(G2072), .B1(G1341), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G1341), .B2(new_n760), .ZN(new_n762));
  NOR2_X1   g337(.A1(G286), .A2(new_n754), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT97), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(KEYINPUT97), .B1(G16), .B2(G21), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT98), .B(G1966), .Z(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n702), .A2(G27), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G164), .B2(new_n702), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT100), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n767), .A2(new_n769), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n753), .A2(new_n758), .A3(new_n762), .A4(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n767), .A2(new_n769), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT99), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n773), .A2(new_n770), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n754), .A2(G5), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G171), .B2(new_n754), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(G1961), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n754), .A2(G20), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT23), .Z(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G299), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1956), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G1961), .B2(new_n780), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n777), .A2(new_n778), .A3(new_n781), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n754), .A2(G22), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT91), .Z(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G166), .B2(new_n754), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1971), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n754), .A2(G23), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n577), .B2(new_n754), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT33), .B(G1976), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT89), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n794), .B(new_n796), .Z(new_n797));
  INV_X1    g372(.A(KEYINPUT90), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n794), .B(new_n796), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(KEYINPUT90), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n792), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n754), .A2(G6), .ZN(new_n803));
  INV_X1    g378(.A(G305), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n754), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT88), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(KEYINPUT88), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT32), .B(G1981), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n806), .A2(new_n807), .ZN(new_n810));
  INV_X1    g385(.A(new_n808), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n802), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT34), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n802), .A2(new_n815), .A3(new_n809), .A4(new_n812), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT92), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n472), .A2(G131), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n474), .A2(G119), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n459), .A2(G107), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  MUX2_X1   g397(.A(G25), .B(new_n822), .S(G29), .Z(new_n823));
  XOR2_X1   g398(.A(KEYINPUT35), .B(G1991), .Z(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT87), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n823), .B(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(G16), .A2(G24), .ZN(new_n827));
  INV_X1    g402(.A(G290), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(G16), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n826), .B1(new_n829), .B2(G1986), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G1986), .B2(new_n829), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n816), .A2(new_n817), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n817), .B1(new_n816), .B2(new_n831), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n814), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n836), .B(new_n814), .C1(new_n832), .C2(new_n833), .ZN(new_n837));
  AOI211_X1 g412(.A(new_n775), .B(new_n788), .C1(new_n835), .C2(new_n837), .ZN(G311));
  NAND2_X1  g413(.A1(new_n835), .A2(new_n837), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n788), .A2(new_n775), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(G150));
  NAND4_X1  g416(.A1(new_n500), .A2(new_n505), .A3(G55), .A4(G543), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n514), .A2(G93), .A3(new_n500), .A4(new_n505), .ZN(new_n843));
  INV_X1    g418(.A(G80), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n511), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n514), .B2(G67), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n842), .B(new_n843), .C1(new_n846), .C2(new_n520), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT102), .B(G860), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n615), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n514), .A2(G56), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n519), .B1(new_n854), .B2(new_n557), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n555), .A2(new_n554), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n514), .A2(G67), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n519), .B1(new_n857), .B2(new_n845), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n843), .A2(new_n842), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n855), .A2(new_n856), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n559), .A2(new_n847), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n853), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT101), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n849), .B1(new_n863), .B2(new_n864), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n851), .B1(new_n866), .B2(new_n867), .ZN(G145));
  XNOR2_X1  g443(.A(new_n734), .B(G164), .ZN(new_n869));
  AOI22_X1  g444(.A1(G130), .A2(new_n474), .B1(new_n472), .B2(G142), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n872));
  INV_X1    g447(.A(G118), .ZN(new_n873));
  AOI22_X1  g448(.A1(new_n871), .A2(new_n872), .B1(new_n873), .B2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n872), .B2(new_n871), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n869), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n747), .B(new_n700), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n822), .B(new_n624), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n877), .B(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n470), .B(G162), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(new_n632), .Z(new_n883));
  AOI21_X1  g458(.A(G37), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(new_n883), .B2(new_n881), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g461(.A(G305), .B(G290), .ZN(new_n887));
  NAND2_X1  g462(.A1(G288), .A2(G166), .ZN(new_n888));
  NAND2_X1  g463(.A1(G303), .A2(new_n577), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n888), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n804), .A2(G290), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n828), .A2(G305), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT42), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n559), .A2(new_n847), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n559), .A2(new_n847), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n618), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n615), .A2(G299), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n612), .A2(new_n602), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n615), .A2(G299), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n612), .A2(new_n602), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n901), .A2(KEYINPUT41), .A3(new_n902), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n905), .B1(new_n900), .B2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n896), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(G868), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(G868), .B2(new_n848), .ZN(G295));
  OAI21_X1  g490(.A(new_n914), .B1(G868), .B2(new_n848), .ZN(G331));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n548), .B2(new_n551), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n899), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n547), .A2(new_n539), .A3(new_n542), .A4(new_n541), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT75), .B1(new_n549), .B2(new_n550), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT105), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n923), .A2(G286), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT105), .B1(new_n921), .B2(new_n922), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n862), .A2(new_n925), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n920), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n924), .B1(new_n920), .B2(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n911), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n923), .A2(G286), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n899), .A2(new_n919), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n862), .A2(new_n925), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n920), .A2(new_n924), .A3(new_n926), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n903), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n890), .A2(new_n894), .ZN(new_n937));
  AOI21_X1  g512(.A(G37), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n929), .A2(new_n895), .A3(new_n935), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n929), .A2(new_n895), .A3(new_n935), .A4(KEYINPUT106), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n938), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  XOR2_X1   g518(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n938), .A2(new_n941), .A3(new_n944), .A4(new_n942), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n917), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT107), .B1(new_n943), .B2(KEYINPUT43), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(KEYINPUT44), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n943), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT108), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n927), .A2(new_n928), .A3(new_n904), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n933), .A2(new_n934), .B1(new_n910), .B2(new_n909), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n937), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G37), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n958), .A3(new_n942), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n939), .A2(new_n940), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT43), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n947), .A2(KEYINPUT44), .ZN(new_n964));
  AND4_X1   g539(.A1(KEYINPUT108), .A2(new_n963), .A3(new_n964), .A4(new_n953), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n949), .B1(new_n954), .B2(new_n965), .ZN(G397));
  NAND3_X1  g541(.A1(new_n461), .A2(G40), .A3(new_n469), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n489), .B2(new_n493), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G2067), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n734), .B(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n972), .B1(new_n974), .B2(new_n701), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT46), .B1(new_n972), .B2(G1996), .ZN(new_n976));
  OR3_X1    g551(.A1(new_n972), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n979));
  XNOR2_X1  g554(.A(new_n978), .B(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n974), .A2(new_n972), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT110), .ZN(new_n982));
  INV_X1    g557(.A(new_n972), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n700), .B(G1996), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n824), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n822), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n729), .A2(new_n973), .A3(new_n733), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n972), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n822), .A2(new_n986), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n983), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n985), .A2(new_n992), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n972), .A2(G1986), .A3(G290), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n994), .B(KEYINPUT48), .Z(new_n995));
  AOI211_X1 g570(.A(new_n980), .B(new_n990), .C1(new_n993), .C2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n967), .B1(new_n969), .B2(new_n971), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n490), .A2(new_n492), .A3(KEYINPUT4), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n998), .A2(new_n484), .A3(new_n481), .A4(new_n488), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT111), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n999), .A2(new_n1002), .A3(KEYINPUT45), .A4(new_n970), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n997), .A2(new_n1001), .A3(new_n770), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n1005));
  INV_X1    g580(.A(G1961), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n971), .A2(KEYINPUT50), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n999), .A2(new_n1008), .A3(new_n970), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(new_n968), .A3(new_n1009), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1004), .A2(new_n1005), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n971), .A2(new_n969), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1012), .A2(new_n968), .A3(new_n1000), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1005), .A2(G2078), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(G301), .A3(new_n1015), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n997), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n1014), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1011), .A2(new_n1018), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1019), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT125), .B1(new_n1019), .B2(G171), .ZN(new_n1021));
  OAI211_X1 g596(.A(KEYINPUT54), .B(new_n1016), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1007), .A2(new_n968), .A3(new_n718), .A4(new_n1009), .ZN(new_n1023));
  OAI211_X1 g598(.A(G168), .B(new_n1023), .C1(new_n1013), .C2(new_n769), .ZN(new_n1024));
  NOR2_X1   g599(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1010), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1012), .A2(new_n968), .A3(new_n1000), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1027), .A2(new_n718), .B1(new_n1028), .B2(new_n768), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT124), .ZN(new_n1030));
  AOI21_X1  g605(.A(G168), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(G8), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT124), .B1(new_n1024), .B2(G8), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT51), .B1(new_n1033), .B2(KEYINPUT123), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1981), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n583), .A2(new_n586), .A3(new_n1036), .A4(new_n587), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT113), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT113), .B1(new_n584), .B2(new_n585), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n582), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1037), .B1(new_n1040), .B2(new_n1036), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT49), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n971), .A2(new_n967), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G8), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n577), .B2(G1976), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(new_n1044), .A3(G8), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n577), .A2(G1976), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1044), .A2(new_n1050), .A3(G8), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n971), .A2(new_n967), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1056), .B(new_n1048), .C1(KEYINPUT52), .C2(new_n1050), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1043), .A2(new_n1046), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n1017), .A2(G1971), .B1(G2090), .B2(new_n1010), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G303), .A2(G8), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1060), .B(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1062), .A3(G8), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1060), .B(KEYINPUT55), .ZN(new_n1064));
  INV_X1    g639(.A(G2090), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n997), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1066));
  INV_X1    g641(.A(G1971), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1065), .A2(new_n1027), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1064), .B1(new_n1068), .B2(new_n1055), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1058), .A2(new_n1063), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1019), .A2(G171), .ZN(new_n1072));
  AOI21_X1  g647(.A(G301), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1022), .A2(new_n1035), .A3(new_n1070), .A4(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n569), .A2(new_n571), .A3(KEYINPUT57), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT116), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n569), .A2(new_n571), .A3(new_n1078), .A4(KEYINPUT57), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n608), .B1(KEYINPUT115), .B2(new_n611), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n569), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1082), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT117), .B1(new_n1080), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n611), .A2(KEYINPUT115), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n571), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1081), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1090), .A2(new_n1091), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1087), .A2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT56), .B(G2072), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1017), .A2(new_n1094), .B1(new_n1010), .B2(new_n785), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1093), .A2(KEYINPUT118), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT118), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1010), .A2(new_n757), .B1(new_n1054), .B2(new_n973), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(new_n602), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1095), .B1(new_n1093), .B2(KEYINPUT119), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1087), .A2(new_n1092), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT120), .B1(new_n1098), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1093), .A2(KEYINPUT119), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1095), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n1107), .A3(new_n1103), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1100), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1093), .A2(KEYINPUT118), .A3(new_n1095), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1110), .A2(new_n1111), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1105), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1112), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1093), .A2(KEYINPUT122), .A3(new_n1095), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1108), .A2(new_n1120), .A3(KEYINPUT61), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1099), .A2(KEYINPUT60), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(new_n615), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n1099), .A2(KEYINPUT60), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT58), .B(G1341), .ZN(new_n1126));
  OAI22_X1  g701(.A1(new_n1066), .A2(G1996), .B1(new_n1054), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n560), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT59), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1130), .A3(new_n560), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1124), .A2(new_n1125), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n1135));
  OAI211_X1 g710(.A(new_n1122), .B(new_n1132), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1075), .B1(new_n1118), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1138), .B1(new_n1035), .B2(KEYINPUT62), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n1140));
  AOI211_X1 g715(.A(KEYINPUT126), .B(new_n1140), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1032), .A2(new_n1034), .A3(new_n1140), .ZN(new_n1142));
  AND4_X1   g717(.A1(new_n1073), .A2(new_n1058), .A3(new_n1069), .A4(new_n1063), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1139), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1146));
  INV_X1    g721(.A(G1976), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(new_n1147), .A3(new_n577), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1045), .B1(new_n1148), .B2(new_n1037), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1063), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(new_n1058), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1029), .A2(new_n1055), .A3(G286), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1058), .A2(new_n1063), .A3(new_n1069), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1151), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n1137), .A2(new_n1145), .A3(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(G290), .A2(G1986), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n994), .B1(new_n983), .B2(new_n1159), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n1160), .B(KEYINPUT109), .Z(new_n1161));
  NAND2_X1  g736(.A1(new_n993), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n996), .B1(new_n1158), .B2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g738(.A(G319), .ZN(new_n1165));
  NOR2_X1   g739(.A1(G227), .A2(new_n1165), .ZN(new_n1166));
  AND3_X1   g740(.A1(new_n692), .A2(new_n693), .A3(new_n1166), .ZN(new_n1167));
  NAND3_X1  g741(.A1(new_n656), .A2(new_n1167), .A3(new_n885), .ZN(new_n1168));
  NOR2_X1   g742(.A1(new_n946), .A2(new_n948), .ZN(new_n1169));
  NOR2_X1   g743(.A1(new_n1168), .A2(new_n1169), .ZN(G308));
  INV_X1    g744(.A(G308), .ZN(G225));
endmodule


