//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G113), .B(G122), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(G104), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G140), .ZN(new_n195));
  AND2_X1   g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  OR2_X1    g010(.A1(KEYINPUT64), .A2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT64), .A2(G146), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(new_n196), .ZN(new_n201));
  INV_X1    g015(.A(G237), .ZN(new_n202));
  INV_X1    g016(.A(G953), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G214), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(G237), .A2(G953), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(G143), .A3(G214), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT18), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n206), .A2(new_n208), .B1(KEYINPUT18), .B2(G131), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n201), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT66), .A2(G131), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT66), .A2(G131), .ZN(new_n216));
  OR2_X1    g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n207), .A2(G143), .A3(G214), .ZN(new_n218));
  AOI21_X1  g032(.A(G143), .B1(new_n207), .B2(G214), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT17), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n215), .A2(new_n216), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n206), .A2(new_n222), .A3(new_n208), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT90), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n220), .A2(new_n223), .A3(KEYINPUT90), .A4(new_n221), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT89), .B1(new_n220), .B2(new_n221), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n193), .A2(new_n195), .A3(KEYINPUT16), .ZN(new_n230));
  OR3_X1    g044(.A1(new_n194), .A2(KEYINPUT16), .A3(G140), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n200), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n231), .A3(G146), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT89), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n209), .A2(new_n235), .A3(KEYINPUT17), .A4(new_n217), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n229), .A2(new_n233), .A3(new_n234), .A4(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n214), .B1(new_n228), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT91), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT91), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n240), .B(new_n214), .C1(new_n228), .C2(new_n237), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n191), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT88), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n190), .B(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n214), .B(new_n244), .C1(new_n228), .C2(new_n237), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n188), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G475), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n220), .A2(new_n223), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT19), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n196), .B(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n197), .A2(new_n198), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n249), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT75), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n234), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT75), .A4(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n214), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n190), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n245), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G475), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n188), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT20), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT20), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n260), .A2(new_n265), .A3(new_n262), .A4(new_n188), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G122), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT92), .B1(new_n268), .B2(G116), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT92), .ZN(new_n270));
  INV_X1    g084(.A(G116), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(G122), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n273), .A2(KEYINPUT14), .B1(G116), .B2(new_n268), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(KEYINPUT14), .B2(new_n273), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G107), .ZN(new_n276));
  INV_X1    g090(.A(G107), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT93), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n268), .A2(G116), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n273), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n278), .B1(new_n273), .B2(new_n279), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n277), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G128), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(G143), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT94), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(KEYINPUT68), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G128), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n286), .B1(new_n290), .B2(new_n205), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT68), .B(G128), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(KEYINPUT94), .A3(G143), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n285), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G134), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI211_X1 g110(.A(G134), .B(new_n285), .C1(new_n291), .C2(new_n293), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n276), .B(new_n283), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT9), .B(G234), .ZN(new_n299));
  INV_X1    g113(.A(G217), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n299), .A2(new_n300), .A3(G953), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n285), .A2(KEYINPUT13), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT94), .B1(new_n292), .B2(G143), .ZN(new_n304));
  AND4_X1   g118(.A1(KEYINPUT94), .A2(new_n287), .A3(new_n289), .A4(G143), .ZN(new_n305));
  OAI22_X1  g119(.A1(new_n304), .A2(new_n305), .B1(KEYINPUT13), .B2(new_n285), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n303), .B1(new_n306), .B2(KEYINPUT95), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n285), .A2(KEYINPUT13), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n291), .B2(new_n293), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT95), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n295), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n294), .A2(new_n295), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n281), .A2(new_n277), .A3(new_n282), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n273), .A2(new_n279), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT93), .ZN(new_n316));
  AOI21_X1  g130(.A(G107), .B1(new_n316), .B2(new_n280), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n313), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n298), .B(new_n301), .C1(new_n312), .C2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n302), .B1(new_n309), .B2(new_n310), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n306), .A2(KEYINPUT95), .ZN(new_n322));
  OAI21_X1  g136(.A(G134), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n316), .A2(G107), .A3(new_n280), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n297), .B1(new_n283), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n301), .B1(new_n326), .B2(new_n298), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n188), .B1(new_n320), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G478), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(KEYINPUT15), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n298), .B1(new_n312), .B2(new_n318), .ZN(new_n332));
  INV_X1    g146(.A(new_n301), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(G902), .B1(new_n334), .B2(new_n319), .ZN(new_n335));
  INV_X1    g149(.A(new_n330), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n248), .A2(new_n267), .A3(new_n331), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(G234), .A2(G237), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(G952), .A3(new_n203), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT96), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n339), .A2(G902), .A3(G953), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT21), .B(G898), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n187), .B1(new_n338), .B2(new_n345), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n247), .A2(G475), .B1(new_n264), .B2(new_n266), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n334), .A2(new_n319), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n336), .B1(new_n348), .B2(new_n188), .ZN(new_n349));
  AOI211_X1 g163(.A(G902), .B(new_n330), .C1(new_n334), .C2(new_n319), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n345), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n347), .A2(new_n351), .A3(KEYINPUT97), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n346), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(G221), .B1(new_n299), .B2(G902), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT77), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n357));
  AND2_X1   g171(.A1(KEYINPUT64), .A2(G146), .ZN(new_n358));
  NOR2_X1   g172(.A1(KEYINPUT64), .A2(G146), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n358), .A2(new_n359), .A3(new_n205), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT65), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n361), .B1(new_n200), .B2(G143), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n205), .A2(KEYINPUT65), .A3(G146), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  AND2_X1   g179(.A1(KEYINPUT0), .A2(G128), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n205), .B1(new_n358), .B2(new_n359), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n200), .A2(G143), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(KEYINPUT0), .A2(G128), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n365), .A2(new_n366), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n277), .B2(G104), .ZN(new_n374));
  INV_X1    g188(.A(G104), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(new_n375), .B2(G107), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n277), .A3(G104), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(KEYINPUT78), .A3(G107), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n374), .A2(new_n376), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G101), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n381), .B1(new_n380), .B2(G101), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n374), .A2(new_n379), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n376), .A2(new_n378), .ZN(new_n385));
  INV_X1    g199(.A(G101), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n383), .A2(KEYINPUT79), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT79), .B1(new_n383), .B2(new_n387), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n372), .B(new_n382), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT80), .B1(new_n375), .B2(G107), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n277), .A3(G104), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n375), .A2(G107), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G101), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n284), .B1(new_n368), .B2(KEYINPUT1), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n362), .A2(new_n363), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n197), .A2(G143), .A3(new_n198), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n284), .A2(KEYINPUT1), .ZN(new_n402));
  AND4_X1   g216(.A1(new_n400), .A2(new_n362), .A3(new_n363), .A4(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n387), .B(new_n397), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n380), .A2(G101), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n386), .B1(new_n394), .B2(new_n395), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT10), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n400), .A2(new_n362), .A3(new_n363), .A4(new_n402), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n292), .B1(new_n400), .B2(KEYINPUT1), .ZN(new_n411));
  INV_X1    g225(.A(new_n368), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n252), .B2(new_n205), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n410), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n404), .A2(new_n405), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT11), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n295), .B2(G137), .ZN(new_n417));
  INV_X1    g231(.A(G137), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(KEYINPUT11), .A3(G134), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n295), .A2(G137), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G131), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n222), .A2(new_n419), .A3(new_n420), .A4(new_n417), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT69), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT69), .B1(new_n422), .B2(new_n423), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n390), .A2(new_n415), .A3(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G110), .B(G140), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n203), .A2(G227), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n428), .B(new_n429), .Z(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n357), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n390), .A2(new_n415), .ZN(new_n433));
  INV_X1    g247(.A(new_n426), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n390), .A2(new_n415), .A3(new_n426), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(KEYINPUT83), .A3(new_n430), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n432), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  OAI221_X1 g252(.A(new_n410), .B1(new_n411), .B2(new_n413), .C1(new_n406), .C2(new_n407), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT82), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n439), .A2(new_n440), .A3(new_n404), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n440), .A2(KEYINPUT12), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(new_n439), .B2(new_n404), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n434), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n439), .A2(new_n404), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n422), .A2(new_n423), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT12), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n436), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n431), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n438), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n188), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G469), .ZN(new_n453));
  INV_X1    g267(.A(G469), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n426), .B1(new_n390), .B2(new_n415), .ZN(new_n455));
  OAI211_X1 g269(.A(KEYINPUT84), .B(new_n431), .C1(new_n427), .C2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n444), .A2(new_n436), .A3(new_n448), .A4(new_n430), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n435), .A2(new_n436), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT84), .B1(new_n459), .B2(new_n431), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n454), .B(new_n188), .C1(new_n458), .C2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n356), .B1(new_n453), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G214), .B1(G237), .B2(G902), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G110), .B(G122), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G113), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n271), .A2(G119), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT5), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G119), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G116), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n271), .A2(G119), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT5), .ZN(new_n475));
  XNOR2_X1  g289(.A(G116), .B(G119), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n468), .A2(KEYINPUT2), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT2), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G113), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n471), .A2(new_n475), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n397), .A2(new_n387), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n397), .B2(new_n387), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n471), .A2(new_n475), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n480), .A2(new_n476), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n488), .B(new_n484), .C1(new_n406), .C2(new_n407), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n467), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n372), .A2(G125), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n414), .A2(new_n194), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n203), .A2(G224), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(KEYINPUT7), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(KEYINPUT7), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n492), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n491), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n480), .B(new_n476), .Z(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n501), .B(new_n382), .C1(new_n388), .C2(new_n389), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n502), .A2(new_n482), .A3(new_n465), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n188), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n502), .A2(new_n482), .ZN(new_n507));
  INV_X1    g321(.A(new_n465), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n502), .A2(new_n482), .A3(new_n465), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(KEYINPUT6), .A3(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n494), .B(new_n495), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n507), .A2(new_n513), .A3(new_n508), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(KEYINPUT87), .B(new_n188), .C1(new_n499), .C2(new_n503), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n506), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G210), .B1(G237), .B2(G902), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n506), .A2(new_n515), .A3(new_n518), .A4(new_n516), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n464), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n354), .A2(new_n462), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n372), .B1(new_n424), .B2(new_n425), .ZN(new_n524));
  INV_X1    g338(.A(new_n421), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n418), .A2(KEYINPUT67), .A3(G134), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT67), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n527), .B1(new_n295), .B2(G137), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n295), .A2(G137), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n525), .A2(new_n222), .B1(new_n530), .B2(G131), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n414), .A2(new_n531), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n524), .A2(new_n500), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n369), .A2(new_n371), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n399), .A2(new_n400), .A3(new_n366), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT69), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n446), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT69), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n414), .A2(new_n531), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT30), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT30), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n446), .A2(new_n535), .A3(new_n534), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n532), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n533), .B1(new_n546), .B2(new_n501), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n202), .A2(new_n203), .A3(G210), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT27), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT70), .ZN(new_n551));
  XOR2_X1   g365(.A(KEYINPUT26), .B(G101), .Z(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT72), .B1(new_n547), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT29), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT72), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n500), .B1(new_n542), .B2(new_n545), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n557), .B(new_n553), .C1(new_n558), .C2(new_n533), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n500), .B1(new_n532), .B2(new_n544), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT28), .B1(new_n533), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT71), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n540), .B2(new_n541), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n524), .A2(KEYINPUT71), .A3(new_n532), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n501), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n561), .B(new_n554), .C1(new_n565), .C2(KEYINPUT28), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n555), .A2(new_n556), .A3(new_n559), .A4(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n500), .B1(new_n524), .B2(new_n532), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT28), .B1(new_n533), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n553), .A2(new_n556), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n569), .B(new_n570), .C1(new_n565), .C2(KEYINPUT28), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n188), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT73), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT73), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n574), .A3(new_n188), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n567), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G472), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT32), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n543), .B1(new_n524), .B2(new_n532), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n532), .A2(new_n543), .A3(new_n544), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n501), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n533), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n554), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT31), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n581), .A2(new_n554), .A3(KEYINPUT31), .A4(new_n582), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n561), .B1(new_n565), .B2(KEYINPUT28), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n553), .ZN(new_n589));
  AOI21_X1  g403(.A(G902), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G472), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n578), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n585), .A2(new_n586), .B1(new_n553), .B2(new_n588), .ZN(new_n593));
  NOR4_X1   g407(.A1(new_n593), .A2(KEYINPUT32), .A3(G472), .A4(G902), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n577), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT22), .B(G137), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n596), .A2(KEYINPUT76), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(KEYINPUT76), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n203), .A2(G221), .A3(G234), .ZN(new_n599));
  OR3_X1    g413(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n599), .B1(new_n597), .B2(new_n598), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT24), .B(G110), .Z(new_n604));
  NAND3_X1  g418(.A1(new_n287), .A2(new_n289), .A3(G119), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n284), .A2(G119), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n230), .A2(G146), .A3(new_n231), .ZN(new_n609));
  AOI21_X1  g423(.A(G146), .B1(new_n230), .B2(new_n231), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT74), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n287), .A2(new_n289), .A3(KEYINPUT23), .A4(G119), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT23), .B1(new_n284), .B2(G119), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n284), .A2(G119), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n612), .B1(new_n617), .B2(G110), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(G110), .ZN(new_n620));
  AOI211_X1 g434(.A(KEYINPUT74), .B(new_n620), .C1(new_n613), .C2(new_n616), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n611), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n613), .A2(new_n620), .A3(new_n616), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n604), .B1(new_n605), .B2(new_n607), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n199), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n257), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n603), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n233), .A2(new_n234), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n629), .B(new_n608), .C1(new_n618), .C2(new_n621), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n606), .B1(new_n292), .B2(G119), .ZN(new_n631));
  OAI22_X1  g445(.A1(new_n617), .A2(G110), .B1(new_n631), .B2(new_n604), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n632), .A2(new_n255), .A3(new_n256), .A4(new_n199), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n630), .A2(new_n633), .A3(new_n602), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n300), .B1(G234), .B2(new_n188), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(G902), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT25), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n630), .A2(new_n633), .A3(new_n602), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n602), .B1(new_n630), .B2(new_n633), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n639), .B(new_n188), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n636), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n639), .B1(new_n635), .B2(new_n188), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n638), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n595), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n523), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(new_n386), .ZN(G3));
  AOI211_X1 g463(.A(new_n345), .B(new_n464), .C1(new_n520), .C2(new_n521), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n248), .A2(new_n267), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT98), .B1(new_n320), .B2(new_n327), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT33), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n348), .A2(KEYINPUT98), .A3(KEYINPUT33), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n329), .A2(G902), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n335), .A2(G478), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n650), .A2(new_n651), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n590), .A2(new_n591), .ZN(new_n664));
  OAI21_X1  g478(.A(G472), .B1(new_n593), .B2(G902), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n664), .A2(new_n646), .A3(new_n665), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n666), .A2(new_n462), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT99), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT34), .B(G104), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G6));
  NOR2_X1   g485(.A1(new_n651), .A2(new_n351), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n522), .A2(new_n352), .A3(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n673), .A2(KEYINPUT100), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(KEYINPUT100), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n667), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT35), .B(G107), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  NAND2_X1  g493(.A1(new_n630), .A2(new_n633), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n602), .A2(KEYINPUT36), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n637), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n683), .B1(new_n643), .B2(new_n644), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n664), .A2(new_n665), .A3(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n354), .A2(new_n685), .A3(new_n462), .A4(new_n522), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  INV_X1    g502(.A(new_n684), .ZN(new_n689));
  AOI211_X1 g503(.A(new_n464), .B(new_n689), .C1(new_n520), .C2(new_n521), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n595), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n356), .ZN(new_n692));
  INV_X1    g506(.A(new_n461), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n454), .B1(new_n451), .B2(new_n188), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(G900), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n342), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n341), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n651), .A2(new_n351), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G128), .ZN(G30));
  XOR2_X1   g516(.A(new_n699), .B(KEYINPUT39), .Z(new_n703));
  NAND2_X1  g517(.A1(new_n462), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT40), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n704), .B(KEYINPUT102), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT40), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n592), .A2(new_n594), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n553), .B1(new_n533), .B2(new_n568), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n583), .A2(G472), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(G472), .A2(G902), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT101), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n520), .A2(new_n521), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT38), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n463), .B1(new_n349), .B2(new_n350), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n347), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n689), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n718), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n708), .A2(new_n710), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT103), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G143), .ZN(G45));
  INV_X1    g542(.A(new_n699), .ZN(new_n729));
  INV_X1    g543(.A(new_n657), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n654), .B2(new_n655), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n651), .B(new_n729), .C1(new_n731), .C2(new_n659), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n696), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G146), .ZN(G48));
  OAI21_X1  g549(.A(new_n188), .B1(new_n458), .B2(new_n460), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(G469), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n737), .A2(new_n692), .A3(new_n461), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n595), .A2(new_n646), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n662), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT41), .B(G113), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  AOI21_X1  g556(.A(new_n739), .B1(new_n674), .B2(new_n675), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n271), .ZN(G18));
  NAND4_X1  g558(.A1(new_n595), .A2(new_n354), .A3(new_n690), .A4(new_n738), .ZN(new_n745));
  XOR2_X1   g559(.A(KEYINPUT104), .B(G119), .Z(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G21));
  NAND4_X1  g561(.A1(new_n737), .A2(new_n692), .A3(new_n461), .A4(new_n352), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n569), .B1(new_n565), .B2(KEYINPUT28), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n553), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n587), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(G472), .A2(G902), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n645), .A2(KEYINPUT105), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n755), .B(new_n638), .C1(new_n643), .C2(new_n644), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n665), .A2(new_n753), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n748), .A2(new_n758), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n719), .A2(KEYINPUT106), .A3(new_n723), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT106), .B1(new_n719), .B2(new_n723), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n665), .A2(new_n753), .A3(new_n684), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n733), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n738), .A2(new_n522), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n764), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n765), .A2(new_n732), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n770), .A2(KEYINPUT107), .A3(new_n522), .A4(new_n738), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G125), .ZN(G27));
  NAND2_X1  g587(.A1(new_n595), .A2(new_n757), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n520), .A2(new_n463), .A3(new_n521), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n733), .A2(new_n462), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT42), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n695), .A2(new_n775), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n732), .A2(KEYINPUT42), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n595), .A3(new_n646), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n211), .ZN(G33));
  NAND4_X1  g597(.A1(new_n779), .A2(new_n595), .A3(new_n646), .A4(new_n700), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G134), .ZN(G36));
  XOR2_X1   g599(.A(new_n775), .B(KEYINPUT108), .Z(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n661), .A2(new_n347), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT43), .Z(new_n789));
  AOI21_X1  g603(.A(new_n689), .B1(new_n664), .B2(new_n665), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n787), .B1(new_n791), .B2(KEYINPUT44), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(KEYINPUT44), .B2(new_n791), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n451), .B(KEYINPUT45), .ZN(new_n794));
  OAI21_X1  g608(.A(G469), .B1(new_n794), .B2(G902), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n693), .B1(new_n795), .B2(KEYINPUT46), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(KEYINPUT46), .B2(new_n795), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n692), .A3(new_n703), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  NAND2_X1  g614(.A1(new_n797), .A2(new_n692), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT47), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n733), .A2(new_n776), .A3(new_n645), .ZN(new_n803));
  OR3_X1    g617(.A1(new_n802), .A2(new_n595), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  INV_X1    g619(.A(new_n341), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n789), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n758), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n721), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n738), .A2(new_n464), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT114), .Z(new_n812));
  NOR3_X1   g626(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n813), .B(new_n814), .Z(new_n815));
  AND2_X1   g629(.A1(new_n737), .A2(new_n461), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n356), .ZN(new_n817));
  AOI211_X1 g631(.A(new_n787), .B(new_n809), .C1(new_n802), .C2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n738), .A2(new_n776), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n807), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n718), .A3(new_n646), .A4(new_n806), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(KEYINPUT116), .Z(new_n823));
  NOR2_X1   g637(.A1(new_n661), .A2(new_n651), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n766), .A2(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n815), .A2(KEYINPUT51), .A3(new_n819), .A4(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n823), .A2(new_n651), .A3(new_n661), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n821), .A2(new_n595), .A3(new_n757), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT48), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n809), .A2(new_n768), .ZN(new_n830));
  INV_X1    g644(.A(G952), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n830), .A2(new_n831), .A3(G953), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n826), .A2(new_n827), .A3(new_n829), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n815), .A2(new_n825), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n834), .B1(new_n835), .B2(new_n818), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT117), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n838), .B(new_n834), .C1(new_n835), .C2(new_n818), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n833), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n686), .B1(new_n523), .B2(new_n647), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n740), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n762), .A2(new_n745), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n666), .A2(new_n650), .A3(new_n462), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n651), .B1(new_n731), .B2(new_n659), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT110), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g661(.A(KEYINPUT110), .B(new_n651), .C1(new_n731), .C2(new_n659), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n672), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n739), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n676), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n842), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n338), .A2(new_n689), .A3(new_n699), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n595), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n779), .B1(new_n856), .B2(new_n770), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(new_n778), .A3(new_n781), .A4(new_n784), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT111), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n691), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(new_n462), .C1(new_n700), .C2(new_n733), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n695), .A2(new_n684), .A3(new_n699), .ZN(new_n862));
  OAI221_X1 g676(.A(new_n862), .B1(new_n711), .B2(new_n717), .C1(new_n761), .C2(new_n760), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n772), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n861), .A2(new_n772), .A3(new_n863), .A4(KEYINPUT52), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n743), .A2(new_n841), .A3(new_n740), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n770), .B1(new_n595), .B2(new_n855), .ZN(new_n870));
  INV_X1    g684(.A(new_n779), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n784), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n782), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT111), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n869), .A2(new_n873), .A3(new_n874), .A4(new_n851), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n859), .A2(new_n868), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n876), .B(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT54), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n876), .A2(new_n877), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT112), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT112), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n876), .A2(new_n882), .A3(new_n877), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT113), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n866), .A2(new_n867), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n842), .A2(new_n851), .A3(new_n853), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(KEYINPUT53), .A3(new_n873), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n884), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n854), .A2(new_n877), .A3(new_n858), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n889), .A2(KEYINPUT113), .A3(new_n868), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n881), .A2(new_n883), .A3(new_n891), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n892), .A2(KEYINPUT54), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n840), .A2(new_n879), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(G952), .B2(G953), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n757), .A2(new_n692), .A3(new_n463), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n788), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n810), .B1(new_n897), .B2(KEYINPUT109), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n897), .A2(KEYINPUT109), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n816), .B(KEYINPUT49), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n898), .A2(new_n899), .A3(new_n718), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n895), .A2(new_n901), .ZN(G75));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n892), .A2(G210), .A3(G902), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n511), .A2(new_n514), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n512), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT55), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n903), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n909), .ZN(new_n911));
  AOI211_X1 g725(.A(KEYINPUT118), .B(new_n911), .C1(new_n904), .C2(new_n905), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n905), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n914), .B1(new_n904), .B2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n892), .A2(KEYINPUT119), .A3(G210), .A4(G902), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n203), .A2(G952), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT120), .B1(new_n913), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n919), .B1(new_n916), .B2(new_n917), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n923), .B(new_n924), .C1(new_n910), .C2(new_n912), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n922), .A2(new_n925), .ZN(G51));
  XNOR2_X1  g740(.A(new_n892), .B(KEYINPUT54), .ZN(new_n927));
  NAND2_X1  g741(.A1(G469), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT57), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT121), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n458), .A2(new_n460), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n927), .A2(new_n933), .A3(new_n929), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n892), .A2(G902), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n936), .A2(G469), .A3(new_n794), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n919), .B1(new_n935), .B2(new_n937), .ZN(G54));
  NAND3_X1  g752(.A1(new_n936), .A2(KEYINPUT58), .A3(G475), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n939), .A2(new_n261), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n261), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n941), .A3(new_n919), .ZN(G60));
  NAND2_X1  g756(.A1(new_n893), .A2(new_n879), .ZN(new_n943));
  NAND2_X1  g757(.A1(G478), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT59), .Z(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n656), .B(KEYINPUT122), .Z(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(KEYINPUT123), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n945), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n919), .B1(new_n927), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT123), .B1(new_n947), .B2(new_n949), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(G63));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT60), .Z(new_n957));
  AOI21_X1  g771(.A(new_n635), .B1(new_n892), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(new_n919), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n892), .A2(new_n682), .A3(new_n957), .ZN(new_n960));
  AOI22_X1  g774(.A1(new_n959), .A2(new_n960), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n961));
  NOR2_X1   g775(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G66));
  NAND2_X1  g777(.A1(G224), .A2(G953), .ZN(new_n964));
  OAI22_X1  g778(.A1(new_n854), .A2(G953), .B1(new_n343), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(G898), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n907), .B1(new_n966), .B2(G953), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n965), .B(new_n967), .ZN(G69));
  XNOR2_X1  g782(.A(new_n546), .B(new_n251), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(G900), .B2(G953), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n861), .A2(new_n772), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n799), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n778), .A2(new_n781), .A3(new_n784), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT126), .Z(new_n974));
  NOR2_X1   g788(.A1(new_n760), .A2(new_n761), .ZN(new_n975));
  OR3_X1    g789(.A1(new_n798), .A2(new_n975), .A3(new_n774), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n972), .A2(new_n804), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n970), .B1(new_n977), .B2(G953), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT125), .ZN(new_n979));
  OR4_X1    g793(.A1(new_n647), .A2(new_n709), .A3(new_n775), .A4(new_n849), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n799), .A2(new_n804), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n727), .A2(KEYINPUT62), .A3(new_n971), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n727), .A2(new_n971), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n981), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n986), .A2(G953), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n979), .B1(new_n987), .B2(new_n969), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n979), .B(new_n969), .C1(new_n986), .C2(G953), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n978), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n203), .B1(G227), .B2(G900), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n992), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n994), .B(new_n978), .C1(new_n988), .C2(new_n990), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n993), .A2(new_n995), .ZN(G72));
  NAND2_X1  g810(.A1(new_n986), .A2(new_n886), .ZN(new_n997));
  XNOR2_X1  g811(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(new_n714), .ZN(new_n999));
  AOI211_X1 g813(.A(new_n553), .B(new_n547), .C1(new_n997), .C2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n999), .B1(new_n977), .B2(new_n854), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n1001), .A2(new_n553), .A3(new_n547), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n555), .A2(new_n559), .A3(new_n583), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n878), .A2(new_n999), .A3(new_n1003), .ZN(new_n1004));
  NOR4_X1   g818(.A1(new_n1000), .A2(new_n1002), .A3(new_n919), .A4(new_n1004), .ZN(G57));
endmodule


