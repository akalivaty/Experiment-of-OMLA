//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT72), .ZN(new_n204));
  XNOR2_X1  g003(.A(G71gat), .B(G99gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT71), .ZN(new_n208));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G183gat), .ZN(new_n212));
  INV_X1    g011(.A(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT67), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(G169gat), .A3(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n216), .A2(new_n221), .A3(new_n223), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT25), .ZN(new_n227));
  NOR2_X1   g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  AND2_X1   g027(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(G190gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n209), .A2(KEYINPUT65), .A3(new_n210), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT66), .B1(new_n222), .B2(KEYINPUT23), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G169gat), .ZN(new_n237));
  INV_X1    g036(.A(G176gat), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n237), .A2(new_n238), .A3(KEYINPUT66), .A4(KEYINPUT23), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT25), .B1(G169gat), .B2(G176gat), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n239), .A2(new_n225), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n234), .A2(new_n236), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT26), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n217), .B1(new_n222), .B2(new_n244), .ZN(new_n245));
  NOR3_X1   g044(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n209), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT27), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(G183gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n212), .A2(KEYINPUT27), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n212), .A2(KEYINPUT27), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n249), .A2(G183gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT68), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT28), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(G190gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n252), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n253), .A2(new_n254), .A3(new_n213), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n256), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n247), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n208), .B1(new_n243), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n260), .ZN(new_n263));
  INV_X1    g062(.A(new_n247), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n239), .A2(new_n225), .A3(new_n240), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(new_n235), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n267), .A2(new_n234), .B1(new_n226), .B2(KEYINPUT25), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n268), .A3(KEYINPUT71), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270));
  INV_X1    g069(.A(G113gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(G120gat), .ZN(new_n272));
  INV_X1    g071(.A(G120gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(G113gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n270), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G127gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT70), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G127gat), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n277), .A2(new_n279), .A3(G134gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(new_n276), .B2(G134gat), .ZN(new_n282));
  INV_X1    g081(.A(G134gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n275), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G127gat), .B(G134gat), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n287), .B(new_n270), .C1(new_n272), .C2(new_n274), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n262), .A2(new_n269), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G227gat), .A2(G233gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT64), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n265), .A2(new_n268), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n286), .A2(new_n288), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(new_n208), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n290), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n207), .B1(new_n296), .B2(KEYINPUT32), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT33), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n206), .A2(KEYINPUT33), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n296), .A2(KEYINPUT32), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT73), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n296), .A2(new_n303), .A3(KEYINPUT32), .A4(new_n300), .ZN(new_n304));
  AOI221_X4 g103(.A(KEYINPUT34), .B1(new_n297), .B2(new_n299), .C1(new_n302), .C2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT34), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n302), .A2(new_n304), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n297), .A2(new_n299), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n290), .A2(new_n295), .ZN(new_n310));
  INV_X1    g109(.A(new_n292), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR3_X1   g111(.A1(new_n305), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n312), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n307), .A2(new_n308), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT34), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n307), .A2(new_n306), .A3(new_n308), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n202), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n314), .A3(new_n317), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n312), .B1(new_n305), .B2(new_n309), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT36), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G225gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT4), .ZN(new_n325));
  AND2_X1   g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT78), .ZN(new_n329));
  XNOR2_X1  g128(.A(G141gat), .B(G148gat), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(KEYINPUT2), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n328), .B1(new_n330), .B2(KEYINPUT2), .ZN(new_n332));
  INV_X1    g131(.A(G148gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT79), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT79), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G148gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n336), .A3(G141gat), .ZN(new_n337));
  INV_X1    g136(.A(G141gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G148gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n327), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n341), .B1(new_n342), .B2(KEYINPUT2), .ZN(new_n343));
  AOI22_X1  g142(.A1(KEYINPUT78), .A2(new_n332), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n294), .A2(new_n325), .A3(new_n331), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n343), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n333), .A2(G141gat), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT2), .B1(new_n339), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n342), .A2(new_n341), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT78), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(new_n331), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT4), .B1(new_n351), .B2(new_n289), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n346), .A2(new_n350), .A3(new_n354), .A4(new_n331), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n351), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n289), .B1(new_n358), .B2(new_n354), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n324), .B(new_n353), .C1(new_n357), .C2(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n344), .A2(new_n331), .A3(new_n286), .A4(new_n288), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n351), .A2(new_n289), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n324), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT5), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G1gat), .B(G29gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(KEYINPUT0), .ZN(new_n369));
  XNOR2_X1  g168(.A(G57gat), .B(G85gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n344), .A2(new_n356), .A3(new_n354), .A4(new_n331), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n355), .A2(KEYINPUT80), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n294), .B1(KEYINPUT3), .B2(new_n351), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n374), .A2(new_n375), .B1(new_n345), .B2(new_n352), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(KEYINPUT5), .A3(new_n324), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n367), .A2(new_n371), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT6), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n371), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n374), .A2(new_n375), .ZN(new_n382));
  AND4_X1   g181(.A1(KEYINPUT5), .A2(new_n382), .A3(new_n324), .A4(new_n353), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT5), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n384), .B1(new_n363), .B2(new_n364), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(new_n376), .B2(new_n324), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n381), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n371), .B1(new_n367), .B2(new_n377), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT81), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n380), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  OR2_X1    g191(.A1(new_n378), .A2(new_n379), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n243), .A2(new_n261), .ZN(new_n395));
  INV_X1    g194(.A(G226gat), .ZN(new_n396));
  INV_X1    g195(.A(G233gat), .ZN(new_n397));
  OAI22_X1  g196(.A1(new_n395), .A2(KEYINPUT29), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT22), .ZN(new_n399));
  INV_X1    g198(.A(G211gat), .ZN(new_n400));
  INV_X1    g199(.A(G218gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G197gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT74), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT74), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(G197gat), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n404), .A2(new_n406), .A3(G204gat), .ZN(new_n407));
  AOI21_X1  g206(.A(G204gat), .B1(new_n404), .B2(new_n406), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n402), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(G211gat), .B(G218gat), .Z(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n410), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n412), .B(new_n402), .C1(new_n407), .C2(new_n408), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT75), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n411), .A2(KEYINPUT75), .A3(new_n413), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n396), .A2(new_n397), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT76), .B1(new_n293), .B2(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT76), .B(new_n419), .C1(new_n243), .C2(new_n261), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n398), .B(new_n418), .C1(new_n420), .C2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n419), .B1(new_n243), .B2(new_n261), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n265), .B2(new_n268), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(new_n419), .ZN(new_n426));
  INV_X1    g225(.A(new_n417), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT75), .B1(new_n411), .B2(new_n413), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G8gat), .B(G36gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(G64gat), .B(G92gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  NAND3_X1  g232(.A1(new_n423), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT77), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT30), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n423), .A2(new_n430), .A3(KEYINPUT77), .A4(new_n433), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n433), .B1(new_n423), .B2(new_n430), .ZN(new_n440));
  INV_X1    g239(.A(new_n434), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n440), .B1(new_n441), .B2(KEYINPUT30), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n394), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G78gat), .B(G106gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(G22gat), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT82), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n411), .A2(new_n449), .A3(new_n413), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n409), .A2(KEYINPUT82), .A3(new_n410), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT29), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n354), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n454), .A2(new_n351), .B1(G228gat), .B2(G233gat), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n429), .B(KEYINPUT83), .C1(new_n357), .C2(KEYINPUT29), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT29), .B1(new_n372), .B2(new_n373), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n457), .B1(new_n458), .B2(new_n418), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n455), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT3), .B1(new_n414), .B2(new_n452), .ZN(new_n461));
  OAI22_X1  g260(.A1(new_n458), .A2(new_n418), .B1(new_n358), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(G228gat), .A3(G233gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT31), .B(G50gat), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n460), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n460), .B2(new_n463), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n448), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n460), .A2(new_n463), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n464), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n460), .A2(new_n463), .A3(new_n465), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n447), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n445), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT84), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n376), .A2(new_n324), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT39), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n371), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n361), .A2(new_n324), .A3(new_n362), .ZN(new_n479));
  OAI211_X1 g278(.A(KEYINPUT39), .B(new_n479), .C1(new_n376), .C2(new_n324), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(KEYINPUT40), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n378), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT40), .B1(new_n478), .B2(new_n480), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n473), .B1(new_n443), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n426), .B2(new_n418), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n398), .B(new_n429), .C1(new_n420), .C2(new_n422), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT38), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n433), .A2(new_n486), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n489), .B1(new_n440), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n491), .A2(new_n436), .A3(new_n438), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n440), .A2(new_n490), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n486), .B1(new_n423), .B2(new_n430), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT38), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n492), .A2(new_n392), .A3(new_n393), .A4(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n475), .B1(new_n485), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n473), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n484), .A2(new_n443), .ZN(new_n499));
  AND4_X1   g298(.A1(new_n475), .A2(new_n496), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n323), .B(new_n474), .C1(new_n497), .C2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n313), .A2(new_n318), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT85), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n394), .A2(new_n444), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT35), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n502), .A2(new_n505), .A3(new_n506), .A4(new_n498), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n498), .A2(new_n320), .A3(new_n321), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT35), .B1(new_n508), .B2(new_n504), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n501), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT86), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT86), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n501), .A2(new_n513), .A3(new_n510), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT16), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(G1gat), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(G1gat), .B2(new_n515), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G8gat), .ZN(new_n519));
  INV_X1    g318(.A(G8gat), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n517), .B(new_n520), .C1(G1gat), .C2(new_n515), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G43gat), .B(G50gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT89), .ZN(new_n524));
  OR2_X1    g323(.A1(G43gat), .A2(G50gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n526));
  NAND2_X1  g325(.A1(G43gat), .A2(G50gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(KEYINPUT15), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT14), .ZN(new_n530));
  INV_X1    g329(.A(G29gat), .ZN(new_n531));
  INV_X1    g330(.A(G36gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G29gat), .A2(G36gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT90), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT90), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n538), .A2(G29gat), .A3(G36gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n535), .B(new_n540), .C1(KEYINPUT15), .C2(new_n523), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n529), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n534), .A2(new_n533), .B1(new_n537), .B2(new_n539), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n543), .A2(KEYINPUT15), .A3(new_n528), .A4(new_n524), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n542), .A2(new_n544), .A3(KEYINPUT17), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT17), .B1(new_n542), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n522), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n542), .A2(new_n544), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n519), .A2(new_n521), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n547), .A2(KEYINPUT18), .A3(new_n548), .A4(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n548), .B(KEYINPUT13), .Z(new_n554));
  NOR2_X1   g353(.A1(new_n522), .A2(new_n549), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n550), .A2(new_n551), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n547), .A2(new_n548), .A3(new_n552), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT18), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT92), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(new_n560), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT92), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G169gat), .B(G197gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT12), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT12), .ZN(new_n572));
  INV_X1    g371(.A(new_n569), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n568), .A2(new_n573), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n563), .A2(new_n565), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT91), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT88), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n571), .A2(new_n580), .A3(new_n576), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(new_n571), .B2(new_n576), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n579), .B(new_n583), .C1(new_n561), .C2(new_n558), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n564), .A2(new_n557), .A3(new_n553), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n579), .B1(new_n586), .B2(new_n583), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n578), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n512), .A2(new_n514), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n394), .ZN(new_n590));
  XOR2_X1   g389(.A(G57gat), .B(G64gat), .Z(new_n591));
  INV_X1    g390(.A(KEYINPUT9), .ZN(new_n592));
  INV_X1    g391(.A(G71gat), .ZN(new_n593));
  INV_X1    g392(.A(G78gat), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G71gat), .B(G78gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G127gat), .B(G155gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n522), .B1(new_n599), .B2(new_n598), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT93), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n604), .A2(new_n610), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G99gat), .B(G106gat), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(G85gat), .ZN(new_n616));
  INV_X1    g415(.A(G92gat), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT94), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT94), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(G85gat), .A3(G92gat), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n618), .A2(KEYINPUT7), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  AOI22_X1  g421(.A1(KEYINPUT8), .A2(new_n622), .B1(new_n616), .B2(new_n617), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT7), .ZN(new_n624));
  OAI211_X1 g423(.A(KEYINPUT94), .B(new_n624), .C1(new_n616), .C2(new_n617), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g425(.A(KEYINPUT95), .B(new_n615), .C1(new_n621), .C2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n615), .B1(new_n621), .B2(new_n626), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n618), .A2(KEYINPUT7), .A3(new_n620), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n630), .A2(new_n614), .A3(new_n625), .A4(new_n623), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n627), .B(new_n632), .C1(new_n545), .C2(new_n546), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n627), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n550), .ZN(new_n635));
  NAND3_X1  g434(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G190gat), .B(G218gat), .Z(new_n638));
  OR2_X1    g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  XOR2_X1   g439(.A(G134gat), .B(G162gat), .Z(new_n641));
  AOI21_X1  g440(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT96), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n639), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n639), .A2(new_n640), .B1(KEYINPUT96), .B2(new_n643), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n613), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n613), .A2(new_n647), .A3(KEYINPUT97), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT98), .Z(new_n654));
  NAND3_X1  g453(.A1(new_n632), .A2(new_n598), .A3(new_n627), .ZN(new_n655));
  INV_X1    g454(.A(new_n597), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n596), .B(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(new_n628), .A3(new_n631), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n655), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n634), .A2(KEYINPUT10), .A3(new_n657), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n654), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n655), .A2(new_n658), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n654), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G120gat), .B(G148gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(G176gat), .B(G204gat), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n667), .B(new_n668), .Z(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n663), .A2(new_n665), .A3(new_n669), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n652), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n589), .A2(new_n590), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT99), .B(G1gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1324gat));
  NAND4_X1  g477(.A1(new_n512), .A2(new_n514), .A3(new_n588), .A4(new_n675), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT16), .B(G8gat), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n679), .A2(new_n444), .A3(new_n680), .ZN(new_n681));
  OR3_X1    g480(.A1(new_n681), .A2(KEYINPUT100), .A3(KEYINPUT42), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT100), .B1(new_n681), .B2(KEYINPUT42), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n589), .A2(new_n443), .A3(new_n675), .ZN(new_n684));
  AOI22_X1  g483(.A1(KEYINPUT42), .A2(new_n681), .B1(new_n684), .B2(G8gat), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(G1325gat));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT36), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT36), .B1(new_n320), .B2(new_n321), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n319), .A2(KEYINPUT101), .A3(new_n322), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G15gat), .B1(new_n679), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n502), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n695), .A2(G15gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n679), .B2(new_n696), .ZN(G1326gat));
  OR3_X1    g496(.A1(new_n679), .A2(KEYINPUT102), .A3(new_n498), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT102), .B1(new_n679), .B2(new_n498), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT43), .B(G22gat), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(G1327gat));
  OAI21_X1  g504(.A(new_n474), .B1(new_n497), .B2(new_n500), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n510), .B1(new_n692), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n647), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n647), .A2(new_n710), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n512), .A2(new_n514), .A3(new_n712), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n613), .B(KEYINPUT104), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n673), .B(KEYINPUT105), .Z(new_n716));
  AND3_X1   g515(.A1(new_n715), .A2(new_n588), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n714), .A2(new_n590), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G29gat), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n613), .A2(new_n647), .A3(new_n673), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n512), .A2(new_n514), .A3(new_n588), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n590), .A2(new_n531), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n721), .A2(KEYINPUT103), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT103), .B1(new_n721), .B2(new_n722), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(new_n723), .B2(new_n725), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n719), .B1(new_n726), .B2(new_n727), .ZN(G1328gat));
  NAND4_X1  g527(.A1(new_n711), .A2(new_n713), .A3(new_n443), .A4(new_n717), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n532), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n730), .B2(new_n729), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n443), .A2(new_n532), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT46), .B1(new_n721), .B2(new_n733), .ZN(new_n734));
  OR3_X1    g533(.A1(new_n721), .A2(KEYINPUT46), .A3(new_n733), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(G1329gat));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n711), .A2(new_n713), .A3(new_n692), .A4(new_n717), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n738), .A2(G43gat), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n695), .A2(G43gat), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n589), .A2(new_n740), .A3(new_n720), .A4(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n741), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT107), .B1(new_n721), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n737), .B1(new_n739), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n738), .A2(G43gat), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n747), .A2(KEYINPUT47), .A3(new_n744), .A4(new_n742), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(G1330gat));
  NAND4_X1  g548(.A1(new_n711), .A2(new_n713), .A3(new_n473), .A4(new_n717), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G50gat), .ZN(new_n751));
  OR3_X1    g550(.A1(new_n721), .A2(G50gat), .A3(new_n498), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT48), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n751), .A2(KEYINPUT48), .A3(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(G1331gat));
  INV_X1    g556(.A(new_n588), .ZN(new_n758));
  INV_X1    g557(.A(new_n716), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n652), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n707), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n590), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g563(.A1(new_n761), .A2(KEYINPUT108), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n707), .B2(new_n760), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n765), .A2(new_n444), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  AND2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n768), .B2(new_n769), .ZN(G1333gat));
  NAND2_X1  g571(.A1(new_n762), .A2(new_n766), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n774));
  INV_X1    g573(.A(new_n767), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n692), .A2(G71gat), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n773), .A2(new_n774), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n765), .A2(new_n767), .A3(new_n776), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n707), .A2(new_n502), .A3(new_n760), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT109), .B1(new_n780), .B2(new_n593), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n778), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT50), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n778), .B(new_n784), .C1(new_n779), .C2(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1334gat));
  NOR3_X1   g585(.A1(new_n765), .A2(new_n498), .A3(new_n767), .ZN(new_n787));
  XOR2_X1   g586(.A(KEYINPUT110), .B(G78gat), .Z(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1335gat));
  INV_X1    g588(.A(new_n613), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n758), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n674), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n711), .A2(new_n713), .A3(new_n590), .A4(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G85gat), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n793), .A2(new_n794), .ZN(new_n797));
  INV_X1    g596(.A(new_n791), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n707), .A2(new_n708), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n707), .A2(KEYINPUT51), .A3(new_n708), .A4(new_n798), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n590), .A2(new_n616), .A3(new_n673), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n796), .A2(new_n797), .B1(new_n804), .B2(new_n805), .ZN(G1336gat));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n801), .A2(new_n807), .A3(new_n802), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n799), .A2(KEYINPUT112), .A3(new_n800), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n716), .A2(G92gat), .A3(new_n444), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n711), .A2(new_n713), .A3(new_n443), .A4(new_n792), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G92gat), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT52), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT52), .B1(new_n803), .B2(new_n810), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(G1337gat));
  NAND3_X1  g617(.A1(new_n714), .A2(new_n692), .A3(new_n792), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(G99gat), .ZN(new_n820));
  OR3_X1    g619(.A1(new_n695), .A2(G99gat), .A3(new_n674), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n804), .B2(new_n821), .ZN(G1338gat));
  NOR3_X1   g621(.A1(new_n716), .A2(new_n498), .A3(G106gat), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT113), .Z(new_n824));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n711), .A2(new_n713), .A3(new_n473), .A4(new_n792), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G106gat), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT53), .B1(new_n803), .B2(new_n824), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n827), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(G1339gat));
  NAND2_X1  g631(.A1(new_n588), .A2(new_n271), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT118), .ZN(new_n834));
  INV_X1    g633(.A(new_n672), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n660), .A2(new_n654), .A3(new_n661), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n836), .A2(new_n662), .A3(new_n837), .ZN(new_n838));
  AOI211_X1 g637(.A(KEYINPUT54), .B(new_n654), .C1(new_n660), .C2(new_n661), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT114), .B1(new_n839), .B2(new_n669), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n662), .A2(new_n837), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n842), .A3(new_n670), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n838), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n835), .B1(new_n844), .B2(KEYINPUT55), .ZN(new_n845));
  INV_X1    g644(.A(new_n838), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n842), .B1(new_n841), .B2(new_n670), .ZN(new_n847));
  AOI211_X1 g646(.A(KEYINPUT114), .B(new_n669), .C1(new_n662), .C2(new_n837), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n845), .A2(new_n588), .A3(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n555), .A2(new_n556), .A3(new_n554), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n548), .B1(new_n547), .B2(new_n552), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n570), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n578), .A2(new_n673), .A3(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n708), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n578), .A2(new_n855), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n859), .A2(new_n845), .A3(new_n708), .A4(new_n851), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT115), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n583), .B1(new_n561), .B2(new_n558), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT91), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n584), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n866), .A2(new_n578), .B1(new_n849), .B2(new_n850), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n856), .B1(new_n867), .B2(new_n845), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n863), .B(new_n860), .C1(new_n868), .C2(new_n708), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n862), .A2(new_n869), .A3(new_n715), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n652), .A2(new_n758), .A3(new_n674), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n508), .A2(new_n394), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n443), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n872), .A2(KEYINPUT116), .A3(new_n873), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n876), .A2(KEYINPUT117), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT117), .B1(new_n876), .B2(new_n877), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n834), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n874), .A2(new_n443), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G113gat), .B1(new_n882), .B2(new_n758), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n883), .ZN(G1340gat));
  AOI21_X1  g683(.A(new_n273), .B1(new_n881), .B2(new_n759), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT119), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n273), .B(new_n673), .C1(new_n878), .C2(new_n879), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1341gat));
  NAND2_X1  g687(.A1(new_n277), .A2(new_n279), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n889), .B1(new_n882), .B2(new_n715), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n876), .A2(new_n877), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n613), .A2(new_n277), .A3(new_n279), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(G1342gat));
  NAND2_X1  g692(.A1(new_n708), .A2(new_n283), .ZN(new_n894));
  OR3_X1    g693(.A1(new_n891), .A2(KEYINPUT56), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G134gat), .B1(new_n882), .B2(new_n647), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT56), .B1(new_n891), .B2(new_n894), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G1343gat));
  AOI21_X1  g697(.A(new_n498), .B1(new_n870), .B2(new_n871), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n652), .A2(new_n758), .A3(new_n674), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n852), .A2(new_n857), .A3(KEYINPUT120), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n647), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT120), .B1(new_n852), .B2(new_n857), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n860), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n902), .B1(new_n906), .B2(new_n790), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT57), .B1(new_n907), .B2(new_n498), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n394), .A2(new_n443), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n692), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n901), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G141gat), .B1(new_n912), .B2(new_n758), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n899), .A2(new_n911), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n758), .A2(G141gat), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n914), .A2(new_n915), .B1(KEYINPUT121), .B2(KEYINPUT58), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT122), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n917), .B(new_n919), .ZN(G1344gat));
  NAND2_X1  g719(.A1(new_n334), .A2(new_n336), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n914), .A2(new_n922), .A3(new_n673), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n925), .B1(new_n692), .B2(new_n910), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n690), .A2(new_n691), .A3(KEYINPUT123), .A4(new_n909), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n673), .A3(new_n927), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n907), .A2(KEYINPUT57), .A3(new_n498), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n900), .B1(new_n872), .B2(new_n473), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n333), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n929), .A2(new_n930), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT124), .B1(new_n934), .B2(new_n928), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n924), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n912), .A2(new_n674), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(KEYINPUT59), .A3(new_n922), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n923), .B1(new_n936), .B2(new_n938), .ZN(G1345gat));
  OAI21_X1  g738(.A(G155gat), .B1(new_n912), .B2(new_n715), .ZN(new_n940));
  INV_X1    g739(.A(G155gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n914), .A2(new_n941), .A3(new_n613), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(G1346gat));
  OAI21_X1  g742(.A(G162gat), .B1(new_n912), .B2(new_n647), .ZN(new_n944));
  INV_X1    g743(.A(G162gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n914), .A2(new_n945), .A3(new_n708), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(G1347gat));
  NOR3_X1   g746(.A1(new_n508), .A2(new_n590), .A3(new_n444), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n872), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n949), .A2(new_n758), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(new_n237), .ZN(G1348gat));
  OAI21_X1  g750(.A(G176gat), .B1(new_n949), .B2(new_n716), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n673), .A2(new_n238), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n949), .B2(new_n953), .ZN(G1349gat));
  OAI21_X1  g753(.A(G183gat), .B1(new_n949), .B2(new_n715), .ZN(new_n955));
  NAND2_X1  g754(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n613), .A2(new_n252), .A3(new_n255), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n955), .B(new_n956), .C1(new_n949), .C2(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n959));
  XOR2_X1   g758(.A(new_n958), .B(new_n959), .Z(G1350gat));
  OAI22_X1  g759(.A1(new_n949), .A2(new_n647), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n961));
  NAND2_X1  g760(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n961), .B(new_n962), .ZN(G1351gat));
  NOR3_X1   g762(.A1(new_n692), .A2(new_n590), .A3(new_n444), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n964), .A2(new_n899), .ZN(new_n965));
  AOI21_X1  g764(.A(G197gat), .B1(new_n965), .B2(new_n588), .ZN(new_n966));
  INV_X1    g765(.A(new_n964), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n934), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n758), .A2(new_n403), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(G1352gat));
  INV_X1    g769(.A(G204gat), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n971), .B1(new_n968), .B2(new_n759), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n965), .A2(new_n971), .A3(new_n673), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT62), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n972), .A2(new_n974), .ZN(G1353gat));
  NAND3_X1  g774(.A1(new_n965), .A2(new_n400), .A3(new_n613), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n929), .A2(new_n930), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n977), .A2(new_n613), .A3(new_n964), .ZN(new_n978));
  AND2_X1   g777(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n979));
  OAI21_X1  g778(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n978), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n979), .B1(new_n978), .B2(new_n981), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n976), .B1(new_n982), .B2(new_n983), .ZN(G1354gat));
  NAND3_X1  g783(.A1(new_n965), .A2(new_n401), .A3(new_n708), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n934), .A2(new_n647), .A3(new_n967), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n985), .B1(new_n986), .B2(new_n401), .ZN(G1355gat));
endmodule


