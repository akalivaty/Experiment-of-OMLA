//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n826, new_n827, new_n828,
    new_n829, new_n831, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  INV_X1    g004(.A(G176gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n203), .B(new_n204), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT25), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT24), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G183gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n212), .B1(new_n217), .B2(G190gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n219));
  XOR2_X1   g018(.A(new_n219), .B(KEYINPUT65), .Z(new_n220));
  OAI21_X1  g019(.A(new_n209), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n222));
  INV_X1    g021(.A(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n213), .A2(new_n223), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n212), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n222), .B1(new_n207), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229));
  INV_X1    g028(.A(G120gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G113gat), .B(G120gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT71), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n236));
  INV_X1    g035(.A(new_n228), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n232), .A2(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT28), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT27), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT67), .B1(new_n213), .B2(KEYINPUT27), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT27), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(new_n244), .A3(G183gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n245), .A3(new_n223), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n240), .B1(new_n241), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(G183gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n213), .A2(KEYINPUT27), .ZN(new_n249));
  AND4_X1   g048(.A1(KEYINPUT28), .A2(new_n248), .A3(new_n249), .A4(new_n223), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n247), .A2(KEYINPUT68), .A3(new_n251), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n202), .A2(KEYINPUT69), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT26), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n257), .A2(new_n258), .B1(G169gat), .B2(G176gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n202), .A2(KEYINPUT69), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT26), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n262), .A2(new_n210), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n239), .B1(new_n256), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT27), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n265), .A2(new_n223), .A3(new_n245), .A4(new_n242), .ZN(new_n266));
  AOI211_X1 g065(.A(new_n253), .B(new_n250), .C1(new_n266), .C2(new_n240), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT68), .B1(new_n247), .B2(new_n251), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n263), .B(new_n239), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n227), .B(new_n238), .C1(new_n264), .C2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n227), .B1(new_n264), .B2(new_n270), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n232), .A2(new_n235), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n236), .A2(new_n237), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n227), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n263), .B1(new_n267), .B2(new_n268), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT70), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n279), .B1(new_n281), .B2(new_n269), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(KEYINPUT72), .A3(new_n238), .ZN(new_n283));
  NAND2_X1  g082(.A1(G227gat), .A2(G233gat), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n273), .A2(new_n278), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(KEYINPUT34), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT32), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n273), .A2(new_n283), .A3(new_n278), .ZN(new_n288));
  INV_X1    g087(.A(new_n284), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT33), .B1(new_n288), .B2(new_n289), .ZN(new_n291));
  XOR2_X1   g090(.A(G15gat), .B(G43gat), .Z(new_n292));
  XNOR2_X1  g091(.A(G71gat), .B(G99gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n290), .A2(new_n291), .A3(new_n295), .ZN(new_n296));
  AOI221_X4 g095(.A(new_n287), .B1(KEYINPUT33), .B2(new_n294), .C1(new_n288), .C2(new_n289), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n286), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n288), .A2(new_n289), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT33), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n295), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n290), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n285), .B(KEYINPUT34), .Z(new_n304));
  INV_X1    g103(.A(new_n297), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n298), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  OAI211_X1 g107(.A(KEYINPUT73), .B(new_n286), .C1(new_n296), .C2(new_n297), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(G226gat), .A2(G233gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT29), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n274), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT75), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT74), .B(G197gat), .Z(new_n316));
  INV_X1    g115(.A(G204gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT74), .B(G197gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G204gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(G211gat), .B(G218gat), .Z(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n325), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n321), .A2(new_n327), .A3(new_n323), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n280), .A2(new_n227), .A3(new_n312), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n314), .A2(new_n315), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n313), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n330), .B(new_n331), .C1(new_n282), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT75), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n282), .A2(new_n312), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n333), .B1(new_n280), .B2(new_n227), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n330), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n332), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT76), .ZN(new_n341));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n342), .B(new_n343), .Z(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n332), .B(new_n346), .C1(new_n335), .C2(new_n339), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n341), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n340), .A2(new_n344), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT30), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n340), .A2(KEYINPUT30), .A3(new_n344), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT35), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT31), .B(G50gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358));
  INV_X1    g157(.A(G141gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G148gat), .ZN(new_n360));
  INV_X1    g159(.A(G148gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G141gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n360), .A2(new_n362), .B1(KEYINPUT2), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n363), .ZN(new_n365));
  NOR2_X1   g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(KEYINPUT79), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n363), .A2(KEYINPUT78), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(G155gat), .B2(G162gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(G155gat), .A3(G162gat), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n368), .A2(new_n369), .A3(new_n371), .A4(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n367), .B1(new_n364), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n327), .B1(new_n321), .B2(new_n323), .ZN(new_n376));
  AOI211_X1 g175(.A(new_n325), .B(new_n322), .C1(new_n318), .C2(new_n320), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n358), .B(new_n375), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n375), .A2(KEYINPUT3), .ZN(new_n379));
  INV_X1    g178(.A(new_n375), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT29), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n378), .B(new_n379), .C1(new_n382), .C2(new_n329), .ZN(new_n383));
  NAND2_X1  g182(.A1(G228gat), .A2(G233gat), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n383), .A2(KEYINPUT85), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT85), .B1(new_n383), .B2(new_n384), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n382), .A2(new_n329), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n387), .A2(new_n384), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n358), .B1(new_n376), .B2(new_n377), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n390), .A2(KEYINPUT86), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT3), .B1(new_n390), .B2(KEYINPUT86), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n380), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI22_X1  g192(.A1(new_n385), .A2(new_n386), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G22gat), .ZN(new_n395));
  INV_X1    g194(.A(G22gat), .ZN(new_n396));
  OAI221_X1 g195(.A(new_n396), .B1(new_n389), .B2(new_n393), .C1(new_n385), .C2(new_n386), .ZN(new_n397));
  XNOR2_X1  g196(.A(G78gat), .B(G106gat), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n398), .B(KEYINPUT84), .Z(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n395), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n400), .B1(new_n395), .B2(new_n397), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n357), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n395), .A2(new_n397), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n399), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n395), .A2(new_n397), .A3(new_n400), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n356), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT6), .ZN(new_n409));
  OR2_X1    g208(.A1(new_n374), .A2(new_n364), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n410), .A2(new_n381), .A3(new_n367), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n379), .A2(new_n277), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n410), .A2(new_n275), .A3(new_n276), .A4(new_n367), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n238), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n412), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n418));
  NAND2_X1  g217(.A1(G225gat), .A2(G233gat), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n417), .A2(KEYINPUT82), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT82), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n412), .A2(new_n415), .A3(new_n416), .A4(new_n419), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(KEYINPUT5), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n277), .A2(new_n375), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n413), .ZN(new_n425));
  INV_X1    g224(.A(new_n419), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n418), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n420), .A2(new_n423), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G57gat), .B(G85gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT81), .ZN(new_n430));
  XOR2_X1   g229(.A(KEYINPUT80), .B(KEYINPUT0), .Z(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G1gat), .B(G29gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n409), .B1(new_n428), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n423), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n427), .A2(new_n422), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n437), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT89), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n438), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n434), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n428), .A2(new_n435), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT89), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .A4(new_n409), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(KEYINPUT6), .A3(new_n434), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n440), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n354), .A2(new_n355), .A3(new_n408), .A4(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n311), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT77), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n348), .A2(new_n450), .A3(new_n352), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n442), .A2(new_n409), .A3(new_n443), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n349), .A2(new_n350), .B1(new_n452), .B2(new_n446), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n450), .B1(new_n348), .B2(new_n352), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT83), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n348), .A2(new_n352), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT77), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT83), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n458), .A2(new_n459), .A3(new_n451), .A4(new_n453), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n408), .A2(new_n298), .A3(new_n306), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n456), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT93), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n449), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(KEYINPUT93), .A3(KEYINPUT35), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT92), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT37), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n344), .B1(new_n340), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n314), .A2(new_n329), .A3(new_n331), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT37), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n329), .B1(new_n336), .B2(new_n338), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT90), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n472), .A2(KEYINPUT90), .A3(new_n473), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n468), .B(new_n470), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  AND4_X1   g277(.A1(new_n349), .A2(new_n440), .A3(new_n446), .A4(new_n445), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n341), .A2(KEYINPUT37), .A3(new_n347), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n468), .B1(new_n481), .B2(new_n470), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n408), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n417), .A2(new_n419), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n484), .A2(KEYINPUT39), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n485), .A2(new_n434), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n425), .B2(new_n426), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n424), .A2(KEYINPUT87), .A3(new_n413), .A4(new_n419), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(KEYINPUT39), .A3(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n490), .A2(KEYINPUT88), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(KEYINPUT88), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n484), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n486), .A2(new_n493), .A3(KEYINPUT40), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n486), .A2(new_n493), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n442), .A2(KEYINPUT40), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n353), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n467), .B1(new_n483), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n481), .A2(new_n470), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n478), .B(new_n479), .C1(new_n501), .C2(new_n468), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n502), .A2(KEYINPUT92), .A3(new_n498), .A4(new_n408), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n310), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n298), .A2(new_n306), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT36), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n408), .B1(new_n456), .B2(new_n460), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n465), .A2(new_n466), .B1(new_n504), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT18), .ZN(new_n513));
  INV_X1    g312(.A(G36gat), .ZN(new_n514));
  AND2_X1   g313(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(G29gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n522));
  XNOR2_X1  g321(.A(G43gat), .B(G50gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(new_n522), .B2(new_n523), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT17), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n527), .A2(G1gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT95), .ZN(new_n529));
  AOI21_X1  g328(.A(G8gat), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT16), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n527), .B1(new_n531), .B2(G1gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n530), .B(new_n533), .Z(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n526), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n525), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n513), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n536), .A2(KEYINPUT18), .A3(new_n539), .A4(new_n537), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT96), .B1(new_n534), .B2(new_n525), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(new_n537), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n539), .B(KEYINPUT13), .Z(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G113gat), .B(G141gat), .Z(new_n547));
  XNOR2_X1  g346(.A(G169gat), .B(G197gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT94), .B(KEYINPUT11), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n549), .B(new_n550), .Z(new_n551));
  XOR2_X1   g350(.A(new_n551), .B(KEYINPUT12), .Z(new_n552));
  NAND4_X1  g351(.A1(new_n541), .A2(new_n542), .A3(new_n546), .A4(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT97), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(KEYINPUT97), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n546), .ZN(new_n558));
  INV_X1    g357(.A(new_n552), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G57gat), .B(G64gat), .Z(new_n563));
  NAND2_X1  g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT9), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G71gat), .ZN(new_n567));
  INV_X1    g366(.A(G78gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(new_n564), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n563), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n571), .B(KEYINPUT99), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n569), .B(KEYINPUT98), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n563), .A2(new_n566), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(new_n574), .A3(new_n564), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT100), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G85gat), .ZN(new_n579));
  INV_X1    g378(.A(G92gat), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT101), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT101), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(G85gat), .A3(G92gat), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n583), .A3(KEYINPUT7), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT8), .A2(new_n585), .B1(new_n579), .B2(new_n580), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n584), .B(new_n586), .C1(KEYINPUT7), .C2(new_n581), .ZN(new_n587));
  XNOR2_X1  g386(.A(G99gat), .B(G106gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n587), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT102), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n578), .A2(KEYINPUT10), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n576), .B(new_n590), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n592), .B1(KEYINPUT10), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G230gat), .A2(G233gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n595), .B(KEYINPUT104), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n593), .A2(new_n596), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G120gat), .B(G148gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(G176gat), .B(G204gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT105), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT106), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n606), .B1(new_n604), .B2(new_n605), .ZN(new_n609));
  OAI22_X1  g408(.A1(new_n608), .A2(new_n609), .B1(new_n600), .B2(new_n603), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n604), .A2(new_n605), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT106), .ZN(new_n612));
  INV_X1    g411(.A(new_n600), .ZN(new_n613));
  INV_X1    g412(.A(new_n603), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .A4(new_n607), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT21), .B1(new_n572), .B2(new_n575), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G127gat), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n534), .B1(new_n578), .B2(KEYINPUT21), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G155gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G183gat), .B(G211gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(new_n626), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n591), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n630), .A2(new_n526), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n591), .A2(new_n525), .ZN(new_n632));
  XNOR2_X1  g431(.A(G190gat), .B(G218gat), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT103), .ZN(new_n634));
  AND2_X1   g433(.A1(G232gat), .A2(G233gat), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n633), .A2(new_n634), .B1(KEYINPUT41), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n633), .A2(new_n634), .ZN(new_n638));
  OR3_X1    g437(.A1(new_n631), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n635), .A2(KEYINPUT41), .ZN(new_n640));
  XNOR2_X1  g439(.A(G134gat), .B(G162gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n638), .B1(new_n631), .B2(new_n637), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n639), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n642), .B1(new_n639), .B2(new_n643), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n629), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n616), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n512), .A2(new_n562), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n452), .A2(new_n446), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(KEYINPUT107), .Z(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT108), .B(G1gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1324gat));
  NOR2_X1   g454(.A1(new_n512), .A2(new_n562), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(new_n353), .A3(new_n648), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n657), .A2(G8gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT16), .B(G8gat), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT42), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(KEYINPUT42), .B2(new_n660), .ZN(G1325gat));
  AOI21_X1  g461(.A(G15gat), .B1(new_n650), .B2(new_n310), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n509), .A2(G15gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT109), .Z(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n650), .B2(new_n665), .ZN(G1326gat));
  INV_X1    g465(.A(new_n408), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT43), .B(G22gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  AND4_X1   g469(.A1(new_n656), .A2(new_n629), .A3(new_n646), .A4(new_n616), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(new_n518), .A3(new_n652), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  INV_X1    g474(.A(new_n646), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n675), .B1(new_n512), .B2(new_n676), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n462), .A2(KEYINPUT93), .A3(KEYINPUT35), .ZN(new_n678));
  AOI21_X1  g477(.A(KEYINPUT93), .B1(new_n462), .B2(KEYINPUT35), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n678), .A2(new_n679), .A3(new_n449), .ZN(new_n680));
  INV_X1    g479(.A(new_n509), .ZN(new_n681));
  INV_X1    g480(.A(new_n510), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n681), .A2(new_n504), .A3(new_n682), .ZN(new_n683));
  OAI211_X1 g482(.A(KEYINPUT44), .B(new_n646), .C1(new_n680), .C2(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n616), .A2(new_n561), .A3(new_n629), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n652), .ZN(new_n689));
  OAI21_X1  g488(.A(G29gat), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n690), .ZN(G1328gat));
  NAND3_X1  g490(.A1(new_n671), .A2(new_n514), .A3(new_n353), .ZN(new_n692));
  AND2_X1   g491(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n693));
  NOR2_X1   g492(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(G36gat), .B1(new_n688), .B2(new_n354), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n695), .B(new_n696), .C1(new_n693), .C2(new_n692), .ZN(G1329gat));
  INV_X1    g496(.A(G43gat), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n671), .A2(new_n698), .A3(new_n310), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n677), .A2(new_n509), .A3(new_n684), .A4(new_n687), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(G43gat), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1330gat));
  INV_X1    g503(.A(G50gat), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n671), .A2(new_n705), .A3(new_n667), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n677), .A2(new_n667), .A3(new_n684), .A4(new_n687), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G50gat), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT48), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1331gat));
  NAND2_X1  g510(.A1(new_n465), .A2(new_n466), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n511), .A2(new_n504), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR4_X1   g513(.A1(new_n616), .A2(new_n561), .A3(new_n629), .A4(new_n646), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n652), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g518(.A1(new_n716), .A2(new_n354), .ZN(new_n720));
  NOR2_X1   g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  AND2_X1   g520(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n720), .B2(new_n721), .ZN(G1333gat));
  OAI21_X1  g523(.A(G71gat), .B1(new_n716), .B2(new_n681), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n310), .A2(new_n567), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n716), .B2(new_n726), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g527(.A1(new_n716), .A2(new_n408), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(new_n568), .ZN(G1335gat));
  INV_X1    g529(.A(new_n629), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n561), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n646), .B(new_n732), .C1(new_n680), .C2(new_n683), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n616), .B1(new_n733), .B2(KEYINPUT51), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n714), .A2(new_n735), .A3(new_n646), .A4(new_n732), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n734), .A2(new_n579), .A3(new_n652), .A4(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n616), .A2(new_n731), .A3(new_n561), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n685), .A2(new_n652), .A3(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT112), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G85gat), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n739), .A2(new_n740), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n737), .B1(new_n742), .B2(new_n743), .ZN(G1336gat));
  NAND4_X1  g543(.A1(new_n677), .A2(new_n353), .A3(new_n684), .A4(new_n738), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G92gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n733), .A2(KEYINPUT51), .ZN(new_n747));
  INV_X1    g546(.A(new_n616), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n354), .A2(G92gat), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n747), .A2(new_n748), .A3(new_n736), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT52), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n750), .A2(KEYINPUT114), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n734), .A2(new_n758), .A3(new_n736), .A4(new_n749), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n756), .A2(new_n757), .A3(new_n746), .A4(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n754), .A2(new_n755), .A3(new_n760), .ZN(G1337gat));
  NAND4_X1  g560(.A1(new_n747), .A2(new_n310), .A3(new_n736), .A4(new_n748), .ZN(new_n762));
  INV_X1    g561(.A(G99gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n685), .A2(new_n738), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n509), .A2(G99gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n764), .B(KEYINPUT115), .C1(new_n765), .C2(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1338gat));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n408), .A2(G106gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n734), .A2(new_n736), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n772), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n677), .A2(new_n667), .A3(new_n684), .A4(new_n738), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G106gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n774), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n776), .B(new_n779), .ZN(G1339gat));
  NAND2_X1  g579(.A1(new_n648), .A2(new_n562), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n598), .A2(KEYINPUT54), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(new_n603), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n594), .B2(new_n597), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n592), .B(new_n596), .C1(KEYINPUT10), .C2(new_n593), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n785), .A2(KEYINPUT117), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT117), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n783), .B(KEYINPUT55), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(KEYINPUT118), .A3(new_n604), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT118), .B1(new_n789), .B2(new_n604), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n544), .A2(new_n545), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n540), .B2(new_n538), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n797), .A2(new_n551), .ZN(new_n798));
  INV_X1    g597(.A(new_n556), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n646), .B(new_n798), .C1(new_n799), .C2(new_n554), .ZN(new_n800));
  NOR4_X1   g599(.A1(new_n791), .A2(new_n792), .A3(new_n795), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n789), .A2(new_n604), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n793), .A2(new_n794), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n804), .A2(new_n561), .A3(new_n790), .A4(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n557), .A2(new_n798), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n610), .A2(new_n615), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n801), .B1(new_n809), .B2(new_n676), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n781), .B1(new_n810), .B2(new_n731), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n811), .A2(new_n408), .A3(new_n310), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n689), .A2(new_n353), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G113gat), .B1(new_n814), .B2(new_n562), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n811), .A2(new_n652), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n507), .A2(new_n667), .A3(new_n353), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n562), .A2(G113gat), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT119), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n815), .B1(new_n818), .B2(new_n820), .ZN(G1340gat));
  INV_X1    g620(.A(new_n818), .ZN(new_n822));
  AOI21_X1  g621(.A(G120gat), .B1(new_n822), .B2(new_n748), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n814), .A2(new_n230), .A3(new_n616), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(G1341gat));
  NAND4_X1  g624(.A1(new_n812), .A2(G127gat), .A3(new_n731), .A4(new_n813), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(KEYINPUT120), .ZN(new_n827));
  AOI21_X1  g626(.A(G127gat), .B1(new_n822), .B2(new_n731), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n826), .A2(KEYINPUT120), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(G1342gat));
  OR3_X1    g629(.A1(new_n818), .A2(G134gat), .A3(new_n676), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n831), .A2(KEYINPUT56), .ZN(new_n832));
  OAI21_X1  g631(.A(G134gat), .B1(new_n814), .B2(new_n676), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n831), .A2(KEYINPUT121), .A3(KEYINPUT56), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT121), .B1(new_n831), .B2(KEYINPUT56), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n832), .B(new_n833), .C1(new_n834), .C2(new_n835), .ZN(G1343gat));
  NOR3_X1   g635(.A1(new_n509), .A2(new_n353), .A3(new_n408), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n816), .A2(new_n837), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(G141gat), .A3(new_n562), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n509), .A2(new_n353), .A3(new_n689), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT57), .B1(new_n811), .B2(new_n667), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n667), .A2(KEYINPUT57), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n561), .A2(new_n604), .A3(new_n805), .A4(new_n789), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n646), .B1(new_n808), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n629), .B1(new_n845), .B2(new_n801), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n843), .B1(new_n846), .B2(new_n781), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n841), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G141gat), .B1(new_n848), .B2(new_n562), .ZN(new_n849));
  XNOR2_X1  g648(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n840), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g652(.A(KEYINPUT122), .B(new_n841), .C1(new_n842), .C2(new_n847), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n561), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n839), .B1(new_n855), .B2(G141gat), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n851), .B1(new_n856), .B2(new_n857), .ZN(G1344gat));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  INV_X1    g658(.A(new_n838), .ZN(new_n860));
  AOI211_X1 g659(.A(new_n859), .B(G148gat), .C1(new_n860), .C2(new_n748), .ZN(new_n861));
  INV_X1    g660(.A(new_n843), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n811), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n781), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT57), .B1(new_n864), .B2(new_n667), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n748), .A3(new_n841), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n361), .B1(new_n867), .B2(KEYINPUT59), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n853), .A2(new_n859), .A3(new_n748), .A4(new_n854), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n861), .B1(new_n868), .B2(new_n869), .ZN(G1345gat));
  INV_X1    g669(.A(G155gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n860), .A2(new_n871), .A3(new_n731), .ZN(new_n872));
  INV_X1    g671(.A(new_n853), .ZN(new_n873));
  INV_X1    g672(.A(new_n854), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n873), .A2(new_n874), .A3(new_n629), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n872), .B1(new_n875), .B2(new_n871), .ZN(G1346gat));
  NOR3_X1   g675(.A1(new_n838), .A2(G162gat), .A3(new_n676), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT124), .ZN(new_n878));
  INV_X1    g677(.A(G162gat), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n873), .A2(new_n874), .A3(new_n676), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(G1347gat));
  NOR2_X1   g680(.A1(new_n652), .A2(new_n354), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n812), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(new_n205), .A3(new_n562), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n811), .A2(new_n461), .A3(new_n882), .ZN(new_n885));
  AOI21_X1  g684(.A(G169gat), .B1(new_n885), .B2(new_n561), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n884), .A2(new_n886), .ZN(G1348gat));
  OAI21_X1  g686(.A(G176gat), .B1(new_n883), .B2(new_n616), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n885), .A2(new_n206), .A3(new_n748), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1349gat));
  NAND3_X1  g689(.A1(new_n812), .A2(new_n731), .A3(new_n882), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n731), .A2(new_n248), .A3(new_n249), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n891), .A2(new_n217), .B1(new_n885), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n894), .A2(KEYINPUT60), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n893), .A2(KEYINPUT126), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(KEYINPUT126), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT60), .B1(new_n893), .B2(new_n894), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(G1350gat));
  OAI21_X1  g698(.A(G190gat), .B1(new_n883), .B2(new_n676), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT61), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n885), .A2(new_n223), .A3(new_n646), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1351gat));
  AND2_X1   g702(.A1(new_n811), .A2(new_n667), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n509), .A2(new_n354), .A3(new_n652), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(G197gat), .B1(new_n907), .B2(new_n561), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n905), .B1(new_n863), .B2(new_n865), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n561), .A2(G197gat), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1352gat));
  NOR3_X1   g711(.A1(new_n906), .A2(G204gat), .A3(new_n616), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT62), .ZN(new_n914));
  OAI21_X1  g713(.A(G204gat), .B1(new_n909), .B2(new_n616), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1353gat));
  OR3_X1    g715(.A1(new_n906), .A2(G211gat), .A3(new_n629), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n910), .A2(new_n731), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT63), .B1(new_n918), .B2(G211gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(G1354gat));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n676), .B1(new_n909), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n923), .B1(new_n922), .B2(new_n909), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G218gat), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n676), .A2(G218gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n906), .B2(new_n926), .ZN(G1355gat));
endmodule


