//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G141gat), .ZN(new_n203));
  INV_X1    g002(.A(G148gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT74), .ZN(new_n208));
  OR2_X1    g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(KEYINPUT2), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT74), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n205), .A2(new_n213), .A3(new_n206), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n208), .A2(new_n211), .A3(new_n212), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n211), .A2(KEYINPUT73), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n212), .A2(new_n205), .A3(new_n206), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT73), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n209), .A2(new_n218), .A3(new_n210), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n222));
  XNOR2_X1  g021(.A(G113gat), .B(G120gat), .ZN(new_n223));
  OR2_X1    g022(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G127gat), .B(G134gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n226), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(new_n223), .B2(new_n224), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n220), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n222), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n221), .A2(new_n230), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT76), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT76), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(new_n221), .B2(new_n230), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT4), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n202), .B(new_n233), .C1(new_n238), .C2(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT77), .B(KEYINPUT5), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n221), .A2(new_n230), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n235), .A2(new_n237), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n202), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n242), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G1gat), .B(G29gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT0), .ZN(new_n249));
  XNOR2_X1  g048(.A(G57gat), .B(G85gat), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n249), .B(new_n250), .Z(new_n251));
  INV_X1    g050(.A(new_n233), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n235), .A2(KEYINPUT4), .A3(new_n237), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n239), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n242), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(new_n245), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n247), .A2(new_n251), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT78), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n247), .A2(new_n258), .ZN(new_n261));
  INV_X1    g060(.A(new_n251), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT6), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT78), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n247), .A2(new_n265), .A3(new_n251), .A4(new_n258), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n260), .A2(new_n263), .A3(new_n264), .A4(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n261), .A2(KEYINPUT6), .A3(new_n262), .ZN(new_n268));
  NAND2_X1  g067(.A1(G226gat), .A2(G233gat), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT23), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  OR2_X1    g072(.A1(G183gat), .A2(G190gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(KEYINPUT24), .A3(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n275), .A2(KEYINPUT24), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT64), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT25), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n278), .A2(new_n279), .B1(G169gat), .B2(G176gat), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n273), .A2(new_n276), .A3(new_n277), .A4(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n278), .A2(new_n279), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n277), .A2(new_n280), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n285), .A2(new_n282), .A3(new_n273), .A4(new_n276), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT27), .B(G183gat), .ZN(new_n288));
  INV_X1    g087(.A(G190gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n275), .ZN(new_n293));
  NOR3_X1   g092(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT65), .ZN(new_n295));
  INV_X1    g094(.A(G169gat), .ZN(new_n296));
  INV_X1    g095(.A(G176gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n271), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(KEYINPUT26), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n293), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n270), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n284), .A2(new_n286), .B1(new_n292), .B2(new_n301), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(new_n269), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT69), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT22), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n310), .A2(new_n311), .B1(G211gat), .B2(G218gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(KEYINPUT69), .A2(KEYINPUT22), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G204gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G197gat), .ZN(new_n316));
  INV_X1    g115(.A(G197gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G204gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT68), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n319), .B1(new_n316), .B2(new_n318), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n314), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(KEYINPUT70), .B(new_n314), .C1(new_n320), .C2(new_n321), .ZN(new_n325));
  XNOR2_X1  g124(.A(G211gat), .B(G218gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  AND4_X1   g126(.A1(new_n309), .A2(new_n324), .A3(new_n325), .A4(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n314), .B(new_n326), .C1(new_n320), .C2(new_n321), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT71), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n326), .B1(new_n322), .B2(new_n323), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n330), .B1(new_n331), .B2(new_n325), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n308), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n333), .ZN(new_n335));
  XOR2_X1   g134(.A(KEYINPUT72), .B(KEYINPUT29), .Z(new_n336));
  AOI21_X1  g135(.A(new_n270), .B1(new_n303), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n335), .B1(new_n337), .B2(new_n307), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G8gat), .B(G36gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  OR3_X1    g142(.A1(new_n339), .A2(KEYINPUT30), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n339), .A2(new_n343), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n334), .A2(new_n338), .A3(new_n342), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(KEYINPUT30), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n267), .A2(new_n268), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n317), .A2(G204gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n315), .A2(G197gat), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT68), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n352), .A2(new_n353), .B1(new_n313), .B2(new_n312), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n309), .B1(new_n354), .B2(new_n326), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n327), .B1(new_n354), .B2(KEYINPUT70), .ZN(new_n356));
  INV_X1    g155(.A(new_n325), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n331), .A2(new_n309), .A3(new_n325), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n358), .A2(new_n359), .B1(new_n232), .B2(new_n336), .ZN(new_n360));
  INV_X1    g159(.A(G228gat), .ZN(new_n361));
  INV_X1    g160(.A(G233gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n221), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n358), .A2(new_n304), .A3(new_n359), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n366), .B1(new_n367), .B2(new_n231), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI211_X1 g169(.A(KEYINPUT80), .B(new_n366), .C1(new_n367), .C2(new_n231), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n232), .A2(new_n336), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n372), .B1(new_n328), .B2(new_n332), .ZN(new_n373));
  INV_X1    g172(.A(new_n336), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n322), .A2(new_n327), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n374), .B1(new_n375), .B2(new_n329), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n221), .B1(new_n376), .B2(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT79), .B1(new_n378), .B2(new_n364), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT79), .ZN(new_n380));
  AOI211_X1 g179(.A(new_n380), .B(new_n363), .C1(new_n373), .C2(new_n377), .ZN(new_n381));
  OAI22_X1  g180(.A1(new_n370), .A2(new_n371), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(G22gat), .ZN(new_n383));
  INV_X1    g182(.A(G22gat), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT3), .B1(new_n333), .B2(new_n304), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT80), .B1(new_n385), .B2(new_n366), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n369), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n387), .A3(new_n365), .ZN(new_n388));
  INV_X1    g187(.A(new_n377), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n364), .B1(new_n360), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n380), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n378), .A2(KEYINPUT79), .A3(new_n364), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n384), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT81), .B1(new_n383), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT31), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(G50gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n382), .A2(G22gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n388), .A2(new_n384), .A3(new_n393), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT82), .ZN(new_n405));
  OAI211_X1 g204(.A(KEYINPUT81), .B(new_n398), .C1(new_n383), .C2(new_n394), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n404), .B2(new_n406), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n349), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n404), .A2(new_n406), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OR3_X1    g210(.A1(new_n255), .A2(KEYINPUT39), .A3(new_n202), .ZN(new_n412));
  OR2_X1    g211(.A1(new_n244), .A2(new_n245), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n413), .B(KEYINPUT39), .C1(new_n255), .C2(new_n202), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n414), .A3(new_n251), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT40), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n347), .A2(new_n344), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n415), .A2(new_n416), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT84), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n261), .A2(new_n423), .A3(new_n262), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n241), .A2(new_n246), .B1(new_n255), .B2(new_n257), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT84), .B1(new_n425), .B2(new_n251), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n419), .A2(new_n421), .A3(new_n422), .A4(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n268), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n266), .A2(new_n264), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n265), .B1(new_n425), .B2(new_n251), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n429), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n339), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT37), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n342), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n436), .B1(new_n435), .B2(new_n434), .ZN(new_n437));
  XOR2_X1   g236(.A(KEYINPUT85), .B(KEYINPUT38), .Z(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n435), .B1(new_n308), .B2(new_n335), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n333), .B1(new_n337), .B2(new_n307), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n438), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n433), .A2(new_n346), .A3(new_n439), .A4(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n411), .A2(new_n428), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT36), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n303), .A2(new_n230), .ZN(new_n447));
  INV_X1    g246(.A(new_n230), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n306), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(G227gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(new_n362), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT34), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT34), .ZN(new_n454));
  INV_X1    g253(.A(new_n452), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n447), .A2(new_n449), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(G15gat), .B(G43gat), .Z(new_n458));
  XNOR2_X1  g257(.A(G71gat), .B(G99gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n455), .B1(new_n447), .B2(new_n449), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n460), .B1(new_n461), .B2(KEYINPUT33), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT32), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI221_X4 g264(.A(new_n463), .B1(KEYINPUT33), .B2(new_n460), .C1(new_n450), .C2(new_n452), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n457), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n303), .A2(new_n230), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n306), .A2(new_n448), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n452), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT32), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT33), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n473), .A3(new_n460), .ZN(new_n474));
  INV_X1    g273(.A(new_n457), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n462), .A2(new_n464), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n467), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT67), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n474), .B2(new_n476), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  AOI211_X1 g281(.A(new_n479), .B(new_n457), .C1(new_n474), .C2(new_n476), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n446), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n478), .A2(KEYINPUT36), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n409), .A2(new_n445), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n483), .B1(new_n478), .B2(new_n481), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n404), .A2(new_n348), .A3(new_n406), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT35), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT35), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n420), .A2(new_n467), .A3(new_n492), .A4(new_n477), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n433), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(new_n406), .A3(new_n404), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n488), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G190gat), .B(G218gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(G29gat), .A2(G36gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(G43gat), .B(G50gat), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n501), .A2(KEYINPUT15), .ZN(new_n502));
  NOR2_X1   g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(KEYINPUT14), .ZN(new_n504));
  AOI211_X1 g303(.A(new_n500), .B(new_n502), .C1(KEYINPUT87), .C2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(KEYINPUT87), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT86), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G43gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(G50gat), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT15), .B1(new_n510), .B2(KEYINPUT86), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n506), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n502), .B1(new_n504), .B2(new_n500), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n513), .A2(KEYINPUT17), .A3(new_n514), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT7), .ZN(new_n519));
  INV_X1    g318(.A(G85gat), .ZN(new_n520));
  OAI21_X1  g319(.A(G92gat), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G92gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n522), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n521), .A2(new_n523), .B1(new_n519), .B2(new_n520), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT8), .ZN(new_n525));
  NAND2_X1  g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT93), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(new_n527), .B2(new_n526), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(G99gat), .B(G106gat), .Z(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n518), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(new_n513), .B2(new_n514), .ZN(new_n534));
  AND3_X1   g333(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n499), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n499), .A3(new_n536), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT94), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT94), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n533), .A2(new_n540), .A3(new_n536), .A4(new_n499), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT95), .B1(new_n539), .B2(new_n541), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G134gat), .B(G162gat), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n543), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n548), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n542), .B1(new_n544), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(G57gat), .B(G64gat), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G71gat), .B(G78gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n532), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n532), .A2(new_n558), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n553), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(KEYINPUT96), .Z(new_n562));
  INV_X1    g361(.A(new_n553), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT10), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n559), .A2(new_n564), .A3(new_n560), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G120gat), .B(G148gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(G176gat), .B(G204gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n572), .B(new_n573), .Z(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n562), .A2(new_n574), .A3(new_n568), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G15gat), .B(G22gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT16), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(G1gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT88), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n582), .B(new_n583), .C1(G1gat), .C2(new_n580), .ZN(new_n584));
  INV_X1    g383(.A(G8gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT21), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n586), .B1(new_n587), .B2(new_n558), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT92), .ZN(new_n589));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT91), .ZN(new_n591));
  XOR2_X1   g390(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n589), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n558), .A2(new_n587), .ZN(new_n595));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G183gat), .B(G211gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n552), .A2(new_n579), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n586), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n515), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G229gat), .A2(G233gat), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n606), .B(KEYINPUT13), .Z(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(KEYINPUT89), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n515), .A2(new_n604), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n586), .B1(new_n514), .B2(new_n513), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT89), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n517), .A2(new_n586), .A3(new_n518), .ZN(new_n615));
  INV_X1    g414(.A(new_n610), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n606), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT18), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G113gat), .B(G141gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G197gat), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT11), .B(G169gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n615), .A2(KEYINPUT18), .A3(new_n606), .A4(new_n616), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n614), .A2(new_n619), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT90), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n608), .A2(new_n613), .B1(new_n617), .B2(new_n618), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n630), .A2(KEYINPUT90), .A3(new_n625), .A4(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n626), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n629), .A2(new_n631), .B1(new_n632), .B2(new_n624), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n603), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n497), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n267), .A2(new_n268), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g439(.A(new_n585), .B1(new_n636), .B2(new_n421), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT16), .B(G8gat), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n635), .A2(new_n420), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT42), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n644), .B1(KEYINPUT42), .B2(new_n643), .ZN(G1325gat));
  INV_X1    g444(.A(new_n478), .ZN(new_n646));
  AOI21_X1  g445(.A(G15gat), .B1(new_n636), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT99), .B1(new_n485), .B2(new_n486), .ZN(new_n648));
  INV_X1    g447(.A(new_n486), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n649), .B(new_n650), .C1(new_n489), .C2(new_n446), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(G15gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n654), .B(KEYINPUT100), .Z(new_n655));
  AOI21_X1  g454(.A(new_n647), .B1(new_n636), .B2(new_n655), .ZN(G1326gat));
  NOR2_X1   g455(.A1(new_n407), .A2(new_n408), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n635), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT43), .B(G22gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  AOI21_X1  g459(.A(new_n552), .B1(new_n488), .B2(new_n496), .ZN(new_n661));
  INV_X1    g460(.A(G29gat), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n633), .A2(new_n602), .A3(new_n578), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n638), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT45), .ZN(new_n665));
  INV_X1    g464(.A(new_n663), .ZN(new_n666));
  INV_X1    g465(.A(new_n552), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n497), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT44), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n409), .A2(new_n445), .A3(new_n652), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n496), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n491), .A2(new_n495), .A3(KEYINPUT101), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n552), .A2(KEYINPUT44), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n666), .B1(new_n669), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n677), .A2(new_n638), .ZN(new_n678));
  OAI211_X1 g477(.A(KEYINPUT102), .B(new_n665), .C1(new_n678), .C2(new_n662), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT102), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n662), .B1(new_n677), .B2(new_n638), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n664), .B(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n680), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n679), .A2(new_n684), .ZN(G1328gat));
  NAND2_X1  g484(.A1(new_n677), .A2(new_n421), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n677), .A2(KEYINPUT104), .A3(new_n421), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(G36gat), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691));
  AOI21_X1  g490(.A(G36gat), .B1(new_n691), .B2(KEYINPUT46), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n661), .A2(new_n421), .A3(new_n663), .A4(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n691), .A2(KEYINPUT46), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n690), .A2(new_n695), .ZN(G1329gat));
  AND2_X1   g495(.A1(new_n674), .A2(new_n675), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n497), .B2(new_n667), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n653), .B(new_n663), .C1(new_n697), .C2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n676), .B1(new_n698), .B2(new_n661), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n703), .A2(KEYINPUT105), .A3(new_n653), .A4(new_n663), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(G43gat), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n661), .A2(new_n663), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n706), .A2(G43gat), .A3(new_n478), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n509), .B1(new_n677), .B2(new_n653), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n708), .B1(new_n711), .B2(new_n707), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(G1330gat));
  NOR3_X1   g512(.A1(new_n706), .A2(G50gat), .A3(new_n657), .ZN(new_n714));
  INV_X1    g513(.A(new_n657), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n677), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n714), .B1(new_n716), .B2(G50gat), .ZN(new_n717));
  INV_X1    g516(.A(G50gat), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n677), .B2(new_n410), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  OAI22_X1  g520(.A1(new_n717), .A2(KEYINPUT48), .B1(new_n719), .B2(new_n721), .ZN(G1331gat));
  INV_X1    g521(.A(new_n633), .ZN(new_n723));
  INV_X1    g522(.A(new_n602), .ZN(new_n724));
  NOR4_X1   g523(.A1(new_n667), .A2(new_n723), .A3(new_n724), .A4(new_n579), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n674), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n637), .B(KEYINPUT106), .Z(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n729), .B(G57gat), .Z(G1332gat));
  NAND2_X1  g529(.A1(new_n726), .A2(KEYINPUT107), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n674), .A2(new_n732), .A3(new_n725), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n420), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  AND2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n735), .B2(new_n736), .ZN(G1333gat));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741));
  INV_X1    g540(.A(G71gat), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n652), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n731), .A2(new_n741), .A3(new_n733), .A4(new_n743), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n731), .A2(new_n733), .A3(new_n743), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(new_n726), .B2(new_n478), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT108), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n740), .B(new_n744), .C1(new_n745), .C2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n731), .A2(new_n733), .A3(new_n743), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(KEYINPUT108), .A3(new_n746), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n740), .B1(new_n751), .B2(new_n744), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n749), .A2(new_n752), .ZN(G1334gat));
  NOR2_X1   g552(.A1(new_n734), .A2(new_n657), .ZN(new_n754));
  XOR2_X1   g553(.A(KEYINPUT109), .B(G78gat), .Z(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1335gat));
  NOR3_X1   g555(.A1(new_n723), .A2(new_n552), .A3(new_n602), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n674), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT51), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n579), .A2(G85gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n638), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n723), .A2(new_n602), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n578), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n669), .B2(new_n676), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n520), .B1(new_n765), .B2(new_n638), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT110), .B1(new_n762), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n703), .A2(new_n578), .A3(new_n763), .ZN(new_n768));
  OAI21_X1  g567(.A(G85gat), .B1(new_n768), .B2(new_n637), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n758), .B(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(new_n638), .A3(new_n760), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n769), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n767), .A2(new_n774), .ZN(G1336gat));
  NOR2_X1   g574(.A1(new_n579), .A2(G92gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n421), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n759), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n522), .B1(new_n765), .B2(new_n421), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT52), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(G92gat), .B1(new_n768), .B2(new_n420), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n772), .A2(new_n421), .A3(new_n776), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n780), .A2(new_n784), .ZN(G1337gat));
  OAI21_X1  g584(.A(G99gat), .B1(new_n768), .B2(new_n652), .ZN(new_n786));
  OR3_X1    g585(.A1(new_n579), .A2(G99gat), .A3(new_n478), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n759), .B2(new_n787), .ZN(G1338gat));
  NAND2_X1  g587(.A1(new_n765), .A2(new_n715), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n411), .A2(G106gat), .A3(new_n579), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n789), .A2(G106gat), .B1(new_n772), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  INV_X1    g591(.A(G106gat), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n765), .B2(new_n410), .ZN(new_n794));
  XOR2_X1   g593(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n795));
  INV_X1    g594(.A(new_n790), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(new_n759), .B2(new_n796), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n791), .A2(new_n792), .B1(new_n794), .B2(new_n797), .ZN(G1339gat));
  NOR2_X1   g597(.A1(new_n605), .A2(new_n607), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT112), .Z(new_n800));
  AOI21_X1  g599(.A(new_n606), .B1(new_n615), .B2(new_n616), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n623), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n629), .A2(new_n631), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n803), .A3(new_n578), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n565), .A2(new_n563), .A3(new_n566), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n568), .A2(KEYINPUT54), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n574), .B1(new_n567), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n806), .A2(KEYINPUT55), .A3(new_n808), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n577), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n804), .B1(new_n633), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n552), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n802), .A2(new_n803), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(new_n552), .A3(new_n813), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n602), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n603), .A2(new_n723), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n728), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n411), .A2(new_n489), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n420), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT114), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n633), .A2(G113gat), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n633), .A2(new_n813), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n667), .B1(new_n829), .B2(new_n804), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n724), .B1(new_n830), .B2(new_n817), .ZN(new_n831));
  INV_X1    g630(.A(new_n820), .ZN(new_n832));
  AOI211_X1 g631(.A(new_n715), .B(new_n478), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n637), .A2(new_n421), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(G113gat), .B1(new_n835), .B2(new_n633), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(KEYINPUT113), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(KEYINPUT113), .ZN(new_n838));
  OAI22_X1  g637(.A1(new_n827), .A2(new_n828), .B1(new_n837), .B2(new_n838), .ZN(G1340gat));
  OAI21_X1  g638(.A(G120gat), .B1(new_n835), .B2(new_n579), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n579), .A2(G120gat), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n827), .B2(new_n841), .ZN(G1341gat));
  OR3_X1    g641(.A1(new_n825), .A2(G127gat), .A3(new_n724), .ZN(new_n843));
  OAI21_X1  g642(.A(G127gat), .B1(new_n835), .B2(new_n724), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1342gat));
  OR3_X1    g644(.A1(new_n825), .A2(G134gat), .A3(new_n552), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n833), .A2(new_n667), .A3(new_n834), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n846), .A2(KEYINPUT56), .B1(G134gat), .B2(new_n847), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n825), .A2(G134gat), .A3(new_n552), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT56), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n849), .A2(KEYINPUT115), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT115), .B1(new_n849), .B2(new_n850), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(G1343gat));
  NAND2_X1  g652(.A1(new_n652), .A2(new_n834), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n821), .B2(new_n411), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n831), .A2(new_n832), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(KEYINPUT57), .A3(new_n715), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n854), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n203), .B1(new_n859), .B2(new_n723), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n653), .A2(new_n421), .A3(new_n411), .ZN(new_n861));
  AND4_X1   g660(.A1(new_n203), .A2(new_n822), .A3(new_n723), .A4(new_n861), .ZN(new_n862));
  OR3_X1    g661(.A1(new_n860), .A2(KEYINPUT58), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT58), .B1(new_n860), .B2(new_n862), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1344gat));
  NAND4_X1  g664(.A1(new_n822), .A2(new_n204), .A3(new_n578), .A4(new_n861), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT116), .Z(new_n867));
  INV_X1    g666(.A(new_n854), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n821), .A2(new_n855), .A3(new_n657), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT57), .B1(new_n857), .B2(new_n410), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n578), .B(new_n868), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n872), .A3(G148gat), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n854), .A2(new_n579), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n552), .A2(new_n813), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n816), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT117), .B1(new_n552), .B2(new_n813), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n877), .A2(new_n878), .B1(new_n814), .B2(new_n552), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n832), .B1(new_n879), .B2(new_n602), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT57), .B1(new_n880), .B2(new_n715), .ZN(new_n881));
  OAI211_X1 g680(.A(KEYINPUT57), .B(new_n410), .C1(new_n819), .C2(new_n820), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n874), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n872), .B1(new_n884), .B2(G148gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n873), .B1(new_n885), .B2(KEYINPUT118), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  AOI211_X1 g686(.A(new_n887), .B(new_n872), .C1(new_n884), .C2(G148gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n867), .B1(new_n886), .B2(new_n888), .ZN(G1345gat));
  AND2_X1   g688(.A1(new_n822), .A2(new_n861), .ZN(new_n890));
  INV_X1    g689(.A(G155gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n891), .A3(new_n602), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n859), .A2(new_n602), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n891), .ZN(G1346gat));
  NOR2_X1   g693(.A1(new_n552), .A2(G162gat), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT119), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n859), .A2(new_n667), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT120), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G162gat), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n898), .A2(KEYINPUT120), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(G1347gat));
  NAND2_X1  g701(.A1(new_n823), .A2(new_n421), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n821), .A2(new_n638), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(G169gat), .B1(new_n904), .B2(new_n723), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n727), .A2(new_n420), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n833), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n633), .A2(new_n296), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(G1348gat));
  AOI21_X1  g709(.A(G176gat), .B1(new_n904), .B2(new_n578), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT121), .Z(new_n912));
  NOR3_X1   g711(.A1(new_n907), .A2(new_n297), .A3(new_n579), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(G1349gat));
  OAI21_X1  g713(.A(G183gat), .B1(new_n907), .B2(new_n724), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n904), .A2(new_n288), .A3(new_n602), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n904), .A2(new_n289), .A3(new_n667), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n289), .B1(new_n908), .B2(new_n667), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(G1351gat));
  AOI21_X1  g723(.A(new_n638), .B1(new_n831), .B2(new_n832), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n652), .A2(new_n421), .A3(new_n410), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n925), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(G197gat), .B1(new_n930), .B2(new_n723), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n881), .A2(new_n883), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n906), .A2(new_n652), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT123), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n633), .A2(new_n317), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(G1352gat));
  NAND3_X1  g736(.A1(new_n932), .A2(new_n578), .A3(new_n934), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n930), .A2(new_n315), .A3(new_n578), .ZN(new_n939));
  AOI22_X1  g738(.A1(new_n938), .A2(G204gat), .B1(KEYINPUT62), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n939), .A2(KEYINPUT62), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n939), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(G1353gat));
  INV_X1    g744(.A(G211gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n946), .A3(new_n602), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n602), .B(new_n934), .C1(new_n881), .C2(new_n883), .ZN(new_n948));
  AND4_X1   g747(.A1(KEYINPUT125), .A2(new_n948), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n949));
  OAI21_X1  g748(.A(G211gat), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  AOI22_X1  g750(.A1(new_n948), .A2(new_n951), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n947), .B1(new_n949), .B2(new_n952), .ZN(G1354gat));
  INV_X1    g752(.A(G218gat), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n552), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n934), .B(new_n955), .C1(new_n881), .C2(new_n883), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n925), .A2(new_n929), .A3(new_n667), .A4(new_n928), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n957), .A2(KEYINPUT126), .A3(new_n954), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT126), .B1(new_n957), .B2(new_n954), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g761(.A(KEYINPUT127), .B(new_n956), .C1(new_n958), .C2(new_n959), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1355gat));
endmodule


