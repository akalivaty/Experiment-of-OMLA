//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT22), .ZN(new_n207));
  INV_X1    g006(.A(G211gat), .ZN(new_n208));
  INV_X1    g007(.A(G218gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(G211gat), .B(G218gat), .Z(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT69), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n212), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AND2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G141gat), .B(G148gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n219), .B1(new_n220), .B2(KEYINPUT2), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT29), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT78), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT72), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n226), .B(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT77), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n214), .A2(new_n238), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n214), .A2(new_n238), .B1(new_n212), .B2(new_n211), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT29), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n237), .B1(new_n241), .B2(KEYINPUT3), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n234), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G228gat), .A2(G233gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G22gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n228), .B1(new_n216), .B2(KEYINPUT29), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n226), .ZN(new_n248));
  INV_X1    g047(.A(new_n244), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n249), .A3(new_n232), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n245), .A2(new_n246), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n249), .B1(new_n234), .B2(new_n242), .ZN(new_n252));
  INV_X1    g051(.A(new_n250), .ZN(new_n253));
  OAI21_X1  g052(.A(G22gat), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(KEYINPUT76), .B(KEYINPUT31), .Z(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n255), .B1(new_n251), .B2(new_n254), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n205), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n258), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(new_n204), .A3(new_n256), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT27), .B(G183gat), .ZN(new_n263));
  INV_X1    g062(.A(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n265), .B(KEYINPUT28), .Z(new_n266));
  AND2_X1   g065(.A1(G183gat), .A2(G190gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n269), .A2(KEYINPUT26), .ZN(new_n270));
  AND2_X1   g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n269), .B1(new_n271), .B2(KEYINPUT26), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n267), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT23), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n271), .B1(new_n269), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT24), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n277), .A2(new_n267), .B1(new_n268), .B2(KEYINPUT23), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n276), .B(new_n278), .C1(new_n267), .C2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT25), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n274), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(G113gat), .B(G120gat), .Z(new_n284));
  INV_X1    g083(.A(KEYINPUT1), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G127gat), .B(G134gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT65), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n283), .B(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G227gat), .A2(G233gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n296), .B(KEYINPUT64), .Z(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT33), .ZN(new_n299));
  XNOR2_X1  g098(.A(G15gat), .B(G43gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(KEYINPUT68), .ZN(new_n301));
  XOR2_X1   g100(.A(G71gat), .B(G99gat), .Z(new_n302));
  XOR2_X1   g101(.A(new_n301), .B(new_n302), .Z(new_n303));
  OAI211_X1 g102(.A(new_n298), .B(KEYINPUT32), .C1(new_n299), .C2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n305), .B1(new_n298), .B2(new_n299), .ZN(new_n306));
  INV_X1    g105(.A(new_n297), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n294), .A2(new_n307), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n308), .A2(KEYINPUT66), .A3(KEYINPUT33), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n298), .A2(KEYINPUT67), .A3(KEYINPUT32), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT67), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT32), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n303), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n304), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  OR3_X1    g116(.A1(new_n295), .A2(KEYINPUT34), .A3(new_n297), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n294), .A2(new_n296), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT34), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n321), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n323), .B(new_n304), .C1(new_n310), .C2(new_n316), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n291), .A2(new_n226), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n291), .A2(new_n226), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT5), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n293), .A2(new_n236), .A3(KEYINPUT4), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n226), .A2(KEYINPUT3), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n229), .A2(new_n291), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT4), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n331), .B1(new_n327), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n334), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  OR2_X1    g138(.A1(new_n339), .A2(KEYINPUT73), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(KEYINPUT73), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n333), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n336), .B1(new_n337), .B2(new_n327), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT4), .B1(new_n293), .B2(new_n236), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n345), .A2(KEYINPUT5), .A3(new_n331), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G1gat), .B(G29gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT0), .ZN(new_n350));
  XNOR2_X1  g149(.A(G57gat), .B(G85gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT6), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(new_n347), .B2(new_n352), .ZN(new_n357));
  NOR4_X1   g156(.A1(new_n342), .A2(new_n346), .A3(KEYINPUT74), .A4(new_n353), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n354), .B(new_n355), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(KEYINPUT6), .B(new_n353), .C1(new_n342), .C2(new_n346), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT75), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G226gat), .A2(G233gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n283), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n230), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(new_n274), .B2(new_n282), .ZN(new_n366));
  OR3_X1    g165(.A1(new_n364), .A2(new_n216), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n216), .B1(new_n364), .B2(new_n366), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G8gat), .B(G36gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n369), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(new_n372), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n376), .B2(KEYINPUT30), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT71), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT70), .B1(new_n369), .B2(new_n373), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT70), .ZN(new_n380));
  AOI211_X1 g179(.A(new_n380), .B(new_n372), .C1(new_n367), .C2(new_n368), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR4_X1   g183(.A1(new_n379), .A2(new_n381), .A3(KEYINPUT71), .A4(KEYINPUT30), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n377), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n262), .A2(new_n326), .A3(new_n362), .A4(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT35), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n389), .B(new_n377), .C1(new_n384), .C2(new_n385), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n352), .B(KEYINPUT79), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n348), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n393), .B(new_n355), .C1(new_n357), .C2(new_n358), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n390), .B1(new_n361), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n325), .B1(new_n261), .B2(new_n259), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n388), .A2(KEYINPUT35), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n262), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n362), .A2(new_n387), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n373), .B1(new_n375), .B2(KEYINPUT37), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT38), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT37), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n403), .B1(new_n369), .B2(new_n404), .ZN(new_n405));
  AOI211_X1 g204(.A(KEYINPUT82), .B(KEYINPUT37), .C1(new_n367), .C2(new_n368), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n401), .B(new_n402), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n382), .ZN(new_n408));
  INV_X1    g207(.A(new_n405), .ZN(new_n409));
  INV_X1    g208(.A(new_n406), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n402), .B1(new_n411), .B2(new_n401), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n413), .A2(new_n394), .A3(new_n361), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n343), .A2(new_n344), .ZN(new_n415));
  OR3_X1    g214(.A1(new_n415), .A2(KEYINPUT39), .A3(new_n330), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n330), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n327), .A2(new_n330), .A3(new_n328), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT80), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n419), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(KEYINPUT39), .A3(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n416), .B(new_n391), .C1(new_n417), .C2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT40), .ZN(new_n424));
  OR3_X1    g223(.A1(new_n423), .A2(KEYINPUT81), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT81), .B1(new_n423), .B2(new_n424), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n348), .A2(new_n392), .B1(new_n423), .B2(new_n424), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n386), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n414), .A2(new_n262), .A3(KEYINPUT83), .A4(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT36), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n325), .B(new_n431), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n400), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n262), .A3(new_n429), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT83), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n397), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n246), .A2(G15gat), .ZN(new_n438));
  INV_X1    g237(.A(G15gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(G22gat), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT16), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n438), .A2(new_n440), .A3(KEYINPUT87), .ZN(new_n443));
  INV_X1    g242(.A(G1gat), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G15gat), .B(G22gat), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n446), .B(KEYINPUT87), .C1(new_n441), .C2(G1gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G8gat), .ZN(new_n449));
  INV_X1    g248(.A(G8gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  OR3_X1    g252(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G29gat), .A2(G36gat), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(G43gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n203), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT15), .ZN(new_n461));
  NAND2_X1  g260(.A1(G43gat), .A2(G50gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n460), .A2(KEYINPUT86), .A3(new_n461), .A4(new_n462), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n468));
  INV_X1    g267(.A(new_n462), .ZN(new_n469));
  NOR2_X1   g268(.A1(G43gat), .A2(G50gat), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n460), .A2(KEYINPUT85), .A3(new_n462), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n458), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n457), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n471), .A2(new_n472), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(new_n461), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n474), .A2(KEYINPUT17), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT17), .B1(new_n474), .B2(new_n477), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n453), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT88), .ZN(new_n481));
  NAND2_X1  g280(.A1(G229gat), .A2(G233gat), .ZN(new_n482));
  XOR2_X1   g281(.A(new_n482), .B(KEYINPUT89), .Z(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n485), .B(new_n453), .C1(new_n478), .C2(new_n479), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n445), .A2(new_n447), .A3(new_n450), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n450), .B1(new_n445), .B2(new_n447), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n474), .B(new_n477), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT90), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT90), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n452), .A2(new_n491), .A3(new_n474), .A4(new_n477), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n481), .A2(new_n484), .A3(new_n486), .A4(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT18), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n474), .A2(new_n477), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT17), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n474), .A2(new_n477), .A3(KEYINPUT17), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n452), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n501), .A2(new_n485), .B1(new_n490), .B2(new_n492), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n502), .A2(KEYINPUT18), .A3(new_n484), .A4(new_n481), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n453), .A2(new_n497), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n493), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n483), .B(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n496), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(G113gat), .B(G141gat), .Z(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT11), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(G169gat), .ZN(new_n512));
  XOR2_X1   g311(.A(KEYINPUT84), .B(G197gat), .Z(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G169gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n511), .B(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n513), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n515), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n515), .B2(new_n518), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n509), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n496), .A2(new_n503), .A3(new_n508), .A4(new_n522), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n524), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n505), .A2(new_n507), .ZN(new_n532));
  AND4_X1   g331(.A1(new_n484), .A2(new_n481), .A3(new_n486), .A4(new_n493), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(KEYINPUT18), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n534), .A2(KEYINPUT92), .A3(new_n496), .A4(new_n522), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n525), .A2(new_n526), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(KEYINPUT93), .A3(new_n524), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G183gat), .B(G211gat), .Z(new_n541));
  XNOR2_X1  g340(.A(G71gat), .B(G78gat), .ZN(new_n542));
  XOR2_X1   g341(.A(G57gat), .B(G64gat), .Z(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(KEYINPUT9), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT94), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT94), .ZN(new_n546));
  XNOR2_X1  g345(.A(G57gat), .B(G64gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT9), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n546), .B1(new_n549), .B2(new_n542), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G71gat), .ZN(new_n552));
  INV_X1    g351(.A(G78gat), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n548), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n543), .A2(new_n542), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT95), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n543), .A2(KEYINPUT95), .A3(new_n542), .A4(new_n554), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n551), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(KEYINPUT96), .B(KEYINPUT21), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G231gat), .A2(G233gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n565), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n551), .A2(KEYINPUT21), .A3(new_n559), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n453), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n569), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n566), .A2(new_n567), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n572), .B1(new_n570), .B2(new_n574), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n541), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n577), .ZN(new_n579));
  INV_X1    g378(.A(new_n541), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n575), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G134gat), .B(G162gat), .Z(new_n583));
  AND2_X1   g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT41), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n583), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(KEYINPUT98), .B(G92gat), .Z(new_n588));
  INV_X1    g387(.A(G85gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(G99gat), .A2(G106gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n588), .A2(new_n589), .B1(KEYINPUT8), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT97), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT7), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n592), .B(KEYINPUT97), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT7), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n591), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G99gat), .B(G106gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n591), .A2(new_n595), .A3(new_n598), .A4(new_n600), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(new_n497), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(KEYINPUT41), .B2(new_n584), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n604), .B1(new_n478), .B2(new_n479), .ZN(new_n607));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT99), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n606), .A2(new_n607), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n612), .A2(new_n613), .B1(new_n614), .B2(new_n608), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT100), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n587), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n612), .A2(new_n613), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n608), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT100), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(KEYINPUT100), .A3(new_n587), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n604), .A2(new_n560), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n602), .A2(new_n559), .A3(new_n551), .A4(new_n603), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n628), .A2(KEYINPUT102), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(KEYINPUT102), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n626), .A2(new_n636), .A3(new_n627), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n627), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n625), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT101), .ZN(new_n641));
  INV_X1    g440(.A(new_n625), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n642), .B1(new_n637), .B2(new_n638), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n631), .A2(new_n635), .A3(new_n641), .A4(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n640), .A2(new_n629), .A3(new_n630), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n634), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n582), .A2(new_n624), .A3(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n437), .A2(new_n540), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n362), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G1gat), .ZN(G1324gat));
  INV_X1    g453(.A(KEYINPUT103), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n436), .A2(new_n430), .A3(new_n400), .A4(new_n432), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n388), .A2(KEYINPUT35), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n396), .A2(new_n395), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n650), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n660), .A2(new_n386), .A3(new_n539), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT16), .B(G8gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT104), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n655), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT42), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n662), .A2(G8gat), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(new_n665), .B2(KEYINPUT42), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT105), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n665), .A2(KEYINPUT42), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n671), .A2(new_n672), .A3(new_n666), .A4(new_n668), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(G1325gat));
  INV_X1    g473(.A(new_n651), .ZN(new_n675));
  OAI21_X1  g474(.A(G15gat), .B1(new_n675), .B2(new_n432), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n651), .A2(new_n439), .A3(new_n326), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(G1326gat));
  NAND2_X1  g477(.A1(new_n651), .A2(new_n398), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n437), .B2(new_n624), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n624), .B1(new_n656), .B2(new_n659), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT44), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n582), .B(KEYINPUT106), .ZN(new_n686));
  INV_X1    g485(.A(new_n529), .ZN(new_n687));
  INV_X1    g486(.A(new_n649), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n683), .A2(new_n685), .A3(new_n652), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G29gat), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n582), .A2(new_n624), .A3(new_n688), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n362), .A2(G29gat), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n660), .A2(new_n539), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT45), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT107), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n691), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(G1328gat));
  XNOR2_X1  g499(.A(new_n684), .B(new_n682), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n386), .A3(new_n689), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G36gat), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n387), .A2(G36gat), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n660), .A2(new_n539), .A3(new_n692), .A4(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n707), .A2(KEYINPUT46), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT46), .B1(new_n707), .B2(new_n708), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n703), .B1(new_n709), .B2(new_n710), .ZN(G1329gat));
  NOR2_X1   g510(.A1(new_n432), .A2(new_n459), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n683), .A2(new_n685), .A3(new_n689), .A4(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n660), .A2(new_n539), .A3(new_n692), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n459), .B1(new_n714), .B2(new_n325), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1330gat));
  NAND4_X1  g517(.A1(new_n701), .A2(G50gat), .A3(new_n398), .A4(new_n689), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n203), .B1(new_n714), .B2(new_n262), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n719), .A2(KEYINPUT48), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT48), .B1(new_n719), .B2(new_n720), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(G1331gat));
  INV_X1    g522(.A(new_n582), .ZN(new_n724));
  INV_X1    g523(.A(new_n624), .ZN(new_n725));
  NOR4_X1   g524(.A1(new_n724), .A2(new_n725), .A3(new_n529), .A4(new_n649), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n660), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n362), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT110), .B(G57gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1332gat));
  INV_X1    g529(.A(new_n727), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n387), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT111), .Z(new_n735));
  XNOR2_X1  g534(.A(new_n733), .B(new_n735), .ZN(G1333gat));
  OAI21_X1  g535(.A(G71gat), .B1(new_n727), .B2(new_n432), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n326), .A2(new_n552), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n727), .B2(new_n738), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g539(.A1(new_n727), .A2(new_n262), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(new_n553), .ZN(G1335gat));
  NOR3_X1   g541(.A1(new_n582), .A2(new_n529), .A3(new_n649), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n701), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G85gat), .B1(new_n744), .B2(new_n362), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n582), .A2(new_n529), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT51), .B1(new_n684), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n684), .A2(KEYINPUT51), .A3(new_n746), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n748), .A2(KEYINPUT112), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT112), .B1(new_n748), .B2(new_n749), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n688), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n652), .A2(new_n589), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n745), .B1(new_n752), .B2(new_n753), .ZN(G1336gat));
  OR2_X1    g553(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n683), .A2(new_n685), .A3(new_n386), .A4(new_n743), .ZN(new_n756));
  INV_X1    g555(.A(new_n588), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n387), .A2(G92gat), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n684), .A2(KEYINPUT51), .A3(new_n746), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n688), .B(new_n759), .C1(new_n760), .C2(new_n747), .ZN(new_n761));
  NAND2_X1  g560(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n762));
  AND4_X1   g561(.A1(new_n755), .A2(new_n758), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  AOI22_X1  g562(.A1(new_n756), .A2(new_n757), .B1(KEYINPUT113), .B2(KEYINPUT52), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n755), .B1(new_n764), .B2(new_n761), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n763), .A2(new_n765), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n744), .B2(new_n432), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n325), .A2(G99gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n752), .B2(new_n768), .ZN(G1338gat));
  INV_X1    g568(.A(G106gat), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n701), .A2(KEYINPUT114), .A3(new_n398), .A4(new_n743), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n683), .A2(new_n685), .A3(new_n398), .A4(new_n743), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n770), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n262), .A2(G106gat), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n688), .B(new_n776), .C1(new_n760), .C2(new_n747), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n772), .A2(G106gat), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(new_n777), .ZN(new_n781));
  OAI22_X1  g580(.A1(new_n775), .A2(new_n779), .B1(new_n781), .B2(new_n778), .ZN(G1339gat));
  NOR2_X1   g581(.A1(new_n650), .A2(new_n529), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n484), .B1(new_n502), .B2(new_n481), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n505), .A2(new_n507), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n515), .B(new_n518), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n537), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n649), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n637), .A2(new_n638), .A3(new_n642), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n641), .A2(KEYINPUT54), .A3(new_n645), .A4(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  AOI211_X1 g592(.A(new_n792), .B(new_n635), .C1(new_n643), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n643), .A2(new_n793), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT115), .B1(new_n795), .B2(new_n634), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n791), .B(KEYINPUT55), .C1(new_n794), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n646), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT116), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n646), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n795), .A2(new_n634), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n792), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n795), .A2(KEYINPUT115), .A3(new_n634), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT55), .B1(new_n805), .B2(new_n791), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n799), .A2(new_n801), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n789), .B1(new_n808), .B2(new_n687), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n624), .ZN(new_n810));
  INV_X1    g609(.A(new_n787), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n806), .B1(new_n798), .B2(KEYINPUT116), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n725), .A2(new_n811), .A3(new_n801), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n686), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n783), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(new_n362), .A3(new_n386), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n396), .ZN(new_n818));
  OAI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n540), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n819), .B(KEYINPUT117), .Z(new_n820));
  XNOR2_X1  g619(.A(new_n818), .B(KEYINPUT118), .ZN(new_n821));
  INV_X1    g620(.A(G113gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n822), .A3(new_n529), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n823), .ZN(G1340gat));
  OAI21_X1  g623(.A(G120gat), .B1(new_n818), .B2(new_n649), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT119), .ZN(new_n826));
  INV_X1    g625(.A(G120gat), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n821), .A2(new_n827), .A3(new_n688), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(G1341gat));
  NOR3_X1   g628(.A1(new_n818), .A2(KEYINPUT120), .A3(new_n724), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(G127gat), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT120), .B1(new_n818), .B2(new_n724), .ZN(new_n832));
  INV_X1    g631(.A(new_n818), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n686), .A2(G127gat), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n831), .A2(new_n832), .B1(new_n833), .B2(new_n834), .ZN(G1342gat));
  AOI21_X1  g634(.A(new_n624), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n817), .A2(new_n396), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n837), .B(new_n838), .Z(G1343gat));
  AND3_X1   g638(.A1(new_n432), .A2(new_n652), .A3(new_n387), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n262), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n783), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n798), .A2(new_n806), .ZN(new_n844));
  AOI221_X4 g643(.A(new_n530), .B1(new_n509), .B2(new_n523), .C1(new_n535), .C2(new_n536), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT93), .B1(new_n537), .B2(new_n524), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n725), .B1(new_n847), .B2(new_n789), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n808), .A2(new_n624), .A3(new_n787), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n724), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n843), .B1(new_n850), .B2(KEYINPUT121), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n788), .B1(new_n539), .B2(new_n844), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n813), .B1(new_n853), .B2(new_n725), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n852), .B1(new_n854), .B2(new_n724), .ZN(new_n855));
  OAI211_X1 g654(.A(KEYINPUT122), .B(new_n842), .C1(new_n851), .C2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n841), .B1(new_n816), .B2(new_n262), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n850), .A2(KEYINPUT121), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n854), .A2(new_n852), .A3(new_n724), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n860), .A3(new_n843), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT122), .B1(new_n861), .B2(new_n842), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n840), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(G141gat), .B1(new_n863), .B2(new_n540), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n432), .A2(new_n398), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n817), .A2(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n866), .A2(G141gat), .A3(new_n540), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(KEYINPUT58), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n529), .B(new_n840), .C1(new_n858), .C2(new_n862), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n867), .B1(G141gat), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(G1344gat));
  INV_X1    g672(.A(G148gat), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n817), .A2(new_n874), .A3(new_n688), .A4(new_n865), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n688), .B(new_n840), .C1(new_n858), .C2(new_n862), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(KEYINPUT59), .A3(new_n874), .ZN(new_n878));
  XOR2_X1   g677(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n879));
  NOR2_X1   g678(.A1(new_n650), .A2(new_n539), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n262), .B1(new_n850), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT124), .B1(new_n882), .B2(KEYINPUT57), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n880), .B1(new_n854), .B2(new_n724), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n884), .B(new_n841), .C1(new_n885), .C2(new_n262), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n686), .B1(new_n810), .B2(new_n813), .ZN(new_n887));
  OAI211_X1 g686(.A(KEYINPUT57), .B(new_n398), .C1(new_n887), .C2(new_n783), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n883), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n688), .A3(new_n840), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n879), .B1(new_n890), .B2(G148gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n875), .B1(new_n878), .B2(new_n891), .ZN(G1345gat));
  OAI21_X1  g691(.A(G155gat), .B1(new_n863), .B2(new_n815), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n724), .A2(G155gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n866), .B2(new_n894), .ZN(G1346gat));
  OAI211_X1 g694(.A(new_n725), .B(new_n840), .C1(new_n858), .C2(new_n862), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(G162gat), .ZN(new_n897));
  OR3_X1    g696(.A1(new_n866), .A2(G162gat), .A3(new_n624), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n897), .A2(KEYINPUT125), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1347gat));
  NAND2_X1  g702(.A1(new_n814), .A2(new_n815), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n843), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n652), .A2(new_n387), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n905), .A2(new_n396), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(G169gat), .B1(new_n907), .B2(new_n529), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n540), .A2(new_n516), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n907), .B2(new_n909), .ZN(G1348gat));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n688), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g711(.A1(new_n907), .A2(new_n686), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G183gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n907), .A2(new_n263), .A3(new_n582), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g716(.A1(new_n907), .A2(new_n725), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G190gat), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT61), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(G190gat), .B2(new_n918), .ZN(G1351gat));
  AND3_X1   g720(.A1(new_n905), .A2(new_n865), .A3(new_n906), .ZN(new_n922));
  AOI21_X1  g721(.A(G197gat), .B1(new_n922), .B2(new_n529), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n906), .A2(new_n432), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n889), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n539), .A2(G197gat), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1352gat));
  NOR2_X1   g726(.A1(new_n649), .A2(G204gat), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n905), .A2(new_n865), .A3(new_n906), .A4(new_n928), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT62), .Z(new_n930));
  NAND3_X1  g729(.A1(new_n889), .A2(new_n688), .A3(new_n924), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G204gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT126), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n930), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1353gat));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n208), .A3(new_n582), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n889), .A2(new_n582), .A3(new_n924), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(KEYINPUT127), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943));
  AOI211_X1 g742(.A(new_n943), .B(KEYINPUT63), .C1(new_n939), .C2(G211gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n938), .B1(new_n942), .B2(new_n944), .ZN(G1354gat));
  NAND3_X1  g744(.A1(new_n922), .A2(new_n209), .A3(new_n725), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n925), .A2(new_n725), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n947), .B2(new_n209), .ZN(G1355gat));
endmodule


