//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G122), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT92), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G122), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G107), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n190), .A2(new_n195), .A3(new_n192), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT68), .B(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n199), .B(KEYINPUT93), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G128), .ZN(new_n202));
  XNOR2_X1  g016(.A(new_n202), .B(KEYINPUT13), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n197), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT65), .A2(G134), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT65), .A2(G134), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n200), .A2(new_n209), .A3(new_n202), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(new_n196), .A2(KEYINPUT94), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n196), .A2(KEYINPUT94), .ZN(new_n215));
  INV_X1    g029(.A(new_n190), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n192), .B(KEYINPUT14), .ZN(new_n217));
  OAI21_X1  g031(.A(G107), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n214), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n200), .A2(new_n202), .ZN(new_n220));
  OR2_X1    g034(.A1(KEYINPUT65), .A2(G134), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT65), .A2(G134), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n219), .B1(new_n210), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT9), .B(G234), .ZN(new_n227));
  INV_X1    g041(.A(G217), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n227), .A2(new_n228), .A3(G953), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n213), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n229), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n212), .B2(new_n225), .ZN(new_n232));
  AOI21_X1  g046(.A(G902), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G478), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(KEYINPUT15), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n233), .B(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  INV_X1    g052(.A(G140), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G125), .ZN(new_n240));
  INV_X1    g054(.A(G125), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G140), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n240), .A2(new_n242), .A3(KEYINPUT75), .A4(KEYINPUT16), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n240), .A2(new_n242), .A3(KEYINPUT16), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT75), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n245), .B1(new_n240), .B2(KEYINPUT16), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n243), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G146), .ZN(new_n248));
  INV_X1    g062(.A(G146), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n249), .B(new_n243), .C1(new_n244), .C2(new_n246), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G237), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G214), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(new_n201), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT17), .A3(G131), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n254), .B(G143), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n251), .B(new_n256), .C1(KEYINPUT17), .C2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT18), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n257), .B1(new_n261), .B2(new_n258), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n255), .A2(KEYINPUT18), .A3(G131), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n240), .A2(new_n242), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(G146), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G113), .B(G122), .ZN(new_n267));
  INV_X1    g081(.A(G104), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(KEYINPUT91), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n260), .A2(new_n266), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n269), .B1(new_n260), .B2(new_n266), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n238), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G475), .ZN(new_n275));
  INV_X1    g089(.A(new_n264), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT19), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(KEYINPUT90), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT90), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(new_n264), .B2(KEYINPUT19), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n278), .B(new_n280), .C1(new_n277), .C2(new_n276), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n259), .B(new_n248), .C1(G146), .C2(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n282), .A2(new_n266), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n271), .B1(new_n283), .B2(new_n269), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT20), .ZN(new_n285));
  NOR2_X1   g099(.A1(G475), .A2(G902), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n275), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n253), .A2(G952), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(G234), .B2(G237), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT21), .B(G898), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G234), .ZN(new_n295));
  OAI211_X1 g109(.A(G902), .B(G953), .C1(new_n295), .C2(new_n252), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n292), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  XOR2_X1   g111(.A(new_n297), .B(KEYINPUT95), .Z(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n237), .A2(new_n289), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT64), .ZN(new_n301));
  XNOR2_X1  g115(.A(G143), .B(G146), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT0), .B(G128), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n249), .A2(G143), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n201), .A2(G146), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(KEYINPUT0), .A2(G128), .ZN(new_n308));
  OR2_X1    g122(.A1(KEYINPUT0), .A2(G128), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n307), .A2(KEYINPUT64), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n302), .A2(KEYINPUT0), .A3(G128), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n304), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G125), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT1), .B1(new_n201), .B2(G146), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G128), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT68), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT68), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G128), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n305), .A2(KEYINPUT67), .A3(KEYINPUT1), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n316), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n307), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT1), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n302), .A2(new_n325), .A3(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n313), .B1(new_n327), .B2(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT86), .ZN(new_n329));
  INV_X1    g143(.A(G224), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(G953), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT86), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n313), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n329), .A2(KEYINPUT7), .A3(new_n332), .A4(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT7), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n328), .B1(new_n336), .B2(new_n331), .ZN(new_n337));
  XNOR2_X1  g151(.A(G110), .B(G122), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT8), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n195), .A2(G104), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n195), .A2(G104), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n340), .B1(KEYINPUT3), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G101), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n195), .A3(G104), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n342), .A2(KEYINPUT82), .A3(new_n343), .A4(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT3), .B1(new_n268), .B2(G107), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n268), .A2(G107), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n347), .A2(new_n345), .A3(new_n343), .A4(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n341), .A2(new_n348), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n346), .A2(new_n351), .B1(G101), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n191), .A2(G119), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT70), .ZN(new_n355));
  INV_X1    g169(.A(G119), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n355), .B1(new_n356), .B2(G116), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n191), .A2(KEYINPUT70), .A3(G119), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n354), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT5), .ZN(new_n360));
  INV_X1    g174(.A(G113), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT5), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n361), .B1(new_n354), .B2(new_n362), .ZN(new_n363));
  XOR2_X1   g177(.A(KEYINPUT2), .B(G113), .Z(new_n364));
  AOI22_X1  g178(.A1(new_n360), .A2(new_n363), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n353), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n353), .A2(new_n365), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n339), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n335), .A2(new_n337), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT88), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n359), .B(new_n364), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n347), .A2(new_n345), .A3(new_n348), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT81), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n347), .A2(new_n345), .A3(KEYINPUT81), .A4(new_n348), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(G101), .A3(new_n377), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n378), .A2(KEYINPUT4), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n346), .A2(new_n351), .ZN(new_n381));
  AND4_X1   g195(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT4), .A4(new_n378), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(new_n346), .B2(new_n351), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n380), .B1(new_n384), .B2(new_n378), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n373), .B(new_n379), .C1(new_n382), .C2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n338), .A3(new_n366), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n335), .A2(KEYINPUT88), .A3(new_n337), .A4(new_n369), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n372), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n238), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(new_n366), .ZN(new_n391));
  INV_X1    g205(.A(new_n338), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT6), .A3(new_n387), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n395), .A3(new_n392), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n329), .A2(new_n334), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(new_n331), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT87), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n394), .A2(KEYINPUT87), .A3(new_n396), .A4(new_n398), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n390), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(G210), .B1(G237), .B2(G902), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(KEYINPUT89), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n404), .ZN(new_n408));
  AOI211_X1 g222(.A(new_n408), .B(new_n390), .C1(new_n401), .C2(new_n402), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n187), .B(new_n300), .C1(new_n407), .C2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G469), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n412));
  XNOR2_X1  g226(.A(G110), .B(G140), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n253), .A2(G227), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n413), .B(new_n414), .Z(new_n415));
  INV_X1    g229(.A(KEYINPUT71), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n312), .B(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n417), .B(new_n379), .C1(new_n382), .C2(new_n385), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT66), .ZN(new_n419));
  AOI21_X1  g233(.A(G137), .B1(new_n221), .B2(new_n222), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n419), .B1(new_n420), .B2(KEYINPUT11), .ZN(new_n421));
  INV_X1    g235(.A(G137), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n207), .B2(new_n208), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT11), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(KEYINPUT66), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(KEYINPUT11), .A3(G134), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n427), .B1(G137), .B2(new_n209), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n421), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G131), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n421), .A2(new_n425), .A3(new_n428), .A4(new_n258), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT10), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n352), .A2(G101), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n317), .B1(new_n305), .B2(KEYINPUT1), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n326), .B1(new_n436), .B2(new_n302), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n349), .A2(new_n350), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n349), .A2(new_n350), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n435), .B(new_n437), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n434), .B1(new_n324), .B2(new_n326), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n434), .A2(new_n440), .B1(new_n441), .B2(new_n353), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n418), .A2(new_n433), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n433), .B1(new_n418), .B2(new_n442), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n412), .B(new_n415), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n440), .B1(new_n353), .B2(new_n327), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n432), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT12), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(KEYINPUT12), .A3(new_n432), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(KEYINPUT84), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n418), .A2(new_n433), .A3(new_n442), .ZN(new_n452));
  INV_X1    g266(.A(new_n415), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n447), .A2(new_n454), .A3(new_n448), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n451), .A2(new_n452), .A3(new_n453), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n445), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n418), .A2(new_n442), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n432), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n452), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n412), .B1(new_n460), .B2(new_n415), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n411), .B(new_n238), .C1(new_n457), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(G469), .A2(G902), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n451), .A2(new_n452), .A3(new_n455), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n415), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n459), .A2(new_n452), .A3(new_n453), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n462), .B(new_n463), .C1(new_n411), .C2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G221), .ZN(new_n469));
  INV_X1    g283(.A(new_n227), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(new_n238), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n410), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(KEYINPUT23), .B1(new_n317), .B2(G119), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n317), .A2(G119), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT23), .A4(G119), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OR3_X1    g293(.A1(new_n479), .A2(KEYINPUT77), .A3(G110), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n476), .B1(new_n198), .B2(G119), .ZN(new_n481));
  XOR2_X1   g295(.A(KEYINPUT24), .B(G110), .Z(new_n482));
  OR3_X1    g296(.A1(new_n481), .A2(KEYINPUT78), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT77), .B1(new_n479), .B2(G110), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT78), .B1(new_n481), .B2(new_n482), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n480), .A2(new_n483), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n276), .A2(new_n249), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n248), .A3(new_n487), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n248), .A2(new_n250), .B1(new_n481), .B2(new_n482), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n479), .A2(G110), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT74), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT74), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n479), .A2(new_n492), .A3(G110), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n489), .A2(KEYINPUT76), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(KEYINPUT76), .B1(new_n489), .B2(new_n494), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n488), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT22), .B(G137), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n469), .A2(new_n295), .A3(G953), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n498), .B(new_n499), .Z(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n488), .B(new_n500), .C1(new_n495), .C2(new_n496), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n238), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT79), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT25), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n228), .B1(G234), .B2(new_n238), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n506), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n502), .A2(KEYINPUT25), .A3(new_n238), .A4(new_n503), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(KEYINPUT79), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n508), .A2(G902), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n514), .B(KEYINPUT80), .Z(new_n515));
  NAND3_X1  g329(.A1(new_n502), .A2(new_n515), .A3(new_n503), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n324), .A2(new_n326), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n422), .A2(G134), .ZN(new_n519));
  OAI21_X1  g333(.A(G131), .B1(new_n420), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n431), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n518), .B1(new_n521), .B2(KEYINPUT72), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT72), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n431), .A2(new_n523), .A3(new_n520), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n522), .A2(new_n524), .B1(new_n417), .B2(new_n432), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT30), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT69), .ZN(new_n527));
  INV_X1    g341(.A(new_n312), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT66), .B1(new_n423), .B2(new_n424), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n426), .B1(new_n223), .B2(new_n422), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n258), .B1(new_n531), .B2(new_n425), .ZN(new_n532));
  INV_X1    g346(.A(new_n431), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n528), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n327), .A2(new_n431), .A3(new_n520), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT30), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n527), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n312), .B1(new_n430), .B2(new_n431), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n327), .A2(new_n431), .A3(new_n520), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n527), .B(new_n537), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n526), .B(new_n373), .C1(new_n538), .C2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n373), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n525), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n252), .A2(new_n253), .A3(G210), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n546), .B(KEYINPUT27), .Z(new_n547));
  XOR2_X1   g361(.A(KEYINPUT26), .B(G101), .Z(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n543), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT31), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT31), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n543), .A2(new_n552), .A3(new_n545), .A4(new_n549), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n536), .A2(new_n373), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n522), .A2(new_n524), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n417), .A2(new_n432), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n557), .A2(KEYINPUT28), .A3(new_n373), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT28), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(new_n525), .B2(new_n544), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n554), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n549), .B(KEYINPUT73), .Z(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n551), .A2(new_n553), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(G472), .A2(G902), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT32), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT32), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n564), .A2(new_n568), .A3(new_n565), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n557), .A2(new_n373), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(new_n558), .B2(new_n560), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n549), .A2(KEYINPUT29), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n543), .A2(new_n545), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(new_n549), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT29), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n561), .B2(new_n562), .ZN(new_n577));
  OAI221_X1 g391(.A(new_n238), .B1(new_n572), .B2(new_n573), .C1(new_n575), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G472), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n517), .B1(new_n570), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n474), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(G101), .ZN(G3));
  INV_X1    g396(.A(new_n566), .ZN(new_n583));
  INV_X1    g397(.A(G472), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(new_n564), .B2(new_n238), .ZN(new_n585));
  OR2_X1    g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n401), .A2(new_n402), .ZN(new_n587));
  INV_X1    g401(.A(new_n390), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n404), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n187), .B1(new_n589), .B2(new_n409), .ZN(new_n590));
  NOR4_X1   g404(.A1(new_n586), .A2(new_n590), .A3(new_n473), .A4(new_n517), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n230), .A2(new_n232), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT96), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n212), .B2(new_n225), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT33), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n230), .A2(new_n232), .A3(new_n594), .A4(KEYINPUT33), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G478), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n234), .A2(new_n238), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n233), .B2(new_n234), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n289), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(new_n299), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n591), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G104), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G6));
  INV_X1    g421(.A(new_n289), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n237), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n299), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n591), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT35), .B(G107), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G9));
  OR2_X1    g427(.A1(new_n501), .A2(KEYINPUT36), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n497), .B(new_n614), .Z(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n515), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n510), .A2(KEYINPUT79), .A3(new_n511), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n507), .A2(new_n508), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n513), .A2(KEYINPUT98), .A3(new_n616), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n586), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n474), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT37), .B(G110), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G12));
  AOI21_X1  g441(.A(new_n473), .B1(new_n570), .B2(new_n579), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n590), .A2(new_n623), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n292), .B1(new_n296), .B2(G900), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n631), .B(KEYINPUT99), .Z(new_n632));
  NOR2_X1   g446(.A1(new_n609), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G128), .ZN(G30));
  XOR2_X1   g449(.A(new_n632), .B(KEYINPUT39), .Z(new_n636));
  NAND3_X1  g450(.A1(new_n468), .A2(new_n472), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT40), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n407), .A2(new_n409), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT38), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n571), .A2(new_n545), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n584), .B1(new_n641), .B2(new_n562), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n550), .A2(new_n642), .B1(G472), .B2(G902), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n643), .B(KEYINPUT100), .Z(new_n644));
  NAND2_X1  g458(.A1(new_n570), .A2(new_n644), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n509), .A2(new_n512), .B1(new_n515), .B2(new_n615), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n237), .A2(new_n289), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n645), .A2(new_n187), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  OR3_X1    g462(.A1(new_n638), .A2(new_n640), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G143), .ZN(G45));
  INV_X1    g464(.A(new_n632), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n599), .A2(new_n289), .A3(new_n601), .A4(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n630), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G146), .ZN(G48));
  OAI21_X1  g469(.A(new_n238), .B1(new_n457), .B2(new_n461), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(G469), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n657), .A2(new_n472), .A3(new_n462), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n590), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n580), .A2(new_n659), .A3(new_n603), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT41), .B(G113), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G15));
  NAND3_X1  g476(.A1(new_n580), .A2(new_n659), .A3(new_n610), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G116), .ZN(G18));
  NAND2_X1  g478(.A1(new_n570), .A2(new_n579), .ZN(new_n665));
  INV_X1    g479(.A(new_n658), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n629), .A2(new_n665), .A3(new_n300), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G119), .ZN(G21));
  OAI211_X1 g482(.A(new_n187), .B(new_n647), .C1(new_n589), .C2(new_n409), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n565), .B(KEYINPUT101), .Z(new_n671));
  INV_X1    g485(.A(new_n553), .ZN(new_n672));
  AOI22_X1  g486(.A1(new_n550), .A2(KEYINPUT31), .B1(new_n572), .B2(new_n562), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n672), .B1(new_n673), .B2(KEYINPUT102), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n550), .A2(KEYINPUT31), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n572), .A2(new_n562), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n671), .B1(new_n674), .B2(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n679), .A2(new_n517), .A3(new_n585), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n670), .A2(new_n680), .A3(new_n298), .A4(new_n666), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G122), .ZN(G24));
  NOR4_X1   g496(.A1(new_n679), .A2(new_n585), .A3(new_n646), .A4(new_n652), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n659), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G125), .ZN(G27));
  NAND2_X1  g499(.A1(new_n403), .A2(new_n404), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n686), .B(new_n187), .C1(new_n406), .C2(new_n403), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT106), .ZN(new_n688));
  INV_X1    g502(.A(new_n407), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(new_n690), .A3(new_n187), .A4(new_n686), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n466), .A2(KEYINPUT103), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n459), .A2(new_n694), .A3(new_n452), .A4(new_n453), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n693), .A2(G469), .A3(new_n465), .A4(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT104), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n443), .A2(new_n444), .A3(new_n415), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n698), .A2(new_n694), .B1(new_n415), .B2(new_n464), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n699), .A2(new_n700), .A3(G469), .A4(new_n693), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n462), .A2(new_n463), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n702), .A2(KEYINPUT105), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n705));
  INV_X1    g519(.A(new_n703), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n697), .A2(new_n701), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n472), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n692), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n710), .A2(new_n580), .A3(new_n653), .A4(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT105), .B1(new_n702), .B2(new_n703), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n706), .A2(new_n705), .A3(new_n707), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n471), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(new_n580), .A3(new_n691), .A4(new_n688), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n711), .B1(new_n717), .B2(new_n652), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G131), .ZN(G33));
  AND2_X1   g534(.A1(new_n688), .A2(new_n691), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n721), .A2(new_n580), .A3(new_n633), .A4(new_n716), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G134), .ZN(G36));
  NAND3_X1  g537(.A1(new_n699), .A2(KEYINPUT45), .A3(new_n693), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n411), .B1(new_n467), .B2(new_n725), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n724), .A2(new_n726), .B1(G469), .B2(G902), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n727), .A2(KEYINPUT46), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n462), .B1(new_n727), .B2(KEYINPUT46), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n472), .B(new_n636), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n234), .B1(new_n596), .B2(new_n597), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n233), .A2(new_n234), .ZN(new_n732));
  INV_X1    g546(.A(new_n600), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR4_X1   g548(.A1(new_n731), .A2(new_n734), .A3(new_n289), .A4(KEYINPUT43), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n289), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n608), .A2(KEYINPUT108), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(new_n599), .A3(new_n601), .A4(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n735), .B1(new_n739), .B2(KEYINPUT43), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n586), .A3(new_n619), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n721), .ZN(new_n744));
  OR3_X1    g558(.A1(new_n741), .A2(KEYINPUT109), .A3(new_n742), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT109), .B1(new_n741), .B2(new_n742), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n730), .B1(new_n747), .B2(KEYINPUT110), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n748), .B1(KEYINPUT110), .B2(new_n747), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT111), .B(G137), .Z(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G39));
  OAI21_X1  g565(.A(new_n472), .B1(new_n728), .B2(new_n729), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT47), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n653), .A2(new_n517), .ZN(new_n754));
  OR4_X1    g568(.A1(new_n665), .A2(new_n753), .A3(new_n692), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G140), .ZN(G42));
  INV_X1    g570(.A(new_n187), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n739), .A2(new_n471), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n517), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n657), .A2(new_n462), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n758), .B(new_n759), .C1(new_n760), .C2(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(KEYINPUT112), .Z(new_n764));
  AOI21_X1  g578(.A(new_n645), .B1(new_n760), .B2(new_n762), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n640), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n640), .A2(new_n757), .A3(new_n666), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n740), .A2(new_n291), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n680), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT50), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n692), .A2(new_n658), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n768), .ZN(new_n773));
  OR4_X1    g587(.A1(new_n585), .A2(new_n773), .A3(new_n646), .A4(new_n679), .ZN(new_n774));
  INV_X1    g588(.A(new_n772), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n570), .A2(new_n759), .A3(new_n291), .A4(new_n644), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n777), .B(new_n608), .C1(new_n731), .C2(new_n734), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n771), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n753), .B1(new_n472), .B2(new_n761), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n769), .A2(new_n692), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n782), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n780), .A2(KEYINPUT51), .A3(new_n786), .ZN(new_n787));
  XOR2_X1   g601(.A(KEYINPUT118), .B(KEYINPUT51), .Z(new_n788));
  AND2_X1   g602(.A1(new_n781), .A2(new_n784), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n788), .B1(new_n779), .B2(new_n789), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n769), .A2(new_n590), .A3(new_n658), .ZN(new_n791));
  INV_X1    g605(.A(new_n602), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n290), .B(new_n791), .C1(new_n792), .C2(new_n777), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT120), .ZN(new_n794));
  INV_X1    g608(.A(new_n580), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n773), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT48), .Z(new_n797));
  NAND4_X1  g611(.A1(new_n787), .A2(new_n790), .A3(new_n794), .A4(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n716), .A2(new_n683), .A3(new_n691), .A4(new_n688), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n639), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(KEYINPUT113), .A3(new_n187), .A4(new_n603), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n586), .A2(new_n517), .A3(new_n473), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n299), .B1(new_n602), .B2(new_n609), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n805), .B(new_n187), .C1(new_n407), .C2(new_n409), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n803), .B(new_n804), .C1(new_n807), .C2(KEYINPUT113), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n474), .B1(new_n624), .B2(new_n580), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n623), .A2(new_n237), .A3(new_n289), .A4(new_n632), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n628), .A3(new_n691), .A4(new_n688), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n722), .A2(new_n808), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n801), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n628), .B(new_n629), .C1(new_n633), .C2(new_n653), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n646), .A2(new_n651), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n570), .B2(new_n644), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n714), .A2(new_n715), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n817), .A3(new_n472), .A4(new_n670), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n814), .A2(new_n818), .A3(new_n684), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT52), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n814), .A2(new_n818), .A3(new_n821), .A4(new_n684), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n660), .A2(new_n667), .A3(new_n681), .A4(new_n663), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n713), .B2(new_n718), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n813), .A2(new_n823), .A3(KEYINPUT53), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n824), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n719), .A2(new_n829), .A3(new_n820), .A4(new_n822), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(KEYINPUT115), .A3(KEYINPUT53), .A4(new_n813), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n825), .A2(new_n820), .A3(new_n822), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n801), .A2(new_n812), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n828), .A2(new_n831), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT54), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n825), .A2(KEYINPUT116), .A3(new_n820), .A4(new_n822), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n838), .B(KEYINPUT53), .C1(new_n833), .C2(new_n834), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n830), .B(new_n813), .C1(KEYINPUT116), .C2(new_n832), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT117), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n837), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n798), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(G952), .A2(G953), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n766), .B1(new_n848), .B2(new_n849), .ZN(G75));
  NOR2_X1   g664(.A1(new_n253), .A2(G952), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n839), .A2(new_n840), .A3(G210), .A4(G902), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n394), .A2(new_n396), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(new_n398), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT55), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n851), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n839), .A2(new_n840), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(G902), .A3(new_n405), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n857), .A2(KEYINPUT56), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n860), .A2(KEYINPUT121), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT121), .B1(new_n860), .B2(new_n861), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(G51));
  XOR2_X1   g679(.A(new_n463), .B(KEYINPUT57), .Z(new_n866));
  NOR2_X1   g680(.A1(new_n841), .A2(new_n842), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT54), .B1(new_n839), .B2(new_n840), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n461), .B2(new_n457), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n841), .A2(new_n238), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n724), .A3(new_n726), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n851), .B1(new_n870), .B2(new_n872), .ZN(G54));
  NAND3_X1  g687(.A1(new_n871), .A2(KEYINPUT58), .A3(G475), .ZN(new_n874));
  INV_X1    g688(.A(new_n284), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n876), .A2(new_n877), .A3(new_n851), .ZN(G60));
  INV_X1    g692(.A(new_n598), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n600), .B(KEYINPUT59), .Z(new_n880));
  OAI211_X1 g694(.A(new_n879), .B(new_n880), .C1(new_n867), .C2(new_n868), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(G952), .B2(new_n253), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n845), .A2(new_n847), .A3(new_n880), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n882), .B1(new_n883), .B2(new_n598), .ZN(G63));
  NAND2_X1  g698(.A1(G217), .A2(G902), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT60), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n839), .A2(new_n840), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n502), .A2(new_n503), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n851), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n859), .A2(new_n615), .A3(new_n887), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT122), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n892), .B(new_n893), .ZN(G66));
  OAI21_X1  g708(.A(G953), .B1(new_n293), .B2(new_n330), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT123), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n829), .A2(new_n808), .A3(new_n809), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(new_n253), .ZN(new_n898));
  INV_X1    g712(.A(G898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n855), .B1(new_n899), .B2(G953), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n898), .B(new_n900), .ZN(G69));
  AOI21_X1  g715(.A(new_n253), .B1(G227), .B2(G900), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n814), .A2(new_n684), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n649), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n602), .A2(new_n609), .ZN(new_n908));
  OR4_X1    g722(.A1(new_n795), .A2(new_n692), .A3(new_n637), .A4(new_n908), .ZN(new_n909));
  AND4_X1   g723(.A1(new_n749), .A2(new_n907), .A3(new_n755), .A4(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n538), .A2(new_n542), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(KEYINPUT30), .B2(new_n525), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n281), .B(KEYINPUT124), .Z(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n910), .A2(G953), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(G900), .A2(G953), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n580), .A2(new_n670), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n722), .B1(new_n730), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n903), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n749), .A2(new_n755), .A3(new_n719), .A4(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n916), .B1(new_n920), .B2(G953), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n902), .B(new_n915), .C1(new_n921), .C2(new_n914), .ZN(new_n922));
  NAND2_X1  g736(.A1(G227), .A2(G900), .ZN(new_n923));
  AND4_X1   g737(.A1(G953), .A2(new_n921), .A3(new_n923), .A4(new_n914), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n924), .ZN(G72));
  NAND2_X1  g739(.A1(G472), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT63), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT125), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n920), .B2(new_n897), .ZN(new_n929));
  INV_X1    g743(.A(new_n574), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(new_n549), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n851), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n749), .A2(new_n907), .A3(new_n755), .A4(new_n909), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n928), .B1(new_n933), .B2(new_n897), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n934), .A2(new_n930), .A3(new_n549), .ZN(new_n935));
  INV_X1    g749(.A(new_n575), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n927), .B1(new_n936), .B2(new_n550), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n836), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n932), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT126), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n932), .A2(new_n935), .A3(new_n941), .A4(new_n938), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(G57));
endmodule


