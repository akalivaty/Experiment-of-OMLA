//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  AOI21_X1  g006(.A(G1gat), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT93), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n206), .B(new_n209), .C1(new_n207), .C2(G1gat), .ZN(new_n212));
  INV_X1    g011(.A(G8gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n211), .B(new_n212), .C1(KEYINPUT94), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(KEYINPUT94), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(new_n216), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT21), .ZN(new_n220));
  XNOR2_X1  g019(.A(G57gat), .B(G64gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT98), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G71gat), .A2(G78gat), .ZN(new_n224));
  OR2_X1    g023(.A1(G71gat), .A2(G78gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT9), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n224), .B(new_n225), .C1(new_n221), .C2(new_n226), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n219), .B1(new_n220), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(G183gat), .ZN(new_n232));
  INV_X1    g031(.A(G231gat), .ZN(new_n233));
  INV_X1    g032(.A(G233gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G183gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n231), .B(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(G231gat), .A3(G233gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n205), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n230), .A2(new_n220), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n241), .B(new_n242), .Z(new_n243));
  NAND3_X1  g042(.A1(new_n235), .A2(new_n238), .A3(new_n205), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n243), .ZN(new_n246));
  INV_X1    g045(.A(new_n244), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n246), .B1(new_n247), .B2(new_n239), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(G190gat), .B(G218gat), .Z(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT99), .ZN(new_n252));
  XOR2_X1   g051(.A(G134gat), .B(G162gat), .Z(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n251), .A2(KEYINPUT99), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT14), .ZN(new_n257));
  INV_X1    g056(.A(G29gat), .ZN(new_n258));
  INV_X1    g057(.A(G36gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n260), .A2(new_n261), .B1(G29gat), .B2(G36gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(G43gat), .B(G50gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n262), .B1(KEYINPUT15), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(KEYINPUT15), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n264), .B(new_n265), .Z(new_n266));
  INV_X1    g065(.A(KEYINPUT17), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n264), .B(new_n265), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT17), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G85gat), .A2(G92gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT7), .ZN(new_n273));
  INV_X1    g072(.A(G99gat), .ZN(new_n274));
  INV_X1    g073(.A(G106gat), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT8), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n273), .B(new_n276), .C1(G85gat), .C2(G92gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(G99gat), .B(G106gat), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n277), .B(new_n278), .Z(new_n279));
  NAND2_X1  g078(.A1(new_n271), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n277), .B(new_n278), .ZN(new_n281));
  AND2_X1   g080(.A1(G232gat), .A2(G233gat), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n266), .A2(new_n281), .B1(KEYINPUT41), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n256), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n282), .A2(KEYINPUT41), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n284), .A2(new_n286), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n255), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n284), .A2(new_n286), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(new_n287), .A3(new_n254), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G230gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n294), .A2(new_n234), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n230), .ZN(new_n296));
  INV_X1    g095(.A(new_n230), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n281), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT10), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n281), .A3(KEYINPUT10), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n295), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI211_X1 g101(.A(new_n294), .B(new_n234), .C1(new_n296), .C2(new_n298), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n304), .A2(KEYINPUT100), .ZN(new_n305));
  XNOR2_X1  g104(.A(G120gat), .B(G148gat), .ZN(new_n306));
  INV_X1    g105(.A(G176gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G204gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n305), .B(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n249), .A2(new_n293), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT101), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT101), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n249), .A2(new_n314), .A3(new_n293), .A4(new_n311), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n217), .A2(new_n218), .A3(new_n266), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT96), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n219), .A2(new_n270), .A3(new_n268), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT95), .ZN(new_n321));
  NAND2_X1  g120(.A1(G229gat), .A2(G233gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT95), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n271), .A2(new_n323), .A3(new_n219), .ZN(new_n324));
  AND4_X1   g123(.A1(new_n319), .A2(new_n321), .A3(new_n322), .A4(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT18), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n219), .A2(new_n269), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n322), .B(KEYINPUT13), .Z(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n319), .A2(new_n321), .A3(new_n324), .A4(new_n322), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT18), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n326), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT97), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n330), .B(new_n335), .C1(new_n332), .C2(new_n331), .ZN(new_n336));
  XNOR2_X1  g135(.A(G169gat), .B(G197gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT92), .ZN(new_n338));
  XOR2_X1   g137(.A(G113gat), .B(G141gat), .Z(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT12), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n334), .A2(new_n336), .A3(new_n344), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n325), .A2(KEYINPUT18), .B1(new_n328), .B2(new_n329), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n346), .B(new_n333), .C1(new_n335), .C2(new_n343), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT90), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT32), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT33), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n352));
  INV_X1    g151(.A(G169gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n353), .A3(new_n307), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n354), .A2(new_n355), .B1(G169gat), .B2(G176gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n236), .A2(KEYINPUT67), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT67), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G183gat), .ZN(new_n359));
  AOI21_X1  g158(.A(G190gat), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT66), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT24), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(G183gat), .B(G190gat), .C1(KEYINPUT66), .C2(KEYINPUT24), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n356), .B(KEYINPUT25), .C1(new_n360), .C2(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(G183gat), .A2(G190gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n361), .A2(KEYINPUT24), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n363), .A2(G183gat), .A3(G190gat), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT65), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI211_X1 g172(.A(KEYINPUT65), .B(new_n368), .C1(new_n369), .C2(new_n370), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n354), .A2(new_n355), .ZN(new_n375));
  NAND2_X1  g174(.A1(G169gat), .A2(G176gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n373), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n367), .B1(new_n378), .B2(KEYINPUT25), .ZN(new_n379));
  INV_X1    g178(.A(G134gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G127gat), .ZN(new_n381));
  INV_X1    g180(.A(G127gat), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT1), .B1(new_n382), .B2(G134gat), .ZN(new_n383));
  INV_X1    g182(.A(G120gat), .ZN(new_n384));
  INV_X1    g183(.A(G113gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT71), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT71), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G113gat), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n384), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n385), .A2(G120gat), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n381), .B(new_n383), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT1), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n384), .A2(G113gat), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n382), .A2(KEYINPUT70), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT70), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G127gat), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n380), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT69), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(new_n382), .B2(G134gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n380), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n394), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n391), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT27), .B(G183gat), .ZN(new_n406));
  INV_X1    g205(.A(G190gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(KEYINPUT28), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n357), .A2(new_n359), .A3(KEYINPUT27), .ZN(new_n409));
  OR2_X1    g208(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n410));
  AOI21_X1  g209(.A(G190gat), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n408), .B1(new_n411), .B2(KEYINPUT28), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT68), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n353), .A2(new_n307), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT26), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n361), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT26), .B1(new_n353), .B2(new_n307), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n416), .B1(new_n376), .B2(new_n417), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n412), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n413), .B1(new_n412), .B2(new_n418), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n379), .B(new_n405), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT72), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n412), .A2(new_n418), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT68), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n412), .A2(new_n413), .A3(new_n418), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n427), .A2(KEYINPUT72), .A3(new_n405), .A4(new_n379), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n379), .B1(new_n419), .B2(new_n420), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n404), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n423), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT73), .ZN(new_n432));
  NAND2_X1  g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT64), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n432), .B1(new_n431), .B2(new_n434), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n351), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G15gat), .B(G43gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(G71gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(new_n274), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n431), .A2(new_n434), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT73), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n350), .B1(new_n440), .B2(KEYINPUT33), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT74), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(KEYINPUT74), .B(new_n446), .C1(new_n435), .C2(new_n436), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n441), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n431), .A2(KEYINPUT34), .A3(new_n434), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n423), .A2(new_n428), .A3(new_n430), .A4(new_n433), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n453), .A2(KEYINPUT75), .A3(KEYINPUT34), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT75), .B1(new_n453), .B2(KEYINPUT34), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n446), .B1(new_n435), .B2(new_n436), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT74), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n448), .ZN(new_n461));
  INV_X1    g260(.A(new_n456), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n441), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G197gat), .B(G204gat), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT22), .ZN(new_n465));
  INV_X1    g264(.A(G218gat), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n465), .B1(new_n203), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(G211gat), .B(G218gat), .Z(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT76), .ZN(new_n471));
  INV_X1    g270(.A(G155gat), .ZN(new_n472));
  INV_X1    g271(.A(G162gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(G155gat), .A2(G162gat), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT80), .B(KEYINPUT2), .ZN(new_n477));
  INV_X1    g276(.A(G141gat), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(G148gat), .ZN(new_n479));
  INV_X1    g278(.A(G148gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(G141gat), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n477), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT81), .B1(new_n480), .B2(G141gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(new_n478), .A3(G148gat), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n483), .B(new_n485), .C1(new_n478), .C2(G148gat), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n475), .B1(new_n474), .B2(KEYINPUT2), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n476), .A2(new_n482), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT3), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n471), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT29), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n470), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n488), .B1(new_n496), .B2(new_n489), .ZN(new_n497));
  OAI211_X1 g296(.A(G228gat), .B(G233gat), .C1(new_n494), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(G228gat), .A2(G233gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n492), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT3), .B1(new_n470), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n499), .B1(new_n501), .B2(new_n488), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n494), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G22gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n498), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT76), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n470), .B(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(new_n491), .B2(new_n492), .ZN(new_n508));
  INV_X1    g307(.A(new_n497), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n499), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n502), .ZN(new_n511));
  OAI21_X1  g310(.A(G22gat), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n505), .A2(new_n512), .A3(KEYINPUT88), .ZN(new_n513));
  XOR2_X1   g312(.A(G78gat), .B(G106gat), .Z(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n514), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n505), .A2(new_n512), .A3(KEYINPUT88), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT31), .B(G50gat), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n515), .A2(new_n519), .A3(new_n517), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n457), .A2(new_n463), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n525));
  NAND2_X1  g324(.A1(G226gat), .A2(G233gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n429), .A2(new_n500), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n526), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n379), .A2(new_n424), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n471), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT29), .B1(new_n379), .B2(new_n424), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT78), .B1(new_n531), .B2(new_n528), .ZN(new_n532));
  INV_X1    g331(.A(new_n367), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n371), .A2(new_n372), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n371), .A2(new_n372), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n356), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n533), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n424), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n495), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT78), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(new_n526), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n429), .A2(new_n528), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n532), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n530), .B1(new_n544), .B2(new_n471), .ZN(new_n545));
  XOR2_X1   g344(.A(G8gat), .B(G36gat), .Z(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(G64gat), .ZN(new_n547));
  INV_X1    g346(.A(G92gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n525), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n545), .A2(new_n549), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT79), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n544), .A2(new_n471), .ZN(new_n553));
  INV_X1    g352(.A(new_n530), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n552), .B1(new_n555), .B2(KEYINPUT30), .ZN(new_n556));
  NOR4_X1   g355(.A1(new_n545), .A2(KEYINPUT79), .A3(new_n525), .A4(new_n549), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n550), .B(new_n551), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT35), .ZN(new_n560));
  NAND2_X1  g359(.A1(G225gat), .A2(G233gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n486), .A2(new_n487), .ZN(new_n562));
  XOR2_X1   g361(.A(KEYINPUT80), .B(KEYINPUT2), .Z(new_n563));
  XNOR2_X1  g362(.A(G141gat), .B(G148gat), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n476), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT3), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT82), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n391), .A2(new_n403), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n568), .B1(new_n391), .B2(new_n403), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n567), .B(new_n490), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT83), .B(KEYINPUT4), .Z(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n404), .B2(new_n566), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT84), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g374(.A(KEYINPUT84), .B(new_n572), .C1(new_n404), .C2(new_n566), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT85), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n578), .B1(new_n404), .B2(new_n566), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n488), .A2(KEYINPUT85), .A3(new_n403), .A4(new_n391), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT4), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n561), .B(new_n571), .C1(new_n577), .C2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT5), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(new_n579), .A3(new_n580), .ZN(new_n585));
  INV_X1    g384(.A(new_n561), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n583), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OR3_X1    g386(.A1(new_n404), .A2(new_n566), .A3(new_n572), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n579), .A2(KEYINPUT4), .A3(new_n580), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n569), .A2(new_n570), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n490), .A2(new_n567), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n588), .A2(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n586), .A2(KEYINPUT5), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n582), .A2(new_n587), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT0), .B(G57gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G85gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G1gat), .B(G29gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  AOI21_X1  g397(.A(KEYINPUT6), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n587), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n592), .A2(new_n593), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n598), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n594), .A2(new_n598), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT6), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n559), .A2(new_n560), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n349), .B1(new_n524), .B2(new_n609), .ZN(new_n610));
  AOI221_X4 g409(.A(new_n456), .B1(new_n437), .B2(new_n440), .C1(new_n460), .C2(new_n448), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n462), .B1(new_n461), .B2(new_n441), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n608), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n558), .A2(new_n614), .A3(KEYINPUT35), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n613), .A2(KEYINPUT90), .A3(new_n523), .A4(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT87), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n604), .B1(new_n599), .B2(KEYINPUT86), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT86), .ZN(new_n619));
  AOI211_X1 g418(.A(new_n619), .B(KEYINPUT6), .C1(new_n594), .C2(new_n598), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n617), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n600), .A2(new_n598), .A3(new_n601), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n619), .B1(new_n622), .B2(KEYINPUT6), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT6), .ZN(new_n624));
  OAI211_X1 g423(.A(KEYINPUT86), .B(new_n624), .C1(new_n602), .C2(new_n603), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n623), .A2(KEYINPUT87), .A3(new_n604), .A4(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n607), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n559), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(new_n613), .A3(new_n523), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n610), .A2(new_n616), .B1(new_n629), .B2(KEYINPUT35), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n585), .A2(new_n586), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n631), .B(KEYINPUT39), .C1(new_n561), .C2(new_n592), .ZN(new_n632));
  OR3_X1    g431(.A1(new_n592), .A2(KEYINPUT39), .A3(new_n561), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n632), .A2(new_n633), .A3(new_n598), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT40), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n636), .A2(new_n637), .A3(new_n606), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n558), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n553), .A2(new_n554), .ZN(new_n640));
  INV_X1    g439(.A(new_n549), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT38), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n527), .A2(new_n471), .A3(new_n529), .ZN(new_n645));
  OAI211_X1 g444(.A(KEYINPUT37), .B(new_n645), .C1(new_n544), .C2(new_n471), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT89), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT37), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n640), .B2(new_n648), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n545), .A2(KEYINPUT89), .A3(KEYINPUT37), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n642), .B(new_n646), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n644), .B1(new_n651), .B2(new_n549), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n640), .A2(new_n647), .A3(new_n648), .ZN(new_n653));
  OAI21_X1  g452(.A(KEYINPUT89), .B1(new_n545), .B2(KEYINPUT37), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n653), .A2(new_n654), .B1(KEYINPUT37), .B2(new_n545), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n614), .B1(new_n655), .B2(new_n642), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n639), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n523), .ZN(new_n658));
  INV_X1    g457(.A(new_n523), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(new_n627), .A3(new_n559), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT36), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(new_n611), .B2(new_n612), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n457), .A2(KEYINPUT36), .A3(new_n463), .ZN(new_n663));
  AOI22_X1  g462(.A1(new_n658), .A2(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n316), .B(new_n348), .C1(new_n630), .C2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n627), .B(KEYINPUT102), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n667), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g467(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n665), .A2(new_n559), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(KEYINPUT42), .A3(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n672), .A2(KEYINPUT103), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT42), .B1(new_n670), .B2(new_n671), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n665), .A2(new_n559), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n213), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n672), .A2(KEYINPUT103), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n673), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n673), .A2(new_n677), .A3(KEYINPUT104), .A4(new_n678), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(G1325gat));
  INV_X1    g482(.A(new_n613), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n665), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(G15gat), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n611), .A2(new_n612), .A3(new_n661), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT36), .B1(new_n457), .B2(new_n463), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n662), .A2(KEYINPUT105), .A3(new_n663), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n665), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n686), .B1(G15gat), .B2(new_n694), .ZN(G1326gat));
  NOR2_X1   g494(.A1(new_n665), .A2(new_n523), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT43), .B(G22gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  NOR2_X1   g497(.A1(new_n630), .A2(new_n664), .ZN(new_n699));
  INV_X1    g498(.A(new_n249), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(new_n311), .A3(new_n348), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n699), .A2(new_n293), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n666), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n258), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT45), .ZN(new_n705));
  INV_X1    g504(.A(new_n293), .ZN(new_n706));
  OAI22_X1  g505(.A1(new_n649), .A2(new_n650), .B1(new_n648), .B2(new_n640), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n608), .B1(new_n707), .B2(KEYINPUT38), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n646), .A2(new_n642), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n653), .B2(new_n654), .ZN(new_n710));
  OAI22_X1  g509(.A1(new_n710), .A2(new_n641), .B1(new_n640), .B2(new_n643), .ZN(new_n711));
  AOI22_X1  g510(.A1(new_n708), .A2(new_n711), .B1(new_n558), .B2(new_n638), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n660), .B1(new_n712), .B2(new_n659), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n690), .A2(new_n713), .A3(new_n691), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n706), .B1(new_n714), .B2(new_n630), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718));
  OAI211_X1 g517(.A(KEYINPUT44), .B(new_n706), .C1(new_n630), .C2(new_n664), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n701), .B(KEYINPUT106), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n717), .A2(new_n718), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n610), .A2(new_n616), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n629), .A2(KEYINPUT35), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n690), .A2(new_n713), .A3(new_n691), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n293), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n719), .B(new_n720), .C1(new_n726), .C2(KEYINPUT44), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT107), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n666), .B1(new_n721), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n705), .B1(new_n258), .B2(new_n729), .ZN(G1328gat));
  AND2_X1   g529(.A1(new_n727), .A2(KEYINPUT107), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n727), .A2(KEYINPUT107), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n558), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G36gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n702), .A2(new_n259), .A3(new_n558), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(KEYINPUT108), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n736), .A2(KEYINPUT108), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n735), .A2(new_n737), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n734), .A2(KEYINPUT109), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n559), .B1(new_n721), .B2(new_n728), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n739), .B(new_n740), .C1(new_n742), .C2(new_n259), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(new_n745), .ZN(G1329gat));
  INV_X1    g545(.A(new_n702), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n747), .A2(G43gat), .A3(new_n684), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G43gat), .B1(new_n727), .B2(new_n693), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(KEYINPUT47), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n692), .B1(new_n731), .B2(new_n732), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n748), .B1(new_n752), .B2(G43gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n753), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g553(.A1(new_n747), .A2(G50gat), .A3(new_n523), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G50gat), .B1(new_n727), .B2(new_n523), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n756), .A2(KEYINPUT48), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n659), .B1(new_n731), .B2(new_n732), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n755), .B1(new_n759), .B2(G50gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n760), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g560(.A(new_n348), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(new_n249), .A3(new_n293), .ZN(new_n763));
  AOI211_X1 g562(.A(new_n311), .B(new_n763), .C1(new_n724), .C2(new_n725), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n703), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n764), .A2(new_n558), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT110), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1333gat));
  OR2_X1    g570(.A1(new_n684), .A2(KEYINPUT111), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n684), .A2(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(G71gat), .B1(new_n764), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n692), .A2(G71gat), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n764), .B2(new_n777), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n659), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G78gat), .ZN(G1335gat));
  INV_X1    g580(.A(new_n311), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n700), .A2(new_n762), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n706), .B(new_n784), .C1(new_n714), .C2(new_n630), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT51), .B1(new_n726), .B2(new_n784), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n782), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(G85gat), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(new_n791), .A3(new_n703), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n784), .A2(new_n782), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT112), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n794), .B(new_n719), .C1(KEYINPUT44), .C2(new_n726), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(new_n666), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT113), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n792), .B1(new_n797), .B2(new_n791), .ZN(G1336gat));
  OAI21_X1  g597(.A(G92gat), .B1(new_n795), .B2(new_n559), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n558), .A2(new_n548), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n799), .B(new_n800), .C1(new_n789), .C2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n785), .B2(KEYINPUT114), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT114), .B1(new_n803), .B2(KEYINPUT51), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n804), .A2(new_n786), .B1(new_n785), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(new_n548), .A3(new_n782), .A4(new_n558), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n808), .A2(new_n799), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n802), .B1(new_n809), .B2(new_n800), .ZN(G1337gat));
  NAND3_X1  g609(.A1(new_n790), .A2(new_n274), .A3(new_n613), .ZN(new_n811));
  OAI21_X1  g610(.A(G99gat), .B1(new_n795), .B2(new_n693), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1338gat));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n804), .A2(new_n786), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n785), .A2(new_n806), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n523), .A2(G106gat), .A3(new_n311), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G106gat), .B1(new_n795), .B2(new_n523), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n815), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n818), .B1(new_n787), .B2(new_n788), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n815), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n814), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n717), .A2(new_n659), .A3(new_n719), .A4(new_n794), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n807), .A2(new_n818), .B1(G106gat), .B2(new_n826), .ZN(new_n827));
  OAI211_X1 g626(.A(KEYINPUT116), .B(new_n823), .C1(new_n827), .C2(new_n815), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(G1339gat));
  NOR2_X1   g628(.A1(new_n763), .A2(new_n782), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n831));
  INV_X1    g630(.A(new_n310), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n302), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n300), .A2(new_n301), .A3(new_n295), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT54), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n302), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n831), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n836), .A2(new_n302), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n841), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(new_n834), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n304), .A2(new_n832), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n839), .A2(new_n840), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n347), .B2(new_n345), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n326), .A2(new_n330), .A3(new_n343), .A4(new_n333), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n324), .A2(new_n321), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n322), .B1(new_n847), .B2(new_n319), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n328), .A2(new_n329), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n342), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n311), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n293), .B1(new_n845), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n844), .ZN(new_n854));
  INV_X1    g653(.A(new_n851), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n855), .A3(new_n706), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n844), .A2(new_n851), .A3(new_n293), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT118), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n853), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n830), .B1(new_n861), .B2(new_n700), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n558), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n666), .A2(new_n524), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(new_n762), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n386), .A2(new_n388), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(new_n385), .B2(new_n866), .ZN(G1340gat));
  NOR2_X1   g668(.A1(new_n865), .A2(new_n311), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(new_n384), .ZN(G1341gat));
  NOR2_X1   g670(.A1(new_n865), .A2(new_n700), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n395), .A2(new_n397), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n872), .B(new_n873), .ZN(G1342gat));
  NOR2_X1   g673(.A1(new_n865), .A2(new_n293), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n380), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n877), .B(new_n878), .C1(new_n380), .C2(new_n875), .ZN(G1343gat));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n844), .A2(new_n851), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT118), .B1(new_n881), .B2(new_n706), .ZN(new_n882));
  NOR4_X1   g681(.A1(new_n844), .A2(new_n851), .A3(new_n293), .A4(new_n857), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n840), .A2(KEYINPUT119), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n837), .A2(new_n887), .A3(new_n838), .ZN(new_n888));
  AND4_X1   g687(.A1(new_n843), .A2(new_n839), .A3(new_n842), .A4(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n348), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n852), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n706), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n700), .B1(new_n885), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n893), .B1(new_n782), .B2(new_n763), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n880), .B1(new_n894), .B2(new_n659), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n249), .B1(new_n884), .B2(new_n853), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n659), .B1(new_n896), .B2(new_n830), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(KEYINPUT57), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n692), .A2(new_n666), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n559), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n895), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n478), .B1(new_n901), .B2(new_n348), .ZN(new_n902));
  INV_X1    g701(.A(new_n897), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n559), .A3(new_n899), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n348), .A2(new_n478), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n905), .B(KEYINPUT120), .Z(new_n906));
  NOR2_X1   g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  OR3_X1    g706(.A1(new_n902), .A2(KEYINPUT58), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT58), .B1(new_n902), .B2(new_n907), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1344gat));
  INV_X1    g709(.A(new_n904), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n480), .A3(new_n782), .ZN(new_n912));
  AOI211_X1 g711(.A(KEYINPUT59), .B(new_n480), .C1(new_n901), .C2(new_n782), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n700), .B1(new_n892), .B2(new_n859), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n313), .A2(new_n315), .A3(new_n762), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT57), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n897), .A2(KEYINPUT57), .B1(new_n916), .B2(new_n659), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n782), .ZN(new_n918));
  OAI21_X1  g717(.A(G148gat), .B1(new_n918), .B2(new_n900), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n919), .A2(KEYINPUT59), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n912), .B1(new_n913), .B2(new_n920), .ZN(G1345gat));
  NAND3_X1  g720(.A1(new_n901), .A2(G155gat), .A3(new_n249), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n472), .B1(new_n904), .B2(new_n700), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(G1346gat));
  NAND3_X1  g723(.A1(new_n911), .A2(new_n473), .A3(new_n706), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT121), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n901), .A2(new_n706), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n473), .B2(new_n927), .ZN(G1347gat));
  OAI21_X1  g727(.A(new_n666), .B1(new_n896), .B2(new_n830), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n929), .A2(new_n559), .A3(new_n524), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n353), .A3(new_n348), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n862), .A2(new_n703), .A3(new_n559), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n774), .A2(new_n659), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n348), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n932), .B1(new_n937), .B2(G169gat), .ZN(new_n938));
  AOI211_X1 g737(.A(KEYINPUT122), .B(new_n353), .C1(new_n936), .C2(new_n348), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n931), .B1(new_n938), .B2(new_n939), .ZN(G1348gat));
  NOR3_X1   g739(.A1(new_n935), .A2(new_n307), .A3(new_n311), .ZN(new_n941));
  AOI21_X1  g740(.A(G176gat), .B1(new_n930), .B2(new_n782), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(G1349gat));
  NAND4_X1  g742(.A1(new_n930), .A2(KEYINPUT123), .A3(new_n249), .A4(new_n406), .ZN(new_n944));
  INV_X1    g743(.A(new_n524), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n933), .A2(new_n249), .A3(new_n406), .A4(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT60), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n357), .A2(new_n359), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n700), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n949), .B(new_n951), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n950), .A2(KEYINPUT60), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n954), .B(new_n955), .ZN(G1350gat));
  OAI21_X1  g755(.A(G190gat), .B1(new_n935), .B2(new_n293), .ZN(new_n957));
  XOR2_X1   g756(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n957), .A2(new_n959), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n930), .A2(new_n407), .A3(new_n706), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(G1351gat));
  NOR2_X1   g762(.A1(new_n692), .A2(new_n559), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(new_n659), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n929), .B1(new_n965), .B2(KEYINPUT126), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(G197gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n968), .A2(new_n969), .A3(new_n348), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n917), .A2(new_n666), .A3(new_n964), .ZN(new_n971));
  OAI21_X1  g770(.A(G197gat), .B1(new_n971), .B2(new_n762), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1352gat));
  NAND3_X1  g772(.A1(new_n968), .A2(new_n309), .A3(new_n782), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n974), .A2(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(KEYINPUT62), .ZN(new_n976));
  NOR4_X1   g775(.A1(new_n918), .A2(new_n703), .A3(new_n559), .A4(new_n692), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n975), .B(new_n976), .C1(new_n309), .C2(new_n977), .ZN(G1353gat));
  NAND3_X1  g777(.A1(new_n968), .A2(new_n203), .A3(new_n249), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n917), .A2(new_n964), .A3(new_n666), .A4(new_n249), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n980), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT63), .B1(new_n980), .B2(G211gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n979), .B(KEYINPUT127), .C1(new_n981), .C2(new_n982), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1354gat));
  NOR3_X1   g786(.A1(new_n971), .A2(new_n466), .A3(new_n293), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n968), .A2(new_n706), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n988), .B1(new_n466), .B2(new_n989), .ZN(G1355gat));
endmodule


