//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1287, new_n1288, new_n1289, new_n1290, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G250), .B(G257), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G264), .B(G270), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT64), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n231), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n202), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n240), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G200), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n254), .A2(G223), .B1(new_n257), .B2(G77), .ZN(new_n258));
  INV_X1    g0058(.A(G222), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1698), .B1(new_n252), .B2(new_n253), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G1), .A3(G13), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(new_n268), .A3(G274), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n265), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n270), .B1(G226), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n248), .B1(new_n264), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n274), .A2(KEYINPUT70), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(KEYINPUT70), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n264), .A2(new_n273), .ZN(new_n277));
  INV_X1    g0077(.A(G190), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR4_X1   g0079(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT10), .A4(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT65), .A2(G58), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT65), .A2(G58), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT8), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n207), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OR2_X1    g0085(.A1(KEYINPUT8), .A2(G58), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n216), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n290), .A2(new_n292), .B1(new_n202), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n206), .A2(G20), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT66), .B1(new_n294), .B2(new_n292), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n294), .A2(new_n292), .A3(KEYINPUT66), .ZN(new_n299));
  OAI211_X1 g0099(.A(G50), .B(new_n296), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n295), .A2(new_n300), .A3(KEYINPUT9), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT69), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT69), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n295), .A2(new_n300), .A3(new_n303), .A4(KEYINPUT9), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT68), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n295), .A2(new_n300), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT9), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI211_X1 g0108(.A(KEYINPUT68), .B(KEYINPUT9), .C1(new_n295), .C2(new_n300), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n302), .B(new_n304), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n280), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT71), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n279), .A2(new_n274), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n313), .B(KEYINPUT10), .C1(new_n310), .C2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT9), .B1(new_n295), .B2(new_n300), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(new_n305), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n302), .A2(new_n304), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n279), .A2(new_n274), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n313), .B1(new_n321), .B2(KEYINPUT10), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n312), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  XOR2_X1   g0123(.A(KEYINPUT8), .B(G58), .Z(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(new_n288), .B1(G20), .B2(G77), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT15), .B(G87), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n284), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n292), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT67), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n294), .A2(new_n292), .ZN(new_n330));
  INV_X1    g0130(.A(G77), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n206), .B2(G20), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n330), .A2(new_n332), .B1(new_n331), .B2(new_n294), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n254), .A2(G238), .B1(new_n257), .B2(G107), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n233), .B2(new_n261), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n263), .ZN(new_n338));
  INV_X1    g0138(.A(G244), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n338), .B(new_n269), .C1(new_n339), .C2(new_n271), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G200), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n335), .B(new_n341), .C1(new_n278), .C2(new_n340), .ZN(new_n342));
  INV_X1    g0142(.A(G169), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n334), .B(new_n344), .C1(G179), .C2(new_n340), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n283), .A2(new_n286), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n293), .ZN(new_n348));
  INV_X1    g0148(.A(new_n299), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n297), .B1(new_n206), .B2(G20), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n348), .B1(new_n350), .B2(new_n347), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT7), .B1(new_n257), .B2(new_n207), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n253), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(G68), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT78), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT77), .ZN(new_n358));
  INV_X1    g0158(.A(new_n288), .ZN(new_n359));
  INV_X1    g0159(.A(G159), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT65), .B(G58), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n201), .B1(new_n363), .B2(G68), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n358), .B(new_n362), .C1(new_n364), .C2(new_n207), .ZN(new_n365));
  OAI21_X1  g0165(.A(G68), .B1(new_n281), .B2(new_n282), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n207), .B1(new_n366), .B2(new_n213), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT77), .B1(new_n367), .B2(new_n361), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n252), .A2(new_n207), .A3(new_n253), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT7), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n354), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT78), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n373), .A3(G68), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n357), .A2(new_n365), .A3(new_n368), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n368), .A2(new_n365), .A3(KEYINPUT16), .A4(new_n356), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n378), .A2(new_n292), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n352), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n269), .B1(new_n233), .B2(new_n271), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n254), .A2(G226), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n260), .A2(G223), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G33), .A2(G87), .ZN(new_n384));
  XOR2_X1   g0184(.A(new_n384), .B(KEYINPUT79), .Z(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n381), .B1(new_n386), .B2(new_n263), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G179), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n343), .B2(new_n387), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT18), .B1(new_n380), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n373), .B1(new_n372), .B2(G68), .ZN(new_n392));
  AOI211_X1 g0192(.A(KEYINPUT78), .B(new_n242), .C1(new_n371), .C2(new_n354), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n368), .A2(new_n365), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT16), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n378), .A2(new_n292), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n351), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n399), .A3(new_n389), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n386), .A2(new_n263), .ZN(new_n401));
  INV_X1    g0201(.A(new_n381), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n278), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G200), .B2(new_n387), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n380), .A2(KEYINPUT17), .A3(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n351), .B(new_n404), .C1(new_n396), .C2(new_n397), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT17), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n391), .A2(new_n400), .A3(new_n405), .A4(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n346), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n277), .A2(new_n343), .ZN(new_n411));
  INV_X1    g0211(.A(G179), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n264), .A2(new_n412), .A3(new_n273), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n306), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n323), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  XOR2_X1   g0215(.A(KEYINPUT74), .B(KEYINPUT13), .Z(new_n416));
  AOI21_X1  g0216(.A(new_n270), .B1(G238), .B2(new_n272), .ZN(new_n417));
  OAI211_X1 g0217(.A(G226), .B(new_n249), .C1(new_n255), .C2(new_n256), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G97), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT72), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n254), .A2(new_n421), .A3(G232), .ZN(new_n422));
  OAI211_X1 g0222(.A(G232), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT72), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n420), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT73), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n263), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n418), .A2(new_n419), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n421), .B1(new_n254), .B2(G232), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n423), .A2(KEYINPUT72), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(KEYINPUT73), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n416), .B(new_n417), .C1(new_n427), .C2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n417), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n268), .B1(new_n431), .B2(KEYINPUT73), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n425), .A2(new_n426), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT13), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n433), .B(G179), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT76), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n417), .B1(new_n427), .B2(new_n432), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT13), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(G179), .A4(new_n433), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n433), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n435), .A2(new_n436), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n416), .B1(new_n447), .B2(new_n417), .ZN(new_n448));
  OAI21_X1  g0248(.A(G169), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT14), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT14), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n451), .B(G169), .C1(new_n446), .C2(new_n448), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n445), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  OAI22_X1  g0253(.A1(new_n359), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n284), .A2(new_n331), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n292), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT75), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n457), .A2(KEYINPUT11), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(KEYINPUT11), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT12), .B1(new_n293), .B2(G68), .ZN(new_n460));
  OR3_X1    g0260(.A1(new_n293), .A2(KEYINPUT12), .A3(G68), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n242), .B1(new_n206), .B2(G20), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n460), .A2(new_n461), .B1(new_n330), .B2(new_n462), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n458), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n453), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n416), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n441), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n248), .B1(new_n468), .B2(new_n433), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n433), .B(G190), .C1(new_n437), .C2(new_n438), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n470), .A2(new_n471), .A3(new_n464), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n415), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G116), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n206), .A2(new_n477), .A3(G13), .A4(G20), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n478), .B(KEYINPUT83), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT80), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n251), .B2(G1), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n206), .A2(KEYINPUT80), .A3(G33), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n292), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(G116), .A4(new_n293), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n291), .A2(new_n216), .B1(G20), .B2(new_n477), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  INV_X1    g0287(.A(G97), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n207), .C1(G33), .C2(new_n488), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n486), .A2(KEYINPUT20), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT20), .B1(new_n486), .B2(new_n489), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n479), .B(new_n485), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(G264), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT82), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n252), .A2(new_n253), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT82), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n495), .A2(new_n496), .A3(G264), .A4(G1698), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n257), .A2(G303), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n495), .A2(G257), .A3(new_n249), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n494), .A2(new_n497), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n263), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n206), .A2(G45), .ZN(new_n502));
  OR2_X1    g0302(.A1(KEYINPUT5), .A2(G41), .ZN(new_n503));
  NAND2_X1  g0303(.A1(KEYINPUT5), .A2(G41), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G274), .A3(new_n268), .ZN(new_n506));
  INV_X1    g0306(.A(G45), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(G1), .ZN(new_n508));
  INV_X1    g0308(.A(new_n504), .ZN(new_n509));
  NOR2_X1   g0309(.A1(KEYINPUT5), .A2(G41), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(G270), .A3(new_n268), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n501), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n492), .B1(new_n515), .B2(G200), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n278), .B2(new_n515), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n501), .A2(new_n492), .A3(G179), .A4(new_n514), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT84), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n513), .B1(new_n500), .B2(new_n263), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n521), .A2(KEYINPUT84), .A3(G179), .A4(new_n492), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n492), .A2(G169), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT85), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT21), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n524), .A2(new_n521), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n525), .B(new_n526), .C1(new_n524), .C2(new_n521), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n517), .A2(new_n523), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(G250), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n532));
  OAI211_X1 g0332(.A(G244), .B(new_n249), .C1(new_n255), .C2(new_n256), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n487), .B(new_n532), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT4), .B1(new_n260), .B2(G244), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n263), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n511), .A2(G257), .A3(new_n268), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n506), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G190), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n359), .A2(new_n331), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(G107), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n545), .A2(KEYINPUT6), .A3(G97), .ZN(new_n546));
  XNOR2_X1  g0346(.A(G97), .B(G107), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT6), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n544), .B1(new_n549), .B2(new_n207), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n545), .B1(new_n371), .B2(new_n354), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n292), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n293), .A2(G97), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n330), .A2(new_n483), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(G97), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n248), .B1(new_n537), .B2(new_n539), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n540), .A2(new_n343), .B1(new_n552), .B2(new_n555), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n537), .A2(new_n412), .A3(new_n539), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n542), .A2(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n554), .A2(G107), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n293), .A2(G107), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n563), .B(KEYINPUT25), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n207), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT22), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT22), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n495), .A2(new_n568), .A3(new_n207), .A4(G87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G116), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(G20), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT23), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n207), .B2(G107), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n545), .A2(KEYINPUT23), .A3(G20), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT24), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT24), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n570), .A2(new_n579), .A3(new_n576), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n565), .B1(new_n581), .B2(new_n292), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT86), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n254), .A2(new_n583), .A3(G257), .ZN(new_n584));
  OAI211_X1 g0384(.A(G257), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT86), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(G250), .B(new_n249), .C1(new_n255), .C2(new_n256), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G294), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n511), .A2(G264), .A3(new_n268), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n511), .A2(KEYINPUT87), .A3(G264), .A4(new_n268), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n592), .A2(new_n263), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(G200), .B1(new_n597), .B2(new_n506), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n590), .B1(new_n584), .B2(new_n586), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n599), .B(new_n506), .C1(new_n268), .C2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(G190), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n582), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n570), .A2(new_n579), .A3(new_n576), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n579), .B1(new_n570), .B2(new_n576), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n292), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n565), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n597), .A2(new_n412), .A3(new_n506), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n601), .A2(new_n343), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  OR2_X1    g0411(.A1(G238), .A2(G1698), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n339), .A2(G1698), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n612), .B(new_n613), .C1(new_n255), .C2(new_n256), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n268), .B1(new_n614), .B2(new_n571), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT81), .B1(new_n507), .B2(G1), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT81), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(new_n206), .A3(G45), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n268), .A2(new_n616), .A3(new_n618), .A4(G250), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n268), .A2(G274), .A3(new_n508), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G190), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT19), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n207), .B1(new_n419), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(G97), .A2(G107), .ZN(new_n626));
  INV_X1    g0426(.A(G87), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n207), .B(G68), .C1(new_n255), .C2(new_n256), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n624), .B1(new_n284), .B2(new_n488), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n632), .A2(new_n292), .B1(new_n294), .B2(new_n326), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n330), .A2(G87), .A3(new_n483), .ZN(new_n634));
  OAI21_X1  g0434(.A(G200), .B1(new_n615), .B2(new_n621), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n623), .A2(new_n633), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n632), .A2(new_n292), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n326), .A2(new_n294), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n330), .A2(new_n483), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n637), .B(new_n638), .C1(new_n326), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n622), .A2(new_n412), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n343), .B1(new_n615), .B2(new_n621), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n561), .A2(new_n603), .A3(new_n611), .A4(new_n645), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n476), .A2(new_n531), .A3(new_n646), .ZN(G372));
  INV_X1    g0447(.A(new_n414), .ZN(new_n648));
  INV_X1    g0448(.A(new_n323), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n391), .A2(new_n400), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n464), .A2(new_n471), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n345), .B1(new_n651), .B2(new_n470), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n453), .B2(new_n465), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n405), .A2(new_n408), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT92), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n649), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI211_X1 g0457(.A(KEYINPUT92), .B(new_n650), .C1(new_n653), .C2(new_n654), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n648), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n523), .A2(new_n529), .A3(new_n530), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT90), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n523), .A2(new_n529), .A3(KEYINPUT90), .A4(new_n530), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n660), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n643), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT89), .B1(new_n633), .B2(new_n634), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n633), .A2(KEYINPUT89), .A3(new_n634), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT88), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n635), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(KEYINPUT88), .B(G200), .C1(new_n615), .C2(new_n621), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n672), .A2(new_n623), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n666), .B1(new_n670), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n561), .A2(new_n675), .A3(new_n603), .ZN(new_n676));
  INV_X1    g0476(.A(new_n560), .ZN(new_n677));
  INV_X1    g0477(.A(new_n553), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n639), .B2(new_n488), .ZN(new_n679));
  OAI21_X1  g0479(.A(G107), .B1(new_n353), .B2(new_n355), .ZN(new_n680));
  AND2_X1   g0480(.A1(G97), .A2(G107), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n548), .B1(new_n681), .B2(new_n626), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n545), .A2(KEYINPUT6), .A3(G97), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n543), .B1(new_n684), .B2(G20), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n679), .B1(new_n686), .B2(new_n292), .ZN(new_n687));
  AOI21_X1  g0487(.A(G169), .B1(new_n537), .B2(new_n539), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n677), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n635), .A2(new_n671), .B1(new_n622), .B2(G190), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n633), .A2(KEYINPUT89), .A3(new_n634), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n691), .B(new_n673), .C1(new_n692), .C2(new_n667), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n689), .A2(new_n690), .A3(new_n693), .A4(new_n643), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n556), .B(new_n560), .C1(new_n541), .C2(G169), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT26), .B1(new_n695), .B2(new_n644), .ZN(new_n696));
  AND4_X1   g0496(.A1(KEYINPUT91), .A2(new_n694), .A3(new_n643), .A4(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n559), .A2(new_n560), .A3(new_n643), .A4(new_n636), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n666), .B1(new_n698), .B2(KEYINPUT26), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT91), .B1(new_n699), .B2(new_n694), .ZN(new_n700));
  OAI22_X1  g0500(.A1(new_n665), .A2(new_n676), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n659), .B1(new_n476), .B2(new_n702), .ZN(G369));
  NAND3_X1  g0503(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G213), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G343), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n492), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n663), .B2(new_n664), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n531), .B2(new_n710), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT93), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n608), .A2(new_n709), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n660), .B1(new_n603), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n709), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n718), .B1(new_n660), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n661), .A2(new_n719), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n724), .B1(new_n660), .B2(new_n719), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n721), .A2(new_n725), .ZN(G399));
  INV_X1    g0526(.A(new_n210), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G41), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n628), .A2(G116), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n729), .A2(G1), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(new_n214), .B2(new_n729), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT28), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT29), .B1(new_n701), .B2(new_n719), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n661), .A2(new_n660), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n676), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n695), .A2(new_n644), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n666), .B1(new_n737), .B2(new_n690), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n693), .A2(new_n643), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT26), .B1(new_n739), .B2(new_n695), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n719), .B1(new_n736), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(KEYINPUT95), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n740), .B(new_n738), .C1(new_n735), .C2(new_n676), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT95), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n744), .A2(new_n745), .A3(new_n719), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n734), .B1(new_n747), .B2(KEYINPUT29), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G330), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT31), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n540), .A2(new_n615), .A3(new_n621), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n515), .A2(new_n412), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(new_n753), .A3(new_n597), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT30), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n752), .A2(new_n753), .A3(KEYINPUT30), .A4(new_n597), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n622), .A2(G179), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n601), .A2(new_n515), .A3(new_n540), .A4(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n751), .B(new_n719), .C1(new_n758), .C2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n756), .A2(new_n757), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n760), .B(KEYINPUT94), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n709), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n646), .A2(new_n531), .A3(new_n709), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n765), .B1(new_n766), .B2(new_n751), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n750), .B1(new_n762), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n749), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n733), .B1(new_n771), .B2(G1), .ZN(G364));
  AND2_X1   g0572(.A1(new_n207), .A2(G13), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n206), .B1(new_n773), .B2(G45), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n728), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n727), .A2(new_n257), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n778), .A2(G355), .B1(new_n477), .B2(new_n727), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n727), .A2(new_n495), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(G45), .B2(new_n214), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n246), .A2(new_n507), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n216), .B1(G20), .B2(new_n343), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n777), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT96), .ZN(new_n790));
  INV_X1    g0590(.A(new_n787), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n207), .A2(new_n412), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G190), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n278), .A2(G179), .A3(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n207), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n495), .B1(new_n794), .B2(new_n331), .C1(new_n796), .C2(new_n488), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n207), .A2(G179), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(new_n278), .A3(G200), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n545), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n792), .A2(G200), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n278), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n800), .B1(G50), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n801), .A2(G190), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n803), .B1(new_n242), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n792), .A2(G190), .A3(new_n248), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT97), .Z(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n797), .B(new_n806), .C1(new_n363), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n798), .A2(new_n793), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT98), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(KEYINPUT98), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(KEYINPUT99), .B(G159), .Z(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n798), .A2(G190), .A3(G200), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n819), .A2(KEYINPUT100), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(KEYINPUT100), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n818), .A2(KEYINPUT32), .B1(G87), .B2(new_n823), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n810), .B(new_n824), .C1(KEYINPUT32), .C2(new_n818), .ZN(new_n825));
  INV_X1    g0625(.A(new_n802), .ZN(new_n826));
  INV_X1    g0626(.A(G326), .ZN(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n826), .A2(new_n827), .B1(new_n828), .B2(new_n799), .ZN(new_n829));
  OR2_X1    g0629(.A1(KEYINPUT33), .A2(G317), .ZN(new_n830));
  NAND2_X1  g0630(.A1(KEYINPUT33), .A2(G317), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n805), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n796), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n829), .B(new_n832), .C1(G294), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n823), .A2(G303), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n815), .A2(G329), .ZN(new_n836));
  INV_X1    g0636(.A(G311), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n257), .B1(new_n794), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n807), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(G322), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n825), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n786), .B(KEYINPUT101), .Z(new_n843));
  OAI221_X1 g0643(.A(new_n790), .B1(new_n791), .B2(new_n842), .C1(new_n714), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n715), .A2(new_n777), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n714), .A2(G330), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT102), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G396));
  NAND2_X1  g0649(.A1(new_n701), .A2(new_n719), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n342), .B1(new_n335), .B2(new_n719), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n345), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n345), .A2(new_n709), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n850), .B(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(new_n769), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n856), .A2(new_n769), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n776), .B(new_n857), .C1(KEYINPUT104), .C2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(KEYINPUT104), .B2(new_n858), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n787), .A2(new_n784), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n777), .B1(new_n331), .B2(new_n861), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n833), .A2(G97), .B1(new_n839), .B2(G294), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n864), .A2(KEYINPUT103), .B1(new_n823), .B2(G107), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(KEYINPUT103), .B2(new_n864), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n814), .A2(new_n837), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n257), .B1(new_n477), .B2(new_n794), .C1(new_n805), .C2(new_n828), .ZN(new_n868));
  INV_X1    g0668(.A(G303), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n826), .A2(new_n869), .B1(new_n627), .B2(new_n799), .ZN(new_n870));
  NOR4_X1   g0670(.A1(new_n866), .A2(new_n867), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n257), .B1(new_n833), .B2(new_n363), .ZN(new_n872));
  INV_X1    g0672(.A(G132), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n872), .B1(new_n242), .B2(new_n799), .C1(new_n814), .C2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n794), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n802), .A2(G137), .B1(new_n817), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(G150), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n877), .B2(new_n805), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(G143), .B2(new_n809), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n879), .A2(KEYINPUT34), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n874), .B(new_n880), .C1(G50), .C2(new_n823), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(KEYINPUT34), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n871), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n853), .B1(new_n851), .B2(new_n345), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n862), .B1(new_n883), .B2(new_n791), .C1(new_n884), .C2(new_n785), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n860), .A2(new_n885), .ZN(G384));
  OR2_X1    g0686(.A1(new_n684), .A2(KEYINPUT35), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n684), .A2(KEYINPUT35), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n887), .A2(new_n888), .A3(G116), .A4(new_n217), .ZN(new_n889));
  XNOR2_X1  g0689(.A(KEYINPUT105), .B(KEYINPUT36), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n889), .B(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n215), .A2(G77), .A3(new_n366), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n206), .B(G13), .C1(new_n892), .C2(new_n241), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n773), .A2(new_n206), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT108), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n748), .B2(new_n475), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n744), .A2(new_n745), .A3(new_n719), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n745), .B1(new_n744), .B2(new_n719), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT29), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT29), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n850), .A2(new_n901), .ZN(new_n902));
  AND4_X1   g0702(.A1(new_n896), .A2(new_n475), .A3(new_n900), .A4(new_n902), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n659), .ZN(new_n905));
  INV_X1    g0705(.A(new_n707), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n650), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n854), .B1(new_n850), .B2(new_n855), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n464), .A2(new_n719), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n466), .A2(new_n473), .A3(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n465), .B(new_n709), .C1(new_n453), .C2(new_n472), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n368), .A2(new_n365), .A3(new_n356), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n915), .A2(new_n376), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n351), .B1(new_n916), .B2(new_n397), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n906), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n409), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n398), .A2(new_n389), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n398), .A2(new_n906), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT37), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n921), .A2(new_n922), .A3(new_n923), .A4(new_n406), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n917), .A2(new_n389), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n918), .A2(new_n925), .A3(new_n406), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n924), .B1(new_n926), .B2(new_n923), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n920), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT38), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n920), .A2(new_n927), .A3(KEYINPUT38), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n907), .B1(new_n914), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT107), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n920), .A2(new_n927), .A3(KEYINPUT107), .A4(KEYINPUT38), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n380), .A2(new_n707), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n409), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n406), .B1(new_n380), .B2(new_n390), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT37), .B1(new_n941), .B2(new_n939), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n940), .A2(KEYINPUT106), .B1(new_n924), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT106), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n409), .A2(new_n944), .A3(new_n939), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n929), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT39), .B1(new_n938), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n932), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n466), .A2(new_n709), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n934), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n905), .B(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n764), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n719), .B1(new_n758), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(KEYINPUT31), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n767), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n855), .B1(new_n911), .B2(new_n912), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n936), .A2(new_n937), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT38), .B1(new_n943), .B2(new_n945), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n958), .B(new_n959), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT40), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n913), .A2(new_n884), .A3(new_n958), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT40), .B1(new_n930), .B2(new_n931), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n475), .A2(new_n958), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n969), .A2(new_n970), .A3(new_n750), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n895), .B1(new_n954), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT109), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n972), .A2(new_n973), .B1(new_n954), .B2(new_n971), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n894), .B1(new_n974), .B2(new_n975), .ZN(G367));
  AOI21_X1  g0776(.A(new_n257), .B1(new_n875), .B2(G50), .ZN(new_n977));
  INV_X1    g0777(.A(G137), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n977), .B1(new_n877), .B2(new_n807), .C1(new_n814), .C2(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n817), .A2(new_n804), .B1(new_n802), .B2(G143), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n799), .A2(new_n331), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n980), .B(new_n982), .C1(new_n242), .C2(new_n796), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n979), .B(new_n983), .C1(new_n363), .C2(new_n823), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n808), .A2(new_n869), .ZN(new_n985));
  INV_X1    g0785(.A(G317), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n814), .A2(new_n986), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n257), .B1(new_n794), .B2(new_n828), .C1(new_n796), .C2(new_n545), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT46), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n823), .A2(G116), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n990), .B1(new_n991), .B2(KEYINPUT114), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n804), .A2(G294), .ZN(new_n993));
  INV_X1    g0793(.A(new_n799), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(G97), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n993), .B(new_n995), .C1(new_n826), .C2(new_n837), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n989), .A2(new_n992), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n991), .A2(KEYINPUT114), .A3(new_n990), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n984), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(KEYINPUT115), .B(KEYINPUT47), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n787), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n668), .A2(new_n669), .A3(new_n709), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n675), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n643), .B2(new_n1003), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(new_n843), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n780), .A2(new_n230), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n788), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n326), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1008), .B1(new_n727), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n777), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1002), .A2(new_n1006), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n561), .B1(new_n687), .B2(new_n719), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT110), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n689), .A2(new_n709), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n725), .A2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT44), .Z(new_n1018));
  NAND2_X1  g0818(.A1(new_n725), .A2(new_n1016), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT45), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT113), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n721), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n716), .A2(KEYINPUT113), .A3(new_n720), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1022), .B(new_n721), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n720), .B(new_n722), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n715), .B(new_n1028), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(new_n770), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n771), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n728), .B(KEYINPUT41), .Z(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n775), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n724), .A2(new_n1016), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1037), .A2(KEYINPUT42), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT111), .Z(new_n1039));
  OAI21_X1  g0839(.A(new_n695), .B1(new_n1014), .B2(new_n611), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1037), .A2(KEYINPUT42), .B1(new_n719), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(KEYINPUT112), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT112), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1042), .A2(new_n1047), .A3(new_n1043), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1046), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1016), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1049), .A2(new_n1050), .B1(new_n721), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1046), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n721), .A2(new_n1051), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1052), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1012), .B1(new_n1036), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT116), .ZN(G387));
  NAND2_X1  g0861(.A1(new_n1029), .A2(new_n770), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1030), .A2(new_n728), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n730), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n778), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(G107), .B2(new_n210), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n780), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n324), .A2(new_n202), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT50), .Z(new_n1069));
  AOI211_X1 g0869(.A(G45), .B(new_n1064), .C1(G68), .C2(G77), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n236), .A2(G45), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1066), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n776), .B1(new_n1073), .B2(new_n1008), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n796), .A2(new_n326), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1076), .B(new_n995), .C1(new_n360), .C2(new_n826), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G77), .B2(new_n823), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n347), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n804), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n815), .A2(G150), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n495), .B1(new_n807), .B2(new_n202), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G68), .B2(new_n875), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n495), .B1(new_n994), .B2(G116), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n805), .A2(new_n837), .B1(new_n794), .B2(new_n869), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G322), .B2(new_n802), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n986), .B2(new_n808), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT48), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n823), .A2(G294), .B1(G283), .B2(new_n833), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT49), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1085), .B1(new_n827), .B2(new_n814), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1084), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT118), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n791), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1074), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n720), .B2(new_n843), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1063), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1029), .A2(new_n774), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT117), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(G393));
  NAND3_X1  g0906(.A1(new_n1025), .A2(new_n1030), .A3(new_n1026), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1032), .A2(new_n728), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1051), .A2(new_n786), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n788), .B1(new_n488), .B2(new_n210), .C1(new_n1067), .C2(new_n240), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n776), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G150), .A2(new_n802), .B1(new_n839), .B2(G159), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT51), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n823), .A2(G68), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n815), .A2(G143), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n799), .A2(new_n627), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n257), .B(new_n1116), .C1(new_n324), .C2(new_n875), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G77), .A2(new_n833), .B1(new_n804), .B2(G50), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n823), .A2(G283), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n815), .A2(G322), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n495), .B(new_n800), .C1(G294), .C2(new_n875), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G116), .A2(new_n833), .B1(new_n804), .B2(G303), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G317), .A2(new_n802), .B1(new_n839), .B2(G311), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT52), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1113), .A2(new_n1119), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1111), .B1(new_n1127), .B2(new_n787), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1027), .A2(new_n775), .B1(new_n1109), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1108), .A2(new_n1129), .ZN(G390));
  INV_X1    g0930(.A(new_n952), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n914), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n948), .B2(new_n950), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n959), .A2(new_n768), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n952), .B1(new_n938), .B2(new_n947), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n743), .A2(new_n746), .A3(new_n854), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1136), .A2(new_n913), .A3(new_n852), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT119), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n945), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n942), .A2(new_n924), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n944), .B1(new_n409), .B2(new_n939), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n936), .B(new_n937), .C1(new_n1142), .C2(KEYINPUT38), .ZN(new_n1143));
  AND4_X1   g0943(.A1(KEYINPUT119), .A2(new_n1143), .A3(new_n1137), .A4(new_n1131), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1133), .B(new_n1134), .C1(new_n1138), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT119), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1143), .A2(new_n1131), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1137), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1135), .A2(KEYINPUT119), .A3(new_n1137), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1143), .A2(new_n949), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n950), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1149), .A2(new_n1150), .B1(new_n1153), .B2(new_n1132), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n913), .A2(G330), .A3(new_n884), .A4(new_n958), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1145), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1153), .A2(new_n784), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n861), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n776), .B1(new_n1079), .B2(new_n1159), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n805), .A2(new_n545), .B1(new_n826), .B2(new_n828), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n796), .A2(new_n331), .B1(new_n799), .B2(new_n242), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n823), .A2(G87), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n815), .A2(G294), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n257), .B1(new_n807), .B2(new_n477), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G97), .B2(new_n875), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(G128), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n805), .A2(new_n978), .B1(new_n826), .B2(new_n1169), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n796), .A2(new_n360), .B1(new_n799), .B2(new_n202), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(KEYINPUT53), .B1(new_n822), .B2(new_n877), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n815), .A2(G125), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n495), .B1(new_n807), .B2(new_n873), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT54), .B(G143), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1175), .B1(new_n875), .B2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1178), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n822), .A2(KEYINPUT53), .A3(new_n877), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1168), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1160), .B1(new_n1181), .B2(new_n787), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1157), .A2(new_n775), .B1(new_n1158), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n475), .A2(G330), .A3(new_n958), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n659), .B(new_n1184), .C1(new_n897), .C2(new_n903), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n531), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n561), .A2(new_n603), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n660), .A2(new_n644), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .A4(new_n719), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n956), .B1(KEYINPUT31), .B2(new_n1189), .ZN(new_n1190));
  OAI211_X1 g0990(.A(G330), .B(new_n884), .C1(new_n1190), .C2(new_n761), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1155), .B1(new_n1192), .B2(new_n913), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n959), .A2(new_n768), .B1(new_n1136), .B2(new_n852), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n913), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n958), .A2(G330), .A3(new_n884), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1193), .A2(new_n908), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1185), .A2(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1199), .B(new_n1145), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT120), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1200), .A2(new_n1201), .A3(new_n728), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1199), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1156), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1201), .B1(new_n1200), .B2(new_n728), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1183), .B1(new_n1205), .B2(new_n1206), .ZN(G378));
  INV_X1    g1007(.A(new_n1185), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1200), .A2(new_n1208), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n907), .B1(new_n933), .B2(new_n914), .C1(new_n1153), .C2(new_n1131), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n306), .B(new_n906), .C1(new_n649), .C2(new_n648), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n306), .A2(new_n906), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n323), .A2(new_n414), .A3(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1211), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1214), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n967), .B2(G330), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n962), .A2(KEYINPUT40), .B1(new_n964), .B2(new_n965), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1220), .A2(new_n750), .A3(new_n1217), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1210), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n967), .A2(new_n1218), .A3(G330), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1217), .B1(new_n1220), .B2(new_n750), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(new_n1224), .A3(new_n953), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1209), .A2(new_n1226), .A3(KEYINPUT57), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT57), .B1(new_n1209), .B2(new_n1226), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT123), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n728), .B(new_n1227), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1230));
  AOI211_X1 g1030(.A(KEYINPUT123), .B(KEYINPUT57), .C1(new_n1209), .C2(new_n1226), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G150), .A2(new_n833), .B1(new_n802), .B2(G125), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT122), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n839), .A2(G128), .B1(new_n875), .B2(G137), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1235), .B1(new_n873), .B2(new_n805), .C1(new_n822), .C2(new_n1176), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n815), .A2(G124), .ZN(new_n1240));
  AOI211_X1 g1040(.A(G33), .B(G41), .C1(new_n817), .C2(new_n994), .ZN(new_n1241));
  AND4_X1   g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n495), .A2(G41), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1243), .B1(new_n326), .B2(new_n794), .C1(new_n545), .C2(new_n807), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n815), .B2(G283), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n823), .A2(G77), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G68), .A2(new_n833), .B1(new_n804), .B2(G97), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n802), .A2(G116), .B1(new_n994), .B2(new_n363), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  XOR2_X1   g1049(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n1250));
  OR2_X1    g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1251), .B(new_n1252), .C1(new_n1243), .C2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n787), .B1(new_n1242), .B2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1255), .B(new_n776), .C1(G50), .C2(new_n1159), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1217), .B2(new_n784), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1226), .B2(new_n775), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1232), .A2(new_n1258), .ZN(G375));
  NAND2_X1  g1059(.A1(new_n1185), .A2(new_n1198), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1203), .A2(new_n1035), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1195), .A2(new_n784), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT124), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n804), .A2(G116), .B1(new_n802), .B2(G294), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1264), .A2(new_n982), .A3(new_n1076), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n257), .B1(new_n794), .B2(new_n545), .C1(new_n828), .C2(new_n807), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n815), .B2(G303), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1265), .B(new_n1267), .C1(new_n488), .C2(new_n822), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1268), .A2(KEYINPUT125), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(KEYINPUT125), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n363), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n495), .B1(new_n794), .B2(new_n877), .C1(new_n1271), .C2(new_n799), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n815), .B2(G128), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n978), .B2(new_n808), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(G132), .A2(new_n802), .B1(new_n804), .B2(new_n1177), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1275), .B1(new_n202), .B2(new_n796), .C1(new_n360), .C2(new_n822), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1269), .B(new_n1270), .C1(new_n1274), .C2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n787), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n777), .B1(new_n242), .B2(new_n861), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1263), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n774), .B2(new_n1198), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1261), .A2(new_n1282), .ZN(G381));
  NAND3_X1  g1083(.A1(new_n1103), .A2(new_n848), .A3(new_n1105), .ZN(new_n1284));
  OR4_X1    g1084(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1284), .ZN(new_n1285));
  OR4_X1    g1085(.A1(G387), .A2(G378), .A3(G375), .A4(new_n1285), .ZN(G407));
  INV_X1    g1086(.A(G378), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n708), .A2(G213), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1232), .A2(new_n1287), .A3(new_n1258), .A4(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(G407), .A2(G213), .A3(new_n1290), .ZN(G409));
  INV_X1    g1091(.A(KEYINPUT61), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G378), .B(new_n1258), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1209), .A2(new_n1035), .A3(new_n1226), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1258), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1287), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1289), .B1(new_n1293), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1289), .A2(G2897), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT60), .B1(new_n1185), .B2(new_n1198), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n729), .B1(new_n1300), .B2(new_n1260), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1185), .A2(KEYINPUT60), .A3(new_n1198), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1301), .A2(KEYINPUT126), .A3(new_n1302), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1281), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1307), .A2(G384), .ZN(new_n1308));
  INV_X1    g1108(.A(G384), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n1281), .B(new_n1309), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1299), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1306), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT126), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1282), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1309), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1307), .A2(G384), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1315), .A2(new_n1316), .A3(new_n1298), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1311), .A2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1292), .B1(new_n1297), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1288), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1321), .B1(new_n1323), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1060), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(G393), .A2(G396), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1284), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G390), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT116), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1331), .B1(new_n1328), .B2(new_n1284), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1330), .B1(G390), .B2(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1327), .A2(new_n1333), .ZN(new_n1334));
  OR2_X1    g1134(.A1(new_n1332), .A2(G390), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1060), .B1(new_n1335), .B2(new_n1330), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1334), .A2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1297), .A2(KEYINPUT63), .A3(new_n1324), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1320), .A2(new_n1326), .A3(new_n1337), .A4(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT62), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1297), .A2(new_n1340), .A3(new_n1324), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1340), .B1(new_n1297), .B2(new_n1324), .ZN(new_n1342));
  NOR3_X1   g1142(.A1(new_n1341), .A2(new_n1319), .A3(new_n1342), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1339), .B1(new_n1343), .B2(new_n1337), .ZN(G405));
  NAND2_X1  g1144(.A1(new_n1327), .A2(new_n1333), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1335), .A2(new_n1060), .A3(new_n1330), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT127), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(G378), .B1(new_n1232), .B2(new_n1258), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1293), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1324), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(G375), .A2(new_n1287), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1353), .A2(new_n1325), .A3(new_n1293), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1345), .A2(new_n1346), .A3(KEYINPUT127), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1349), .A2(new_n1352), .A3(new_n1354), .A4(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1325), .B1(new_n1353), .B2(new_n1293), .ZN(new_n1357));
  NOR3_X1   g1157(.A1(new_n1350), .A2(new_n1324), .A3(new_n1351), .ZN(new_n1358));
  OAI211_X1 g1158(.A(new_n1348), .B(new_n1347), .C1(new_n1357), .C2(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1356), .A2(new_n1359), .ZN(G402));
endmodule


