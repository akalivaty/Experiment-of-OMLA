//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1322, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n210), .B(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT66), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n212), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n205), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n208), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n230));
  AND3_X1   g0030(.A1(new_n219), .A2(new_n229), .A3(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT67), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G45), .ZN(new_n250));
  AOI21_X1  g0050(.A(G1), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G1), .A3(G13), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(new_n253), .A3(G274), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT69), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n256), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n253), .A2(new_n256), .A3(new_n258), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n255), .B1(new_n262), .B2(G226), .ZN(new_n263));
  OR2_X1    g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1698), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G222), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n265), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G223), .A3(G1698), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n267), .B(new_n269), .C1(new_n205), .C2(new_n268), .ZN(new_n270));
  INV_X1    g0070(.A(new_n253), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n263), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G169), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT8), .B(G58), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT71), .ZN(new_n277));
  INV_X1    g0077(.A(G58), .ZN(new_n278));
  OR3_X1    g0078(.A1(new_n278), .A2(KEYINPUT71), .A3(KEYINPUT8), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G20), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n277), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G150), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n282), .B(new_n284), .C1(new_n204), .C2(new_n214), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n286), .A2(KEYINPUT70), .A3(new_n213), .ZN(new_n287));
  AOI21_X1  g0087(.A(KEYINPUT70), .B1(new_n286), .B2(new_n213), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n286), .A2(new_n213), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT70), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n286), .A2(KEYINPUT70), .A3(new_n213), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n257), .A2(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G50), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n297), .A2(new_n300), .B1(new_n202), .B2(new_n292), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n290), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n263), .A2(new_n272), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n275), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n290), .A2(KEYINPUT9), .A3(new_n301), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT75), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n263), .B2(new_n272), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT76), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n263), .A2(new_n272), .A3(G190), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n310), .A2(new_n313), .A3(new_n314), .A4(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT10), .B1(new_n308), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT75), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n307), .B(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT10), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n315), .A2(new_n314), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT9), .B1(new_n290), .B2(new_n301), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n321), .A2(new_n322), .A3(new_n312), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n319), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n306), .B1(new_n317), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(G232), .A2(G1698), .ZN(new_n326));
  INV_X1    g0126(.A(G238), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(G1698), .ZN(new_n328));
  AND2_X1   g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  NOR2_X1   g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n271), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n268), .A2(G107), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n254), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n221), .B1(new_n260), .B2(new_n261), .ZN(new_n335));
  OAI21_X1  g0135(.A(G200), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n205), .B1(new_n257), .B2(G20), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n297), .A2(new_n337), .B1(new_n205), .B2(new_n292), .ZN(new_n338));
  XOR2_X1   g0138(.A(KEYINPUT8), .B(G58), .Z(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(new_n283), .B1(G20), .B2(G77), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT15), .B(G87), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT72), .A3(new_n281), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT72), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n214), .A2(G33), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n340), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n347), .A2(KEYINPUT73), .A3(new_n289), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT73), .B1(new_n347), .B2(new_n289), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n336), .B(new_n338), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT74), .ZN(new_n351));
  INV_X1    g0151(.A(G190), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n334), .A2(new_n335), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n350), .A2(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n338), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n347), .A2(new_n289), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT73), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n347), .A2(KEYINPUT73), .A3(new_n289), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n355), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT74), .B1(new_n360), .B2(new_n336), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  NOR3_X1   g0162(.A1(new_n334), .A2(new_n335), .A3(G179), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(new_n274), .B2(new_n353), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n338), .B1(new_n348), .B2(new_n349), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n283), .A2(G50), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n369), .B1(new_n214), .B2(G68), .C1(new_n205), .C2(new_n345), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n370), .A2(new_n289), .ZN(new_n371));
  INV_X1    g0171(.A(G68), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n292), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT12), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n373), .A2(KEYINPUT12), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n371), .A2(KEYINPUT11), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(KEYINPUT11), .B2(new_n371), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n297), .A2(G68), .A3(new_n298), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT77), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT14), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G97), .ZN(new_n383));
  INV_X1    g0183(.A(G232), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G1698), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(G226), .B2(G1698), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n383), .B1(new_n386), .B2(new_n331), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n271), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n254), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n327), .B1(new_n260), .B2(new_n261), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT13), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT13), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n255), .B1(new_n387), .B2(new_n271), .ZN(new_n393));
  INV_X1    g0193(.A(new_n261), .ZN(new_n394));
  OAI21_X1  g0194(.A(G238), .B1(new_n394), .B2(new_n259), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n392), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n382), .B(G169), .C1(new_n391), .C2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT13), .B1(new_n389), .B2(new_n390), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(new_n395), .A3(new_n392), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(G179), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n398), .A2(new_n399), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n382), .B1(new_n402), .B2(G169), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n381), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(G200), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n380), .B(new_n405), .C1(new_n352), .C2(new_n402), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n297), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n277), .A2(new_n279), .A3(new_n298), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n277), .A2(new_n279), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n409), .A2(new_n410), .B1(new_n411), .B2(new_n291), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n295), .A2(new_n296), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT7), .B1(new_n331), .B2(new_n214), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT7), .ZN(new_n415));
  NOR4_X1   g0215(.A1(new_n329), .A2(new_n330), .A3(new_n415), .A4(G20), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n278), .A2(new_n372), .ZN(new_n418));
  OAI21_X1  g0218(.A(G20), .B1(new_n418), .B2(new_n201), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n283), .A2(G159), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT16), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n413), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n422), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n412), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OR2_X1    g0227(.A1(G223), .A2(G1698), .ZN(new_n428));
  INV_X1    g0228(.A(G226), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G1698), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n428), .B(new_n430), .C1(new_n329), .C2(new_n330), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G87), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n253), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n253), .A2(G232), .A3(new_n258), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n254), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT78), .B1(new_n436), .B2(new_n303), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT78), .ZN(new_n438));
  NOR4_X1   g0238(.A1(new_n433), .A2(new_n435), .A3(new_n438), .A4(G179), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n437), .A2(new_n439), .B1(G169), .B2(new_n436), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT18), .B1(new_n427), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n415), .B1(new_n268), .B2(G20), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n331), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n372), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n424), .B1(new_n444), .B2(new_n421), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n445), .A2(new_n289), .A3(new_n426), .ZN(new_n446));
  INV_X1    g0246(.A(new_n412), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n436), .A2(G169), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n431), .A2(new_n432), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n271), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(new_n303), .A3(new_n254), .A4(new_n434), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n438), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n436), .A2(KEYINPUT78), .A3(new_n303), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n449), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT18), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n448), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n436), .A2(new_n352), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n311), .B1(new_n433), .B2(new_n435), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n446), .A2(new_n447), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT17), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n446), .A2(KEYINPUT17), .A3(new_n447), .A4(new_n460), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n441), .A2(new_n457), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AND4_X1   g0266(.A1(new_n325), .A2(new_n368), .A3(new_n408), .A4(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT81), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n222), .B1(new_n442), .B2(new_n443), .ZN(new_n470));
  INV_X1    g0270(.A(G97), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(new_n222), .A3(KEYINPUT6), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT6), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G97), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n222), .A2(KEYINPUT79), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT79), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G107), .ZN(new_n477));
  AND4_X1   g0277(.A1(new_n472), .A2(new_n474), .A3(new_n475), .A4(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n472), .A2(new_n474), .B1(new_n475), .B2(new_n477), .ZN(new_n479));
  OAI21_X1  g0279(.A(G20), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n283), .A2(G77), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n470), .B1(new_n482), .B2(KEYINPUT80), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT80), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n484), .A3(new_n481), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n413), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n291), .A2(G97), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n257), .A2(G33), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n291), .B(new_n489), .C1(new_n287), .C2(new_n288), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n488), .B1(new_n490), .B2(new_n471), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n469), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n473), .A2(G97), .A3(G107), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n471), .A2(KEYINPUT6), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n476), .A2(G107), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n222), .A2(KEYINPUT79), .ZN(new_n496));
  OAI22_X1  g0296(.A1(new_n493), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n472), .A2(new_n474), .A3(new_n475), .A4(new_n477), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n214), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n481), .ZN(new_n500));
  OAI21_X1  g0300(.A(KEYINPUT80), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n470), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n485), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n491), .B1(new_n503), .B2(new_n289), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT81), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n257), .B(G45), .C1(new_n249), .C2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT82), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(G41), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n249), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n507), .A2(new_n512), .A3(G274), .A4(new_n253), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n250), .A2(G1), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n509), .A2(G41), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(G257), .A3(new_n253), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT4), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(new_n221), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n266), .A2(new_n521), .B1(G33), .B2(G283), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n520), .B1(new_n331), .B2(new_n221), .ZN(new_n523));
  INV_X1    g0323(.A(G1698), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n520), .B1(new_n268), .B2(G250), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n522), .B(new_n523), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n519), .B1(new_n526), .B2(new_n271), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n352), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(G200), .B2(new_n527), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n492), .A2(new_n505), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n521), .B(new_n524), .C1(new_n330), .C2(new_n329), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n523), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(G250), .B1(new_n329), .B2(new_n330), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n524), .B1(new_n534), .B2(KEYINPUT4), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n271), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT83), .ZN(new_n537));
  INV_X1    g0337(.A(new_n519), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n303), .A4(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n527), .B2(G169), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n537), .B1(new_n527), .B2(new_n303), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n504), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n530), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(G264), .B(G1698), .C1(new_n329), .C2(new_n330), .ZN(new_n546));
  OAI211_X1 g0346(.A(G257), .B(new_n524), .C1(new_n329), .C2(new_n330), .ZN(new_n547));
  INV_X1    g0347(.A(G303), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n546), .B(new_n547), .C1(new_n548), .C2(new_n268), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n271), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n509), .A2(G41), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n253), .B1(new_n506), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G270), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n550), .A2(new_n554), .A3(new_n513), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G200), .ZN(new_n556));
  INV_X1    g0356(.A(G116), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n257), .A2(new_n557), .A3(G13), .A4(G20), .ZN(new_n558));
  OR2_X1    g0358(.A1(new_n558), .A2(KEYINPUT87), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(KEYINPUT87), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n286), .A2(new_n213), .B1(G20), .B2(new_n557), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n531), .B(new_n214), .C1(G33), .C2(new_n471), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n562), .A2(KEYINPUT20), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT20), .B1(new_n562), .B2(new_n563), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT86), .B1(new_n490), .B2(new_n557), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT86), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n297), .A2(new_n568), .A3(G116), .A4(new_n489), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n566), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n549), .A2(new_n271), .B1(new_n553), .B2(G270), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(G190), .A3(new_n513), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n556), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT88), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(G179), .A3(new_n513), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n555), .A2(G169), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT21), .B1(new_n578), .B2(new_n570), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n274), .B1(new_n571), .B2(new_n513), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT21), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n567), .A2(new_n569), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n580), .B(new_n581), .C1(new_n582), .C2(new_n566), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n577), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n575), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n253), .B1(G250), .B2(new_n514), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n250), .A2(G1), .A3(G274), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(G238), .B(new_n524), .C1(new_n329), .C2(new_n330), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G33), .A2(G116), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(G244), .B(G1698), .C1(new_n329), .C2(new_n330), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT84), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n268), .A2(KEYINPUT84), .A3(G244), .A4(G1698), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n589), .B1(new_n597), .B2(new_n253), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n274), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n303), .B(new_n589), .C1(new_n597), .C2(new_n253), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT19), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n214), .B1(new_n383), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(G87), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(new_n471), .A3(new_n222), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n214), .B(G68), .C1(new_n329), .C2(new_n330), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n601), .B1(new_n345), .B2(new_n471), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n608), .A2(new_n289), .B1(new_n292), .B2(new_n341), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n297), .A2(new_n342), .A3(new_n489), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n599), .A2(new_n600), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n413), .A2(G87), .A3(new_n291), .A4(new_n489), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n608), .A2(new_n289), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n341), .A2(new_n292), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n595), .A2(new_n596), .ZN(new_n619));
  INV_X1    g0419(.A(new_n592), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n588), .B1(new_n621), .B2(new_n271), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n618), .B1(new_n622), .B2(new_n311), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT85), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n623), .A2(new_n624), .B1(G190), .B2(new_n622), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n617), .B1(new_n598), .B2(G200), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT85), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n613), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n292), .A2(new_n222), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(KEYINPUT25), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n490), .A2(new_n222), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n214), .B(G87), .C1(new_n329), .C2(new_n330), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT22), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT22), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n268), .A2(new_n635), .A3(new_n214), .A4(G87), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n222), .A2(G20), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT90), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n639), .A3(KEYINPUT23), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n638), .A2(KEYINPUT23), .B1(G20), .B2(new_n591), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n639), .B1(new_n638), .B2(KEYINPUT23), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g0445(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n637), .A2(new_n644), .A3(new_n646), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT91), .B1(new_n650), .B2(new_n289), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n637), .A2(new_n644), .A3(new_n646), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n646), .B1(new_n637), .B2(new_n644), .ZN(new_n653));
  OAI211_X1 g0453(.A(KEYINPUT91), .B(new_n289), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n632), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT92), .B1(new_n552), .B2(new_n223), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT92), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n517), .A2(new_n658), .A3(G264), .A4(new_n253), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(G257), .B(G1698), .C1(new_n329), .C2(new_n330), .ZN(new_n661));
  OAI211_X1 g0461(.A(G250), .B(new_n524), .C1(new_n329), .C2(new_n330), .ZN(new_n662));
  INV_X1    g0462(.A(G294), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n661), .B(new_n662), .C1(new_n280), .C2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n271), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n660), .A2(G179), .A3(new_n513), .A4(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(KEYINPUT93), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT93), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n660), .A2(new_n513), .A3(new_n665), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G169), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n667), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n656), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n632), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n289), .B1(new_n652), .B2(new_n653), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT91), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n674), .B1(new_n677), .B2(new_n654), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n670), .A2(new_n311), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(G190), .B2(new_n670), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n628), .A2(new_n673), .A3(new_n681), .ZN(new_n682));
  NOR4_X1   g0482(.A1(new_n468), .A2(new_n545), .A3(new_n585), .A4(new_n682), .ZN(G372));
  AND2_X1   g0483(.A1(new_n441), .A2(new_n457), .ZN(new_n684));
  INV_X1    g0484(.A(new_n404), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n367), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n406), .A2(new_n463), .A3(new_n464), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n317), .A2(new_n324), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n306), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n667), .ZN(new_n691));
  INV_X1    g0491(.A(new_n671), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(new_n668), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n584), .B1(new_n678), .B2(new_n693), .ZN(new_n694));
  OAI211_X1 g0494(.A(G190), .B(new_n589), .C1(new_n597), .C2(new_n253), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n618), .B(new_n695), .C1(new_n622), .C2(new_n311), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n612), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n678), .B2(new_n680), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n694), .A2(new_n698), .A3(new_n544), .A4(new_n530), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n612), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n598), .A2(new_n274), .B1(new_n610), .B2(new_n609), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n600), .A2(new_n701), .B1(new_n626), .B2(new_n695), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n504), .A2(KEYINPUT81), .ZN(new_n703));
  AOI211_X1 g0503(.A(new_n469), .B(new_n491), .C1(new_n503), .C2(new_n289), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n702), .B(new_n542), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT26), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(KEYINPUT94), .A3(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n540), .A2(new_n504), .A3(new_n541), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n628), .A2(KEYINPUT26), .A3(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n705), .A2(new_n706), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT94), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n700), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n690), .B1(new_n468), .B2(new_n714), .ZN(G369));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  INV_X1    g0516(.A(new_n585), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n257), .A2(new_n214), .A3(G13), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n718), .A2(KEYINPUT27), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(KEYINPUT27), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G213), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G343), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n570), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n717), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n584), .A2(new_n726), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n716), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n673), .A2(new_n681), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n678), .A2(new_n724), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n731), .A2(new_n732), .B1(new_n673), .B2(new_n724), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n673), .A2(new_n681), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n584), .A2(new_n723), .ZN(new_n736));
  INV_X1    g0536(.A(new_n673), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n735), .A2(new_n736), .B1(new_n737), .B2(new_n724), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n734), .A2(new_n738), .ZN(G399));
  INV_X1    g0539(.A(new_n209), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G41), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n604), .A2(G116), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n742), .A2(G1), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(new_n217), .B2(new_n742), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT28), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT26), .B1(new_n628), .B2(new_n708), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n705), .A2(new_n706), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n699), .B(new_n612), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(KEYINPUT29), .A3(new_n724), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n713), .A2(new_n709), .A3(new_n707), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n699), .A2(new_n612), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n723), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n750), .B1(new_n753), .B2(KEYINPUT29), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n628), .A2(new_n673), .A3(new_n681), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n530), .A2(new_n544), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n755), .A2(new_n756), .A3(new_n717), .A4(new_n724), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n536), .A2(new_n571), .A3(new_n538), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n758), .A2(new_n666), .A3(new_n598), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT96), .ZN(new_n760));
  OAI21_X1  g0560(.A(KEYINPUT30), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT30), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n527), .A2(new_n622), .A3(new_n571), .ZN(new_n763));
  OAI211_X1 g0563(.A(KEYINPUT96), .B(new_n762), .C1(new_n763), .C2(new_n666), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n527), .A2(new_n622), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n765), .A2(new_n303), .A3(new_n555), .A4(new_n670), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n761), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n767), .A2(new_n723), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(KEYINPUT31), .B1(new_n767), .B2(new_n723), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n716), .B1(new_n757), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n754), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n746), .B1(new_n774), .B2(G1), .ZN(G364));
  NAND3_X1  g0575(.A1(new_n727), .A2(new_n716), .A3(new_n729), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n585), .A2(new_n725), .ZN(new_n777));
  OAI21_X1  g0577(.A(G330), .B1(new_n777), .B2(new_n728), .ZN(new_n778));
  INV_X1    g0578(.A(G13), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n257), .B1(new_n780), .B2(G45), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n741), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n776), .A2(new_n778), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G13), .A2(G33), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G20), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n727), .A2(new_n729), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n268), .A2(G355), .A3(new_n209), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(G116), .B2(new_n209), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n247), .A2(G45), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n740), .A2(new_n268), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(new_n250), .B2(new_n218), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n791), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n213), .B1(G20), .B2(new_n274), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n788), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n783), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(G20), .A2(G179), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT97), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n802), .A2(G190), .A3(new_n311), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n311), .A2(G190), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(KEYINPUT33), .B(G317), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n804), .A2(G322), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT101), .Z(new_n810));
  NOR2_X1   g0610(.A1(new_n214), .A2(G190), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n811), .A2(new_n303), .A3(G200), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT100), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G283), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR4_X1   g0618(.A1(new_n214), .A2(new_n352), .A3(new_n311), .A4(G179), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  NOR2_X1   g0621(.A1(G190), .A2(G200), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n802), .A2(new_n822), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n331), .B1(new_n820), .B2(new_n548), .C1(new_n821), .C2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(G179), .A2(G200), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT99), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n811), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n818), .B(new_n824), .C1(G329), .C2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n214), .B1(new_n827), .B2(G190), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n802), .A2(G190), .A3(G200), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n832), .A2(G294), .B1(G326), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n810), .A2(new_n830), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n831), .A2(new_n471), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(G50), .B2(new_n834), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n278), .B2(new_n803), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n816), .A2(new_n222), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n806), .A2(new_n372), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n820), .A2(new_n603), .ZN(new_n842));
  NOR4_X1   g0642(.A1(new_n840), .A2(new_n331), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(G159), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n828), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT32), .ZN(new_n846));
  INV_X1    g0646(.A(new_n823), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n847), .A2(KEYINPUT98), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(KEYINPUT98), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n843), .B(new_n846), .C1(new_n205), .C2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n836), .B1(new_n839), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n800), .B1(new_n852), .B2(new_n797), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n789), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n785), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G396));
  NAND2_X1  g0656(.A1(new_n365), .A2(new_n723), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n366), .B(new_n857), .C1(new_n354), .C2(new_n361), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n364), .A2(new_n365), .A3(new_n723), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT102), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n859), .A2(KEYINPUT102), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n724), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n753), .A2(new_n862), .B1(new_n714), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n864), .A2(new_n773), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n783), .B1(new_n864), .B2(new_n773), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n797), .A2(new_n786), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n783), .B1(G77), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n804), .A2(G143), .ZN(new_n870));
  INV_X1    g0670(.A(G137), .ZN(new_n871));
  INV_X1    g0671(.A(G150), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n870), .B1(new_n871), .B2(new_n833), .C1(new_n872), .C2(new_n806), .ZN(new_n873));
  INV_X1    g0673(.A(new_n850), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n873), .B1(G159), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT34), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n268), .B1(new_n820), .B2(new_n202), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n816), .A2(new_n372), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n877), .B(new_n878), .C1(G132), .C2(new_n829), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n278), .B2(new_n831), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n837), .B1(G303), .B2(new_n834), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n663), .B2(new_n803), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n816), .A2(new_n603), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n331), .B1(new_n820), .B2(new_n222), .C1(new_n817), .C2(new_n806), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n883), .B(new_n884), .C1(G311), .C2(new_n829), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n557), .B2(new_n850), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n876), .A2(new_n880), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n869), .B1(new_n887), .B2(new_n797), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n787), .B2(new_n862), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT103), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n867), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(G384));
  NOR2_X1   g0692(.A1(new_n478), .A2(new_n479), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n894), .A2(KEYINPUT35), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(KEYINPUT35), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n895), .A2(G116), .A3(new_n216), .A4(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT36), .ZN(new_n898));
  OAI21_X1  g0698(.A(G77), .B1(new_n278), .B2(new_n372), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n899), .A2(new_n217), .B1(G50), .B2(new_n372), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(G1), .A3(new_n779), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT104), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n467), .B(new_n750), .C1(new_n753), .C2(KEYINPUT29), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n690), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT108), .Z(new_n906));
  NOR2_X1   g0706(.A1(new_n366), .A2(new_n723), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n714), .B2(new_n863), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n427), .A2(new_n721), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n465), .A2(new_n910), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n440), .A2(new_n721), .B1(new_n446), .B2(new_n447), .ZN(new_n912));
  INV_X1    g0712(.A(new_n461), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT37), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n721), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n448), .B1(new_n455), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT37), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n917), .A3(new_n461), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n911), .A2(KEYINPUT38), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT38), .B1(new_n911), .B2(new_n919), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n381), .A2(new_n723), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n404), .A2(new_n406), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n925), .B1(new_n404), .B2(new_n406), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n909), .A2(new_n924), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT39), .B1(new_n920), .B2(new_n922), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT105), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT105), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n933), .B(KEYINPUT39), .C1(new_n920), .C2(new_n922), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n913), .A2(KEYINPUT106), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT106), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n461), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n936), .A2(new_n916), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT107), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT37), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n461), .A2(new_n937), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(new_n912), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n917), .B1(new_n943), .B2(new_n938), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n918), .A2(KEYINPUT107), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n941), .B(new_n911), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT38), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n920), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n932), .A2(new_n934), .B1(new_n935), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n685), .A2(new_n724), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n930), .B1(new_n684), .B2(new_n915), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n906), .B(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n927), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n404), .A2(new_n406), .A3(new_n925), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n859), .B(KEYINPUT102), .Z(new_n955));
  AOI22_X1  g0755(.A1(new_n953), .A2(new_n954), .B1(new_n955), .B2(new_n858), .ZN(new_n956));
  NOR4_X1   g0756(.A1(new_n682), .A2(new_n545), .A3(new_n585), .A4(new_n723), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n767), .A2(KEYINPUT31), .A3(new_n723), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n767), .A2(new_n723), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n958), .B1(new_n959), .B2(new_n768), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n956), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT40), .B1(new_n961), .B2(new_n948), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT40), .B1(new_n921), .B2(new_n923), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n862), .B1(new_n926), .B2(new_n927), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n768), .B1(new_n767), .B2(new_n723), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(KEYINPUT31), .B2(new_n959), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n966), .B2(new_n757), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n962), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n757), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n970), .A2(new_n467), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n716), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n971), .B2(new_n969), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n952), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n257), .B2(new_n780), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n952), .A2(new_n973), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n903), .B1(new_n975), .B2(new_n976), .ZN(G367));
  INV_X1    g0777(.A(KEYINPUT109), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n492), .A2(new_n505), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n979), .A2(new_n542), .A3(new_n723), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n723), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n981), .B1(new_n756), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n736), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n731), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n978), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n756), .A2(new_n982), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n980), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n989), .A2(KEYINPUT109), .A3(new_n985), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(KEYINPUT42), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT42), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n987), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n544), .B1(new_n983), .B2(new_n673), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n724), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n992), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n702), .B1(new_n618), .B2(new_n724), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n613), .A2(new_n617), .A3(new_n723), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT43), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(KEYINPUT43), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n997), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n734), .A2(new_n983), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n991), .A2(KEYINPUT42), .B1(new_n995), .B2(new_n724), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1007), .A2(new_n1002), .A3(new_n1001), .A4(new_n994), .ZN(new_n1008));
  AND3_X1   g0808(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1006), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n741), .B(KEYINPUT41), .Z(new_n1012));
  INV_X1    g0812(.A(KEYINPUT44), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n989), .B2(new_n738), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n731), .A2(new_n984), .B1(new_n673), .B2(new_n723), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n983), .A2(KEYINPUT44), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT45), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n983), .B2(new_n1015), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n989), .A2(new_n738), .A3(KEYINPUT45), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n734), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1017), .A2(new_n1021), .A3(new_n734), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1024), .B1(new_n1026), .B2(KEYINPUT110), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n730), .A2(KEYINPUT111), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n733), .A2(new_n736), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT111), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n778), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n986), .A4(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n986), .B1(new_n733), .B2(new_n736), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1033), .A2(KEYINPUT111), .A3(new_n730), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT110), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1022), .A2(new_n1036), .A3(new_n1023), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1027), .A2(new_n774), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1012), .B1(new_n1038), .B2(new_n774), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1011), .B1(new_n1039), .B2(new_n782), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n816), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(G97), .ZN(new_n1042));
  INV_X1    g0842(.A(G317), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n331), .C1(new_n1043), .C2(new_n828), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT112), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT46), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n820), .B2(new_n557), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n819), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(new_n806), .C2(new_n663), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1044), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n1045), .B2(new_n1049), .C1(new_n817), .C2(new_n850), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n832), .A2(G107), .B1(G311), .B2(new_n834), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n548), .B2(new_n803), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n831), .A2(new_n372), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G143), .B2(new_n834), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n872), .B2(new_n803), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1041), .A2(G77), .B1(new_n829), .B2(G137), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n268), .B1(new_n820), .B2(new_n278), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G159), .B2(new_n807), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1057), .B(new_n1059), .C1(new_n202), .C2(new_n850), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1051), .A2(new_n1053), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT47), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n797), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n235), .A2(new_n794), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n799), .B1(new_n740), .B2(new_n342), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n784), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n788), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1063), .B(new_n1066), .C1(new_n1067), .C2(new_n1000), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1040), .A2(new_n1068), .ZN(G387));
  OR3_X1    g0869(.A1(new_n774), .A2(KEYINPUT116), .A3(new_n1035), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1035), .A2(new_n754), .A3(new_n773), .ZN(new_n1071));
  OAI21_X1  g0871(.A(KEYINPUT116), .B1(new_n774), .B2(new_n1035), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1070), .A2(new_n741), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n733), .A2(new_n1067), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n743), .A2(new_n740), .A3(new_n331), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n222), .B2(new_n740), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT113), .Z(new_n1078));
  NAND2_X1  g0878(.A1(new_n339), .A2(new_n202), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT50), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n743), .B(new_n250), .C1(new_n372), .C2(new_n205), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n793), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n239), .A2(new_n250), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1078), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n784), .B(new_n1075), .C1(new_n798), .C2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1042), .B(new_n268), .C1(new_n205), .C2(new_n820), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G50), .B2(new_n804), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n828), .A2(new_n872), .B1(new_n372), .B2(new_n823), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n411), .B2(new_n807), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n831), .A2(new_n341), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G159), .B2(new_n834), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n803), .A2(new_n1043), .B1(new_n806), .B2(new_n821), .ZN(new_n1093));
  XOR2_X1   g0893(.A(KEYINPUT114), .B(G322), .Z(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n834), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n850), .B2(new_n548), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT48), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n831), .A2(new_n817), .B1(new_n663), .B2(new_n820), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(KEYINPUT49), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n268), .B1(new_n829), .B2(G326), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(new_n557), .C2(new_n816), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT49), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1092), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT115), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1107), .A2(new_n797), .A3(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1085), .A2(new_n1109), .B1(new_n782), .B2(new_n1035), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1073), .A2(new_n1110), .ZN(G393));
  NAND2_X1  g0911(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n1071), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1038), .A2(new_n741), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1024), .A2(new_n782), .A3(new_n1025), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n244), .A2(new_n794), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n798), .B1(new_n471), .B2(new_n209), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n783), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n829), .A2(new_n1094), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n548), .B2(new_n806), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G294), .B2(new_n847), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n268), .B(new_n840), .C1(G283), .C2(new_n819), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(new_n557), .C2(new_n831), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n821), .A2(new_n803), .B1(new_n833), .B2(new_n1043), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1124), .B(KEYINPUT52), .Z(new_n1125));
  AOI211_X1 g0925(.A(new_n331), .B(new_n883), .C1(G68), .C2(new_n819), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n874), .A2(new_n339), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n831), .A2(new_n205), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n829), .A2(G143), .B1(G50), .B2(new_n807), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n872), .A2(new_n833), .B1(new_n803), .B2(new_n844), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT51), .Z(new_n1133));
  OAI22_X1  g0933(.A1(new_n1123), .A2(new_n1125), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1118), .B1(new_n1134), .B2(new_n797), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n989), .B2(new_n1067), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1115), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(KEYINPUT117), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT117), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1115), .A2(new_n1139), .A3(new_n1136), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1114), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(G390));
  AOI21_X1  g0943(.A(new_n929), .B1(new_n772), .B2(new_n862), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n716), .B(new_n964), .C1(new_n757), .C2(new_n966), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n909), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(G330), .B(new_n862), .C1(new_n957), .C2(new_n960), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n928), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n772), .A2(new_n862), .A3(new_n929), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n749), .A2(new_n724), .A3(new_n862), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n908), .A4(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1146), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n970), .A2(G330), .A3(new_n467), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n750), .A2(new_n467), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n707), .A2(new_n709), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT94), .B1(new_n705), .B2(new_n706), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n612), .B(new_n699), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT29), .B1(new_n1157), .B2(new_n724), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n690), .B(new_n1153), .C1(new_n1154), .C2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT118), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n904), .A2(KEYINPUT118), .A3(new_n690), .A4(new_n1153), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1152), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n863), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n907), .B1(new_n1157), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n950), .B1(new_n1165), .B2(new_n928), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n949), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1150), .A2(new_n908), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n929), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n950), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n948), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1167), .A2(new_n1172), .A3(new_n1149), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1145), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n1167), .B2(new_n1172), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1163), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n741), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT119), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1167), .A2(new_n1172), .A3(new_n1149), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1166), .A2(new_n949), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1179), .B1(new_n1180), .B2(new_n1174), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1178), .B1(new_n1181), .B2(new_n1163), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1152), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1167), .A2(new_n1172), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n1145), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1183), .A2(KEYINPUT119), .A3(new_n1179), .A4(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1177), .B1(new_n1182), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n783), .B1(new_n411), .B2(new_n868), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n819), .A2(G150), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT53), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n331), .B(new_n1190), .C1(G132), .C2(new_n804), .ZN(new_n1191));
  XOR2_X1   g0991(.A(KEYINPUT54), .B(G143), .Z(new_n1192));
  NAND2_X1  g0992(.A1(new_n874), .A2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n832), .A2(G159), .B1(G128), .B2(new_n834), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n816), .A2(new_n202), .B1(new_n871), .B2(new_n806), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G125), .B2(new_n829), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .A4(new_n1196), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1129), .B1(new_n557), .B2(new_n803), .C1(new_n817), .C2(new_n833), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n878), .A2(new_n268), .A3(new_n842), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n829), .A2(G294), .B1(G107), .B2(new_n807), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(new_n471), .C2(new_n850), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1197), .B1(new_n1198), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1188), .B1(new_n1202), .B2(new_n797), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n932), .A2(new_n934), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n948), .A2(new_n935), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1203), .B1(new_n1206), .B2(new_n787), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1181), .B2(new_n781), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1187), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(G378));
  INV_X1    g1010(.A(KEYINPUT123), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n308), .A2(new_n316), .A3(KEYINPUT10), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n320), .B1(new_n319), .B2(new_n323), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n305), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n302), .A2(new_n915), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n325), .A2(new_n1215), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1219), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n716), .B(new_n1222), .C1(new_n962), .C2(new_n968), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1222), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n969), .B2(G330), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n951), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n946), .A2(new_n947), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n921), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n967), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1229), .A2(KEYINPUT40), .B1(new_n967), .B2(new_n963), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1222), .B1(new_n1230), .B2(new_n716), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n969), .A2(G330), .A3(new_n1224), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n684), .A2(new_n915), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1206), .B2(new_n1170), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1231), .A2(new_n1232), .B1(new_n1234), .B2(new_n930), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1211), .B1(new_n1226), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n951), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1231), .A2(new_n1234), .A3(new_n930), .A4(new_n1232), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1238), .A3(KEYINPUT123), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n782), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1222), .A2(new_n786), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n783), .B1(G50), .B2(new_n868), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1054), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n807), .A2(G97), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n331), .A2(new_n249), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G77), .B2(new_n819), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n823), .A2(new_n341), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n816), .A2(new_n278), .B1(new_n828), .B2(new_n817), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n803), .A2(new_n222), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1249), .B(new_n1250), .C1(KEYINPUT120), .C2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(KEYINPUT120), .B2(new_n1251), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1248), .B(new_n1253), .C1(G116), .C2(new_n834), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1254), .A2(KEYINPUT58), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n819), .A2(new_n1192), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n823), .B2(new_n871), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G125), .A2(new_n834), .B1(new_n804), .B2(G128), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n872), .B2(new_n831), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1257), .B(new_n1259), .C1(G132), .C2(new_n807), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1261), .A2(KEYINPUT59), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(KEYINPUT59), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1041), .A2(G159), .ZN(new_n1264));
  AOI211_X1 g1064(.A(G33), .B(G41), .C1(new_n829), .C2(G124), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1254), .A2(KEYINPUT58), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1246), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1255), .A2(new_n1266), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1243), .B1(new_n1269), .B2(new_n797), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1242), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT121), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1271), .B(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(KEYINPUT122), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1182), .A2(new_n1186), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(KEYINPUT124), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT57), .B1(new_n1279), .B2(new_n1240), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1277), .B1(new_n1182), .B2(new_n1186), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT57), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n741), .B1(new_n1281), .B2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1241), .B(new_n1274), .C1(new_n1280), .C2(new_n1285), .ZN(G375));
  INV_X1    g1086(.A(new_n1152), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1276), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1012), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n1289), .A3(new_n1163), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n928), .A2(new_n786), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n783), .B1(G68), .B2(new_n868), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n834), .A2(G294), .B1(new_n807), .B2(G116), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(new_n850), .B2(new_n222), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1294), .B(KEYINPUT125), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n268), .B1(new_n819), .B2(G97), .ZN(new_n1296));
  OAI221_X1 g1096(.A(new_n1296), .B1(new_n828), .B2(new_n548), .C1(new_n816), .C2(new_n205), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n1090), .B(new_n1297), .C1(G283), .C2(new_n804), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n834), .A2(G132), .ZN(new_n1300));
  XOR2_X1   g1100(.A(new_n1300), .B(KEYINPUT126), .Z(new_n1301));
  OAI21_X1  g1101(.A(new_n268), .B1(new_n820), .B2(new_n844), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n803), .A2(new_n871), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n1302), .B(new_n1303), .C1(new_n1041), .C2(G58), .ZN(new_n1304));
  INV_X1    g1104(.A(G128), .ZN(new_n1305));
  OAI22_X1  g1105(.A1(new_n828), .A2(new_n1305), .B1(new_n872), .B2(new_n823), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(new_n807), .B2(new_n1192), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1304), .B(new_n1307), .C1(new_n202), .C2(new_n831), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1299), .B1(new_n1301), .B2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1292), .B1(new_n1309), .B2(new_n797), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(new_n1152), .A2(new_n782), .B1(new_n1291), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1290), .A2(new_n1311), .ZN(G381));
  NAND2_X1  g1112(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1274), .B1(new_n1313), .B2(new_n781), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n742), .B1(new_n1279), .B2(new_n1283), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1282), .B1(new_n1281), .B2(new_n1313), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1314), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1040), .A2(new_n1142), .A3(new_n1068), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1073), .A2(new_n855), .A3(new_n1110), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1319), .A2(G381), .A3(G384), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1317), .A2(new_n1209), .A3(new_n1318), .A4(new_n1320), .ZN(G407));
  NAND2_X1  g1121(.A1(new_n1317), .A2(new_n1209), .ZN(new_n1322));
  OAI211_X1 g1122(.A(G407), .B(G213), .C1(G343), .C2(new_n1322), .ZN(G409));
  NAND2_X1  g1123(.A1(G393), .A2(G396), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1319), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1142), .B1(new_n1040), .B2(new_n1068), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1326), .B1(new_n1318), .B2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(G387), .A2(G390), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1040), .A2(new_n1142), .A3(new_n1068), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1329), .A2(new_n1330), .A3(new_n1325), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1328), .A2(new_n1331), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n722), .A2(G213), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n782), .B1(new_n1226), .B2(new_n1235), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1273), .ZN(new_n1335));
  NOR3_X1   g1135(.A1(new_n1187), .A2(new_n1208), .A3(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1279), .A2(new_n1240), .A3(new_n1289), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1333), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1338), .B1(new_n1317), .B2(new_n1209), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1288), .A2(KEYINPUT60), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT60), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1276), .A2(new_n1287), .A3(new_n1341), .ZN(new_n1342));
  AOI211_X1 g1142(.A(new_n742), .B(new_n1183), .C1(new_n1340), .C2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1311), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n891), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1340), .A2(new_n1342), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1346), .A2(new_n741), .A3(new_n1163), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1347), .A2(G384), .A3(new_n1311), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1333), .A2(G2897), .ZN(new_n1349));
  AND3_X1   g1149(.A1(new_n1345), .A2(new_n1348), .A3(new_n1349), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1349), .B1(new_n1345), .B2(new_n1348), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  AOI211_X1 g1152(.A(KEYINPUT61), .B(new_n1332), .C1(new_n1339), .C2(new_n1352), .ZN(new_n1353));
  AND2_X1   g1153(.A1(new_n1345), .A2(new_n1348), .ZN(new_n1354));
  OAI211_X1 g1154(.A(new_n1338), .B(new_n1354), .C1(new_n1317), .C2(new_n1209), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT63), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1357), .A2(KEYINPUT127), .ZN(new_n1358));
  OR2_X1    g1158(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1359));
  INV_X1    g1159(.A(KEYINPUT127), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1355), .A2(new_n1360), .A3(new_n1356), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1353), .A2(new_n1358), .A3(new_n1359), .A4(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(KEYINPUT61), .B1(new_n1339), .B2(new_n1352), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(G375), .A2(G378), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT62), .ZN(new_n1365));
  NAND4_X1  g1165(.A1(new_n1364), .A2(new_n1365), .A3(new_n1338), .A4(new_n1354), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1355), .A2(KEYINPUT62), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1363), .A2(new_n1366), .A3(new_n1367), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1368), .A2(new_n1332), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1362), .A2(new_n1369), .ZN(G405));
  NAND2_X1  g1170(.A1(new_n1364), .A2(new_n1322), .ZN(new_n1371));
  INV_X1    g1171(.A(new_n1332), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1371), .A2(new_n1372), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1364), .A2(new_n1322), .A3(new_n1332), .ZN(new_n1374));
  AND3_X1   g1174(.A1(new_n1373), .A2(new_n1354), .A3(new_n1374), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1354), .B1(new_n1373), .B2(new_n1374), .ZN(new_n1376));
  NOR2_X1   g1176(.A1(new_n1375), .A2(new_n1376), .ZN(G402));
endmodule


