

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(n702), .A2(n1003), .ZN(n697) );
  OR2_X1 U550 ( .A1(n737), .A2(n736), .ZN(n738) );
  BUF_X1 U551 ( .A(n688), .Z(G164) );
  NOR2_X2 U552 ( .A1(G2105), .A2(n534), .ZN(n897) );
  INV_X2 U553 ( .A(G2104), .ZN(n534) );
  AND2_X1 U554 ( .A1(G138), .A2(n900), .ZN(n565) );
  NOR2_X1 U555 ( .A1(n539), .A2(n538), .ZN(G160) );
  AND2_X1 U556 ( .A1(G102), .A2(n897), .ZN(n517) );
  XOR2_X1 U557 ( .A(KEYINPUT14), .B(n591), .Z(n518) );
  OR2_X1 U558 ( .A1(n1008), .A2(n696), .ZN(n702) );
  NOR2_X1 U559 ( .A1(G1966), .A2(n779), .ZN(n751) );
  NAND2_X1 U560 ( .A1(n798), .A2(n689), .ZN(n720) );
  NAND2_X1 U561 ( .A1(G8), .A2(n720), .ZN(n779) );
  NOR2_X1 U562 ( .A1(n567), .A2(n517), .ZN(n568) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n533) );
  XNOR2_X1 U564 ( .A(n535), .B(KEYINPUT65), .ZN(n893) );
  AND2_X1 U565 ( .A1(n571), .A2(n570), .ZN(n688) );
  XOR2_X1 U566 ( .A(KEYINPUT69), .B(n529), .Z(G171) );
  XOR2_X1 U567 ( .A(G543), .B(KEYINPUT0), .Z(n639) );
  NOR2_X1 U568 ( .A1(G651), .A2(n639), .ZN(n651) );
  NAND2_X1 U569 ( .A1(n651), .A2(G52), .ZN(n521) );
  XOR2_X1 U570 ( .A(G651), .B(KEYINPUT66), .Z(n522) );
  NOR2_X1 U571 ( .A1(G543), .A2(n522), .ZN(n519) );
  XOR2_X2 U572 ( .A(KEYINPUT1), .B(n519), .Z(n658) );
  NAND2_X1 U573 ( .A1(G64), .A2(n658), .ZN(n520) );
  NAND2_X1 U574 ( .A1(n521), .A2(n520), .ZN(n528) );
  NOR2_X2 U575 ( .A1(n639), .A2(n522), .ZN(n654) );
  NAND2_X1 U576 ( .A1(G77), .A2(n654), .ZN(n523) );
  XNOR2_X1 U577 ( .A(n523), .B(KEYINPUT68), .ZN(n525) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n650) );
  NAND2_X1 U579 ( .A1(G90), .A2(n650), .ZN(n524) );
  NAND2_X1 U580 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U581 ( .A(KEYINPUT9), .B(n526), .Z(n527) );
  NOR2_X1 U582 ( .A1(n528), .A2(n527), .ZN(n529) );
  AND2_X1 U583 ( .A1(G2105), .A2(G2104), .ZN(n891) );
  NAND2_X1 U584 ( .A1(n891), .A2(G113), .ZN(n532) );
  NAND2_X1 U585 ( .A1(G101), .A2(n897), .ZN(n530) );
  XOR2_X1 U586 ( .A(KEYINPUT23), .B(n530), .Z(n531) );
  NAND2_X1 U587 ( .A1(n532), .A2(n531), .ZN(n539) );
  XOR2_X2 U588 ( .A(KEYINPUT17), .B(n533), .Z(n900) );
  NAND2_X1 U589 ( .A1(G137), .A2(n900), .ZN(n537) );
  NAND2_X1 U590 ( .A1(n534), .A2(G2105), .ZN(n535) );
  NAND2_X1 U591 ( .A1(G125), .A2(n893), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U593 ( .A(G2446), .B(G2430), .Z(n541) );
  XNOR2_X1 U594 ( .A(G2451), .B(KEYINPUT106), .ZN(n540) );
  XNOR2_X1 U595 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U596 ( .A(n542), .B(G2427), .Z(n544) );
  XNOR2_X1 U597 ( .A(G1341), .B(G1348), .ZN(n543) );
  XNOR2_X1 U598 ( .A(n544), .B(n543), .ZN(n548) );
  XOR2_X1 U599 ( .A(G2443), .B(G2435), .Z(n546) );
  XNOR2_X1 U600 ( .A(G2438), .B(G2454), .ZN(n545) );
  XNOR2_X1 U601 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U602 ( .A(n548), .B(n547), .Z(n549) );
  AND2_X1 U603 ( .A1(G14), .A2(n549), .ZN(G401) );
  AND2_X1 U604 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U605 ( .A1(G111), .A2(n891), .ZN(n551) );
  NAND2_X1 U606 ( .A1(G99), .A2(n897), .ZN(n550) );
  NAND2_X1 U607 ( .A1(n551), .A2(n550), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n893), .A2(G123), .ZN(n552) );
  XOR2_X1 U609 ( .A(KEYINPUT18), .B(n552), .Z(n553) );
  NOR2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n900), .A2(G135), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n975) );
  XNOR2_X1 U613 ( .A(G2096), .B(n975), .ZN(n557) );
  OR2_X1 U614 ( .A1(G2100), .A2(n557), .ZN(G156) );
  NAND2_X1 U615 ( .A1(n651), .A2(G53), .ZN(n559) );
  NAND2_X1 U616 ( .A1(G65), .A2(n658), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U618 ( .A1(G91), .A2(n650), .ZN(n561) );
  NAND2_X1 U619 ( .A1(G78), .A2(n654), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U621 ( .A1(n563), .A2(n562), .ZN(n712) );
  INV_X1 U622 ( .A(n712), .ZN(G299) );
  INV_X1 U623 ( .A(KEYINPUT88), .ZN(n564) );
  XNOR2_X1 U624 ( .A(n565), .B(n564), .ZN(n571) );
  NAND2_X1 U625 ( .A1(G126), .A2(n893), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G114), .A2(n891), .ZN(n566) );
  XNOR2_X1 U627 ( .A(KEYINPUT87), .B(n566), .ZN(n567) );
  AND2_X1 U628 ( .A1(n569), .A2(n568), .ZN(n570) );
  INV_X1 U629 ( .A(G120), .ZN(G236) );
  INV_X1 U630 ( .A(G69), .ZN(G235) );
  INV_X1 U631 ( .A(G108), .ZN(G238) );
  NAND2_X1 U632 ( .A1(n650), .A2(G89), .ZN(n573) );
  XNOR2_X1 U633 ( .A(n573), .B(KEYINPUT4), .ZN(n575) );
  NAND2_X1 U634 ( .A1(G76), .A2(n654), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U636 ( .A(n576), .B(KEYINPUT5), .ZN(n581) );
  NAND2_X1 U637 ( .A1(n651), .A2(G51), .ZN(n578) );
  NAND2_X1 U638 ( .A1(G63), .A2(n658), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U640 ( .A(KEYINPUT6), .B(n579), .Z(n580) );
  NAND2_X1 U641 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U642 ( .A(n582), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U643 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U644 ( .A1(G7), .A2(G661), .ZN(n583) );
  XNOR2_X1 U645 ( .A(n583), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U646 ( .A(G223), .ZN(n834) );
  NAND2_X1 U647 ( .A1(n834), .A2(G567), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT11), .B(n584), .Z(G234) );
  XOR2_X1 U649 ( .A(G860), .B(KEYINPUT72), .Z(n608) );
  XNOR2_X1 U650 ( .A(KEYINPUT71), .B(KEYINPUT13), .ZN(n590) );
  NAND2_X1 U651 ( .A1(G81), .A2(n650), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n585), .B(KEYINPUT70), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n586), .B(KEYINPUT12), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G68), .A2(n654), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U656 ( .A(n590), .B(n589), .ZN(n592) );
  NAND2_X1 U657 ( .A1(G56), .A2(n658), .ZN(n591) );
  NOR2_X1 U658 ( .A1(n592), .A2(n518), .ZN(n594) );
  NAND2_X1 U659 ( .A1(n651), .A2(G43), .ZN(n593) );
  NAND2_X1 U660 ( .A1(n594), .A2(n593), .ZN(n1008) );
  OR2_X1 U661 ( .A1(n608), .A2(n1008), .ZN(G153) );
  NAND2_X1 U662 ( .A1(G868), .A2(G171), .ZN(n603) );
  NAND2_X1 U663 ( .A1(n651), .A2(G54), .ZN(n596) );
  NAND2_X1 U664 ( .A1(G66), .A2(n658), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U666 ( .A1(G92), .A2(n650), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G79), .A2(n654), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U669 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U670 ( .A(n601), .B(KEYINPUT15), .ZN(n1003) );
  INV_X1 U671 ( .A(n1003), .ZN(n616) );
  INV_X1 U672 ( .A(G868), .ZN(n669) );
  NAND2_X1 U673 ( .A1(n616), .A2(n669), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U675 ( .A(n604), .B(KEYINPUT73), .ZN(G284) );
  NOR2_X1 U676 ( .A1(G286), .A2(n669), .ZN(n606) );
  NOR2_X1 U677 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U679 ( .A(KEYINPUT74), .B(n607), .ZN(G297) );
  NAND2_X1 U680 ( .A1(G559), .A2(n608), .ZN(n609) );
  XOR2_X1 U681 ( .A(KEYINPUT75), .B(n609), .Z(n610) );
  NAND2_X1 U682 ( .A1(n610), .A2(n616), .ZN(n611) );
  XNOR2_X1 U683 ( .A(n611), .B(KEYINPUT16), .ZN(n612) );
  XNOR2_X1 U684 ( .A(KEYINPUT76), .B(n612), .ZN(G148) );
  NOR2_X1 U685 ( .A1(G868), .A2(n1008), .ZN(n615) );
  NAND2_X1 U686 ( .A1(G868), .A2(n616), .ZN(n613) );
  NOR2_X1 U687 ( .A1(G559), .A2(n613), .ZN(n614) );
  NOR2_X1 U688 ( .A1(n615), .A2(n614), .ZN(G282) );
  XNOR2_X1 U689 ( .A(n1008), .B(KEYINPUT77), .ZN(n618) );
  NAND2_X1 U690 ( .A1(n616), .A2(G559), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n618), .B(n617), .ZN(n667) );
  XOR2_X1 U692 ( .A(n667), .B(KEYINPUT78), .Z(n619) );
  NOR2_X1 U693 ( .A1(G860), .A2(n619), .ZN(n627) );
  NAND2_X1 U694 ( .A1(G93), .A2(n650), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G55), .A2(n651), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U697 ( .A1(G80), .A2(n654), .ZN(n622) );
  XNOR2_X1 U698 ( .A(KEYINPUT79), .B(n622), .ZN(n623) );
  NOR2_X1 U699 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U700 ( .A1(G67), .A2(n658), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n670) );
  XOR2_X1 U702 ( .A(n627), .B(n670), .Z(G145) );
  NAND2_X1 U703 ( .A1(G85), .A2(n650), .ZN(n629) );
  NAND2_X1 U704 ( .A1(G72), .A2(n654), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U706 ( .A1(G60), .A2(n658), .ZN(n630) );
  XNOR2_X1 U707 ( .A(KEYINPUT67), .B(n630), .ZN(n631) );
  NOR2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n651), .A2(G47), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(G290) );
  NAND2_X1 U711 ( .A1(G49), .A2(n651), .ZN(n636) );
  NAND2_X1 U712 ( .A1(G74), .A2(G651), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U714 ( .A(KEYINPUT80), .B(n637), .ZN(n638) );
  NOR2_X1 U715 ( .A1(n658), .A2(n638), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n639), .A2(G87), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(G288) );
  NAND2_X1 U718 ( .A1(G75), .A2(n654), .ZN(n642) );
  XOR2_X1 U719 ( .A(KEYINPUT81), .B(n642), .Z(n644) );
  NAND2_X1 U720 ( .A1(n650), .A2(G88), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U722 ( .A(KEYINPUT82), .B(n645), .ZN(n649) );
  NAND2_X1 U723 ( .A1(n651), .A2(G50), .ZN(n647) );
  NAND2_X1 U724 ( .A1(G62), .A2(n658), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U726 ( .A1(n649), .A2(n648), .ZN(G166) );
  NAND2_X1 U727 ( .A1(G86), .A2(n650), .ZN(n653) );
  NAND2_X1 U728 ( .A1(G48), .A2(n651), .ZN(n652) );
  NAND2_X1 U729 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U730 ( .A1(n654), .A2(G73), .ZN(n655) );
  XOR2_X1 U731 ( .A(KEYINPUT2), .B(n655), .Z(n656) );
  NOR2_X1 U732 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U733 ( .A1(G61), .A2(n658), .ZN(n659) );
  NAND2_X1 U734 ( .A1(n660), .A2(n659), .ZN(G305) );
  XNOR2_X1 U735 ( .A(n712), .B(G290), .ZN(n666) );
  XNOR2_X1 U736 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n662) );
  XNOR2_X1 U737 ( .A(G288), .B(G166), .ZN(n661) );
  XNOR2_X1 U738 ( .A(n662), .B(n661), .ZN(n663) );
  XOR2_X1 U739 ( .A(n663), .B(G305), .Z(n664) );
  XNOR2_X1 U740 ( .A(n670), .B(n664), .ZN(n665) );
  XNOR2_X1 U741 ( .A(n666), .B(n665), .ZN(n908) );
  XNOR2_X1 U742 ( .A(n667), .B(n908), .ZN(n668) );
  NAND2_X1 U743 ( .A1(n668), .A2(G868), .ZN(n672) );
  NAND2_X1 U744 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U745 ( .A1(n672), .A2(n671), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n673) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n673), .Z(n674) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U750 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U752 ( .A1(G235), .A2(G236), .ZN(n677) );
  XNOR2_X1 U753 ( .A(n677), .B(KEYINPUT85), .ZN(n678) );
  NOR2_X1 U754 ( .A1(G238), .A2(n678), .ZN(n679) );
  NAND2_X1 U755 ( .A1(G57), .A2(n679), .ZN(n838) );
  NAND2_X1 U756 ( .A1(G567), .A2(n838), .ZN(n685) );
  NAND2_X1 U757 ( .A1(G132), .A2(G82), .ZN(n680) );
  XNOR2_X1 U758 ( .A(n680), .B(KEYINPUT22), .ZN(n681) );
  XNOR2_X1 U759 ( .A(n681), .B(KEYINPUT84), .ZN(n682) );
  NOR2_X1 U760 ( .A1(G218), .A2(n682), .ZN(n683) );
  NAND2_X1 U761 ( .A1(G96), .A2(n683), .ZN(n839) );
  NAND2_X1 U762 ( .A1(G2106), .A2(n839), .ZN(n684) );
  NAND2_X1 U763 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U764 ( .A(KEYINPUT86), .B(n686), .Z(G319) );
  INV_X1 U765 ( .A(G319), .ZN(n914) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n687) );
  NOR2_X1 U767 ( .A1(n914), .A2(n687), .ZN(n837) );
  NAND2_X1 U768 ( .A1(n837), .A2(G36), .ZN(G176) );
  XNOR2_X1 U769 ( .A(KEYINPUT89), .B(G166), .ZN(G303) );
  XNOR2_X1 U770 ( .A(G1981), .B(G305), .ZN(n1014) );
  NOR2_X2 U771 ( .A1(n688), .A2(G1384), .ZN(n798) );
  NAND2_X1 U772 ( .A1(G160), .A2(G40), .ZN(n797) );
  INV_X1 U773 ( .A(n797), .ZN(n689) );
  INV_X1 U774 ( .A(G1996), .ZN(n690) );
  NOR2_X1 U775 ( .A1(n720), .A2(n690), .ZN(n693) );
  XNOR2_X1 U776 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n691) );
  XNOR2_X1 U777 ( .A(n691), .B(KEYINPUT64), .ZN(n692) );
  XNOR2_X1 U778 ( .A(n693), .B(n692), .ZN(n695) );
  BUF_X2 U779 ( .A(n720), .Z(n726) );
  NAND2_X1 U780 ( .A1(n726), .A2(G1341), .ZN(n694) );
  NAND2_X1 U781 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U782 ( .A(n697), .B(KEYINPUT96), .Z(n701) );
  INV_X1 U783 ( .A(n726), .ZN(n717) );
  NOR2_X1 U784 ( .A1(n717), .A2(G1348), .ZN(n699) );
  NOR2_X1 U785 ( .A1(G2067), .A2(n726), .ZN(n698) );
  NOR2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U787 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U788 ( .A1(n702), .A2(n1003), .ZN(n703) );
  NAND2_X1 U789 ( .A1(n704), .A2(n703), .ZN(n710) );
  NAND2_X1 U790 ( .A1(n717), .A2(G2072), .ZN(n705) );
  XNOR2_X1 U791 ( .A(KEYINPUT27), .B(n705), .ZN(n708) );
  NAND2_X1 U792 ( .A1(G1956), .A2(n726), .ZN(n706) );
  XOR2_X1 U793 ( .A(KEYINPUT94), .B(n706), .Z(n707) );
  NOR2_X1 U794 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U795 ( .A1(n712), .A2(n711), .ZN(n709) );
  NAND2_X1 U796 ( .A1(n710), .A2(n709), .ZN(n715) );
  NOR2_X1 U797 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U798 ( .A(n713), .B(KEYINPUT28), .Z(n714) );
  NAND2_X1 U799 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U800 ( .A(n716), .B(KEYINPUT29), .ZN(n747) );
  XNOR2_X1 U801 ( .A(KEYINPUT25), .B(G2078), .ZN(n952) );
  NOR2_X1 U802 ( .A1(n726), .A2(n952), .ZN(n719) );
  INV_X1 U803 ( .A(G1961), .ZN(n923) );
  NOR2_X1 U804 ( .A1(n717), .A2(n923), .ZN(n718) );
  NOR2_X1 U805 ( .A1(n719), .A2(n718), .ZN(n730) );
  AND2_X1 U806 ( .A1(G171), .A2(n730), .ZN(n746) );
  NOR2_X1 U807 ( .A1(G1971), .A2(n779), .ZN(n722) );
  NOR2_X1 U808 ( .A1(G2090), .A2(n726), .ZN(n721) );
  NOR2_X1 U809 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U810 ( .A1(n723), .A2(G303), .ZN(n735) );
  INV_X1 U811 ( .A(n735), .ZN(n724) );
  NOR2_X1 U812 ( .A1(n724), .A2(G286), .ZN(n737) );
  OR2_X1 U813 ( .A1(n746), .A2(n737), .ZN(n725) );
  OR2_X1 U814 ( .A1(n747), .A2(n725), .ZN(n739) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n726), .ZN(n744) );
  NOR2_X1 U816 ( .A1(n751), .A2(n744), .ZN(n727) );
  NAND2_X1 U817 ( .A1(G8), .A2(n727), .ZN(n728) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n728), .ZN(n729) );
  NOR2_X1 U819 ( .A1(G168), .A2(n729), .ZN(n732) );
  NOR2_X1 U820 ( .A1(G171), .A2(n730), .ZN(n731) );
  NOR2_X1 U821 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U822 ( .A(n733), .B(KEYINPUT97), .ZN(n734) );
  XNOR2_X1 U823 ( .A(n734), .B(KEYINPUT31), .ZN(n748) );
  AND2_X1 U824 ( .A1(n748), .A2(n735), .ZN(n736) );
  NAND2_X1 U825 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U826 ( .A(n740), .B(KEYINPUT98), .ZN(n741) );
  NAND2_X1 U827 ( .A1(n741), .A2(G8), .ZN(n743) );
  XOR2_X1 U828 ( .A(KEYINPUT32), .B(KEYINPUT99), .Z(n742) );
  XNOR2_X1 U829 ( .A(n743), .B(n742), .ZN(n755) );
  NAND2_X1 U830 ( .A1(G8), .A2(n744), .ZN(n745) );
  XOR2_X1 U831 ( .A(KEYINPUT93), .B(n745), .Z(n753) );
  OR2_X1 U832 ( .A1(n747), .A2(n746), .ZN(n749) );
  AND2_X1 U833 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U834 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U835 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U836 ( .A1(n755), .A2(n754), .ZN(n769) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n763) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U839 ( .A1(n763), .A2(n756), .ZN(n1016) );
  NAND2_X1 U840 ( .A1(n769), .A2(n1016), .ZN(n757) );
  XNOR2_X1 U841 ( .A(n757), .B(KEYINPUT100), .ZN(n760) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n1001) );
  INV_X1 U843 ( .A(n1001), .ZN(n758) );
  NOR2_X1 U844 ( .A1(n779), .A2(n758), .ZN(n759) );
  AND2_X1 U845 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U846 ( .A1(n761), .A2(KEYINPUT33), .ZN(n762) );
  NOR2_X1 U847 ( .A1(n1014), .A2(n762), .ZN(n768) );
  NAND2_X1 U848 ( .A1(KEYINPUT33), .A2(n763), .ZN(n764) );
  XOR2_X1 U849 ( .A(KEYINPUT101), .B(n764), .Z(n765) );
  NOR2_X1 U850 ( .A1(n779), .A2(n765), .ZN(n766) );
  XOR2_X1 U851 ( .A(KEYINPUT102), .B(n766), .Z(n767) );
  NAND2_X1 U852 ( .A1(n768), .A2(n767), .ZN(n775) );
  NOR2_X1 U853 ( .A1(G2090), .A2(G303), .ZN(n770) );
  NAND2_X1 U854 ( .A1(G8), .A2(n770), .ZN(n771) );
  NAND2_X1 U855 ( .A1(n769), .A2(n771), .ZN(n772) );
  NAND2_X1 U856 ( .A1(n779), .A2(n772), .ZN(n773) );
  XOR2_X1 U857 ( .A(KEYINPUT103), .B(n773), .Z(n774) );
  NAND2_X1 U858 ( .A1(n775), .A2(n774), .ZN(n822) );
  NOR2_X1 U859 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U860 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  XNOR2_X1 U861 ( .A(KEYINPUT92), .B(n777), .ZN(n778) );
  NOR2_X1 U862 ( .A1(n779), .A2(n778), .ZN(n820) );
  XOR2_X1 U863 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n804) );
  NAND2_X1 U864 ( .A1(G117), .A2(n891), .ZN(n781) );
  NAND2_X1 U865 ( .A1(G129), .A2(n893), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U867 ( .A1(n897), .A2(G105), .ZN(n782) );
  XOR2_X1 U868 ( .A(KEYINPUT38), .B(n782), .Z(n783) );
  NOR2_X1 U869 ( .A1(n784), .A2(n783), .ZN(n786) );
  NAND2_X1 U870 ( .A1(n900), .A2(G141), .ZN(n785) );
  NAND2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n879) );
  NOR2_X1 U872 ( .A1(n879), .A2(G1996), .ZN(n787) );
  XNOR2_X1 U873 ( .A(n787), .B(KEYINPUT104), .ZN(n982) );
  NAND2_X1 U874 ( .A1(G95), .A2(n897), .ZN(n789) );
  NAND2_X1 U875 ( .A1(G119), .A2(n893), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U877 ( .A1(G107), .A2(n891), .ZN(n790) );
  XNOR2_X1 U878 ( .A(KEYINPUT91), .B(n790), .ZN(n791) );
  NOR2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U880 ( .A1(n900), .A2(G131), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n880) );
  AND2_X1 U882 ( .A1(n880), .A2(G1991), .ZN(n796) );
  AND2_X1 U883 ( .A1(n879), .A2(G1996), .ZN(n795) );
  NOR2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n980) );
  NOR2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n826) );
  INV_X1 U886 ( .A(n826), .ZN(n799) );
  NOR2_X1 U887 ( .A1(n980), .A2(n799), .ZN(n823) );
  NOR2_X1 U888 ( .A1(G1991), .A2(n880), .ZN(n978) );
  NOR2_X1 U889 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NOR2_X1 U890 ( .A1(n978), .A2(n800), .ZN(n801) );
  NOR2_X1 U891 ( .A1(n823), .A2(n801), .ZN(n802) );
  NOR2_X1 U892 ( .A1(n982), .A2(n802), .ZN(n803) );
  XNOR2_X1 U893 ( .A(n804), .B(n803), .ZN(n815) );
  XNOR2_X1 U894 ( .A(G2067), .B(KEYINPUT37), .ZN(n816) );
  XNOR2_X1 U895 ( .A(KEYINPUT90), .B(KEYINPUT34), .ZN(n808) );
  NAND2_X1 U896 ( .A1(G140), .A2(n900), .ZN(n806) );
  NAND2_X1 U897 ( .A1(G104), .A2(n897), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U899 ( .A(n808), .B(n807), .ZN(n813) );
  NAND2_X1 U900 ( .A1(G116), .A2(n891), .ZN(n810) );
  NAND2_X1 U901 ( .A1(G128), .A2(n893), .ZN(n809) );
  NAND2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n811) );
  XOR2_X1 U903 ( .A(KEYINPUT35), .B(n811), .Z(n812) );
  NOR2_X1 U904 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U905 ( .A(KEYINPUT36), .B(n814), .ZN(n904) );
  NOR2_X1 U906 ( .A1(n816), .A2(n904), .ZN(n989) );
  NAND2_X1 U907 ( .A1(n826), .A2(n989), .ZN(n824) );
  NAND2_X1 U908 ( .A1(n815), .A2(n824), .ZN(n817) );
  NAND2_X1 U909 ( .A1(n816), .A2(n904), .ZN(n986) );
  NAND2_X1 U910 ( .A1(n817), .A2(n986), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n818), .A2(n826), .ZN(n830) );
  INV_X1 U912 ( .A(n830), .ZN(n819) );
  OR2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n832) );
  INV_X1 U915 ( .A(n823), .ZN(n825) );
  AND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(n828) );
  XNOR2_X1 U917 ( .A(G1986), .B(G290), .ZN(n1000) );
  NAND2_X1 U918 ( .A1(n1000), .A2(n826), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n828), .A2(n827), .ZN(n829) );
  AND2_X1 U920 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U921 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U922 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U925 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U927 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U929 ( .A(G132), .ZN(G219) );
  INV_X1 U930 ( .A(G82), .ZN(G220) );
  NOR2_X1 U931 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  XOR2_X1 U933 ( .A(G1966), .B(G1971), .Z(n841) );
  XNOR2_X1 U934 ( .A(G1986), .B(G1976), .ZN(n840) );
  XNOR2_X1 U935 ( .A(n841), .B(n840), .ZN(n851) );
  XOR2_X1 U936 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n843) );
  XNOR2_X1 U937 ( .A(G1996), .B(G2474), .ZN(n842) );
  XNOR2_X1 U938 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U939 ( .A(G1956), .B(G1961), .Z(n845) );
  XNOR2_X1 U940 ( .A(G1991), .B(G1981), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U942 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U943 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n848) );
  XNOR2_X1 U944 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U945 ( .A(n851), .B(n850), .Z(G229) );
  XOR2_X1 U946 ( .A(G2678), .B(KEYINPUT107), .Z(n853) );
  XNOR2_X1 U947 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n852) );
  XNOR2_X1 U948 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U949 ( .A(KEYINPUT42), .B(G2090), .Z(n855) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U952 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U953 ( .A(G2096), .B(G2100), .ZN(n858) );
  XNOR2_X1 U954 ( .A(n859), .B(n858), .ZN(n861) );
  XOR2_X1 U955 ( .A(G2078), .B(G2084), .Z(n860) );
  XNOR2_X1 U956 ( .A(n861), .B(n860), .ZN(G227) );
  NAND2_X1 U957 ( .A1(n900), .A2(G136), .ZN(n868) );
  NAND2_X1 U958 ( .A1(G112), .A2(n891), .ZN(n863) );
  NAND2_X1 U959 ( .A1(G100), .A2(n897), .ZN(n862) );
  NAND2_X1 U960 ( .A1(n863), .A2(n862), .ZN(n866) );
  NAND2_X1 U961 ( .A1(n893), .A2(G124), .ZN(n864) );
  XOR2_X1 U962 ( .A(KEYINPUT44), .B(n864), .Z(n865) );
  NOR2_X1 U963 ( .A1(n866), .A2(n865), .ZN(n867) );
  NAND2_X1 U964 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U965 ( .A(KEYINPUT112), .B(n869), .Z(G162) );
  NAND2_X1 U966 ( .A1(G142), .A2(n900), .ZN(n871) );
  NAND2_X1 U967 ( .A1(G106), .A2(n897), .ZN(n870) );
  NAND2_X1 U968 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U969 ( .A(n872), .B(KEYINPUT45), .ZN(n874) );
  NAND2_X1 U970 ( .A1(G130), .A2(n893), .ZN(n873) );
  NAND2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n877) );
  NAND2_X1 U972 ( .A1(G118), .A2(n891), .ZN(n875) );
  XNOR2_X1 U973 ( .A(KEYINPUT113), .B(n875), .ZN(n876) );
  NOR2_X1 U974 ( .A1(n877), .A2(n876), .ZN(n890) );
  XNOR2_X1 U975 ( .A(G164), .B(G162), .ZN(n878) );
  XNOR2_X1 U976 ( .A(n878), .B(n975), .ZN(n883) );
  XOR2_X1 U977 ( .A(G160), .B(n879), .Z(n881) );
  XOR2_X1 U978 ( .A(n881), .B(n880), .Z(n882) );
  XOR2_X1 U979 ( .A(n883), .B(n882), .Z(n888) );
  XOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT117), .Z(n885) );
  XNOR2_X1 U981 ( .A(KEYINPUT118), .B(KEYINPUT48), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U983 ( .A(KEYINPUT116), .B(n886), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U985 ( .A(n890), .B(n889), .ZN(n906) );
  NAND2_X1 U986 ( .A1(n891), .A2(G115), .ZN(n892) );
  XOR2_X1 U987 ( .A(KEYINPUT115), .B(n892), .Z(n895) );
  NAND2_X1 U988 ( .A1(n893), .A2(G127), .ZN(n894) );
  NAND2_X1 U989 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U990 ( .A(n896), .B(KEYINPUT47), .ZN(n899) );
  NAND2_X1 U991 ( .A1(G103), .A2(n897), .ZN(n898) );
  NAND2_X1 U992 ( .A1(n899), .A2(n898), .ZN(n903) );
  NAND2_X1 U993 ( .A1(n900), .A2(G139), .ZN(n901) );
  XOR2_X1 U994 ( .A(KEYINPUT114), .B(n901), .Z(n902) );
  NOR2_X1 U995 ( .A1(n903), .A2(n902), .ZN(n971) );
  XNOR2_X1 U996 ( .A(n904), .B(n971), .ZN(n905) );
  XNOR2_X1 U997 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U998 ( .A1(G37), .A2(n907), .ZN(G395) );
  XNOR2_X1 U999 ( .A(G286), .B(n908), .ZN(n911) );
  XNOR2_X1 U1000 ( .A(KEYINPUT119), .B(n1003), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(n909), .B(n1008), .ZN(n910) );
  XNOR2_X1 U1002 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1003 ( .A(n912), .B(G171), .ZN(n913) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n913), .ZN(G397) );
  NOR2_X1 U1005 ( .A1(n914), .A2(G401), .ZN(n915) );
  XOR2_X1 U1006 ( .A(KEYINPUT120), .B(n915), .Z(n919) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n916) );
  XOR2_X1 U1008 ( .A(KEYINPUT121), .B(n916), .Z(n917) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1010 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1011 ( .A(KEYINPUT122), .B(n920), .ZN(n922) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1013 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G96), .ZN(G221) );
  INV_X1 U1016 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1017 ( .A(n923), .B(G5), .ZN(n943) );
  XOR2_X1 U1018 ( .A(G1966), .B(G21), .Z(n934) );
  XOR2_X1 U1019 ( .A(G1981), .B(G6), .Z(n927) );
  XNOR2_X1 U1020 ( .A(G1956), .B(G20), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(G19), .B(G1341), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(KEYINPUT126), .B(n928), .ZN(n931) );
  XOR2_X1 U1025 ( .A(KEYINPUT59), .B(G1348), .Z(n929) );
  XNOR2_X1 U1026 ( .A(G4), .B(n929), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(KEYINPUT60), .B(n932), .ZN(n933) );
  NAND2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n941) );
  XNOR2_X1 U1030 ( .A(G1976), .B(G23), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(G1971), .B(G22), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n938) );
  XOR2_X1 U1033 ( .A(G1986), .B(G24), .Z(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(KEYINPUT58), .B(n939), .ZN(n940) );
  NOR2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(n944), .B(KEYINPUT127), .ZN(n945) );
  XOR2_X1 U1039 ( .A(KEYINPUT61), .B(n945), .Z(n947) );
  XOR2_X1 U1040 ( .A(G16), .B(KEYINPUT125), .Z(n946) );
  NOR2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n970) );
  INV_X1 U1042 ( .A(KEYINPUT55), .ZN(n994) );
  XNOR2_X1 U1043 ( .A(G2090), .B(G35), .ZN(n961) );
  XOR2_X1 U1044 ( .A(G1991), .B(G25), .Z(n948) );
  NAND2_X1 U1045 ( .A1(n948), .A2(G28), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(n949), .B(KEYINPUT124), .ZN(n958) );
  XNOR2_X1 U1047 ( .A(G2067), .B(G26), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(G1996), .B(G32), .ZN(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n956) );
  XOR2_X1 U1050 ( .A(n952), .B(G27), .Z(n954) );
  XNOR2_X1 U1051 ( .A(G2072), .B(G33), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT53), .B(n959), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n964) );
  XOR2_X1 U1057 ( .A(G2084), .B(G34), .Z(n962) );
  XNOR2_X1 U1058 ( .A(KEYINPUT54), .B(n962), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(n994), .B(n965), .ZN(n967) );
  INV_X1 U1061 ( .A(G29), .ZN(n966) );
  NAND2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n968), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n998) );
  XOR2_X1 U1065 ( .A(G2072), .B(n971), .Z(n973) );
  XOR2_X1 U1066 ( .A(G164), .B(G2078), .Z(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1068 ( .A(KEYINPUT50), .B(n974), .Z(n992) );
  XNOR2_X1 U1069 ( .A(G160), .B(G2084), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n985) );
  XOR2_X1 U1073 ( .A(G2090), .B(G162), .Z(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(n983), .B(KEYINPUT51), .ZN(n984) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(KEYINPUT123), .B(n990), .ZN(n991) );
  NOR2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(KEYINPUT52), .B(n993), .ZN(n995) );
  NAND2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n996), .A2(G29), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n1023) );
  XOR2_X1 U1085 ( .A(G16), .B(KEYINPUT56), .Z(n1021) );
  XNOR2_X1 U1086 ( .A(G171), .B(G1961), .ZN(n1012) );
  XNOR2_X1 U1087 ( .A(G1956), .B(G299), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(G1348), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  NAND2_X1 U1092 ( .A1(G1971), .A2(G303), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(G1341), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1096 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XOR2_X1 U1097 ( .A(G1966), .B(G168), .Z(n1013) );
  NOR2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1099 ( .A(KEYINPUT57), .B(n1015), .Z(n1017) );
  NAND2_X1 U1100 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1101 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1102 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1103 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1104 ( .A(n1024), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
  INV_X1 U1106 ( .A(G171), .ZN(G301) );
endmodule

