//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n558, new_n560,
    new_n561, new_n562, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1143, new_n1144, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(new_n455), .B(KEYINPUT66), .Z(G261));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT70), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n468), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n472), .A2(G137), .A3(new_n463), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n467), .A2(new_n474), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  NAND3_X1  g058(.A1(new_n472), .A2(new_n463), .A3(new_n473), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n484), .B(new_n485), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n472), .A2(G2105), .A3(new_n473), .ZN(new_n490));
  INV_X1    g065(.A(G124), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n487), .A2(new_n492), .ZN(G162));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR4_X1   g069(.A1(new_n478), .A2(KEYINPUT4), .A3(new_n494), .A4(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n472), .A2(G138), .A3(new_n463), .A4(new_n473), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n495), .B1(KEYINPUT4), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n463), .A2(G114), .ZN(new_n500));
  OAI22_X1  g075(.A1(new_n490), .A2(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n497), .A2(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G651), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n509), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n504), .A2(KEYINPUT73), .A3(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n508), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n508), .A2(new_n512), .A3(KEYINPUT74), .A4(new_n513), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G88), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n520), .A2(new_n506), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n508), .A2(new_n512), .A3(G543), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n519), .A2(new_n521), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND2_X1  g101(.A1(new_n523), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n516), .A2(G89), .A3(new_n517), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n529), .A2(KEYINPUT75), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(KEYINPUT75), .B1(new_n529), .B2(new_n531), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n527), .B(new_n528), .C1(new_n533), .C2(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND2_X1  g111(.A1(new_n518), .A2(G90), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n523), .A2(G52), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT76), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n537), .A2(new_n538), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT5), .B(G543), .Z(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n547), .A2(KEYINPUT77), .A3(G651), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n550), .B2(new_n506), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n516), .A2(G81), .A3(new_n517), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n523), .A2(G43), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  XOR2_X1   g134(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n560));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(new_n518), .A2(G91), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n522), .A2(new_n565), .B1(KEYINPUT79), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g142(.A(KEYINPUT80), .B(G65), .ZN(new_n568));
  NOR3_X1   g143(.A1(new_n545), .A2(new_n568), .A3(new_n506), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n566), .A2(KEYINPUT79), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n508), .A2(new_n512), .A3(G53), .A4(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G78), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(new_n506), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n569), .B1(new_n573), .B2(G543), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n564), .A2(new_n567), .A3(new_n574), .ZN(G299));
  OAI21_X1  g150(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n523), .A2(G49), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n516), .A2(new_n517), .ZN(new_n578));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(new_n523), .A2(G48), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  OAI221_X1 g158(.A(new_n581), .B1(new_n506), .B2(new_n582), .C1(new_n578), .C2(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(new_n518), .A2(G85), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(new_n506), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n523), .A2(G47), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n516), .A2(G92), .A3(new_n517), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT81), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n516), .A2(new_n594), .A3(G92), .A4(new_n517), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G54), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n522), .A2(new_n599), .B1(new_n600), .B2(new_n506), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT82), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n593), .A2(KEYINPUT10), .A3(new_n595), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n598), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n591), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n591), .B1(new_n605), .B2(G868), .ZN(G321));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G299), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n605), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g192(.A(new_n478), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n466), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  INV_X1    g197(.A(G123), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n463), .A2(G111), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT83), .Z(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  OAI22_X1  g201(.A1(new_n490), .A2(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(new_n486), .B2(G135), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n622), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT84), .Z(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT15), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2435), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(KEYINPUT14), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n636), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(G14), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  XOR2_X1   g222(.A(G2067), .B(G2678), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n647), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2100), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n649), .A2(new_n650), .ZN(new_n656));
  AOI21_X1  g231(.A(KEYINPUT18), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n654), .B(new_n657), .Z(G227));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT86), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n662), .B2(new_n663), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n660), .A2(KEYINPUT87), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n665), .B(new_n666), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(new_n663), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n668), .A2(new_n660), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1981), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G1991), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n671), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT88), .B(G1986), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G229));
  INV_X1    g254(.A(G16), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n680), .A2(G6), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(G305), .B2(G16), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT32), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G1981), .ZN(new_n684));
  NAND2_X1  g259(.A1(G166), .A2(G16), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G16), .B2(G22), .ZN(new_n686));
  INV_X1    g261(.A(G1971), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  OAI21_X1  g264(.A(KEYINPUT90), .B1(G16), .B2(G23), .ZN(new_n690));
  OR3_X1    g265(.A1(KEYINPUT90), .A2(G16), .A3(G23), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n690), .B(new_n691), .C1(G288), .C2(new_n680), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT33), .B(G1976), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  NAND4_X1  g269(.A1(new_n684), .A2(new_n688), .A3(new_n689), .A4(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(KEYINPUT34), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(KEYINPUT34), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT36), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G25), .ZN(new_n701));
  INV_X1    g276(.A(G119), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n463), .A2(G107), .ZN(new_n704));
  OAI22_X1  g279(.A1(new_n490), .A2(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n486), .B2(G131), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n701), .B1(new_n706), .B2(new_n700), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT35), .B(G1991), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(G16), .A2(G24), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n589), .B2(G16), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT89), .ZN(new_n712));
  INV_X1    g287(.A(G1986), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n698), .A2(new_n699), .A3(new_n709), .A4(new_n714), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n696), .A2(new_n697), .A3(new_n709), .A4(new_n714), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(KEYINPUT36), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n700), .A2(G35), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n700), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT29), .B(G2090), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n605), .A2(G16), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G4), .B2(G16), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT91), .B(G1348), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n486), .A2(G139), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT92), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n618), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(new_n463), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT25), .Z(new_n734));
  NAND3_X1  g309(.A1(new_n730), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  MUX2_X1   g310(.A(G33), .B(new_n735), .S(G29), .Z(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(G2072), .Z(new_n737));
  NAND3_X1  g312(.A1(new_n680), .A2(KEYINPUT23), .A3(G20), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT23), .ZN(new_n739));
  INV_X1    g314(.A(G20), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(G16), .ZN(new_n741));
  INV_X1    g316(.A(G299), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n738), .B(new_n741), .C1(new_n742), .C2(new_n680), .ZN(new_n743));
  INV_X1    g318(.A(G1956), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n724), .A2(new_n726), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n486), .A2(G141), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT26), .Z(new_n749));
  INV_X1    g324(.A(G105), .ZN(new_n750));
  INV_X1    g325(.A(G129), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n749), .B1(new_n465), .B2(new_n750), .C1(new_n490), .C2(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n747), .A2(new_n752), .ZN(new_n753));
  MUX2_X1   g328(.A(G32), .B(new_n753), .S(G29), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT93), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT27), .B(G1996), .Z(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n737), .A2(new_n745), .A3(new_n746), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n628), .A2(G29), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT30), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(G28), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(G28), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n761), .A2(new_n762), .A3(new_n700), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  AND2_X1   g339(.A1(KEYINPUT24), .A2(G34), .ZN(new_n765));
  NOR2_X1   g340(.A1(KEYINPUT24), .A2(G34), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n765), .A2(new_n766), .A3(G29), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n482), .B2(G29), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n759), .B(new_n763), .C1(new_n764), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n764), .ZN(new_n770));
  NOR2_X1   g345(.A1(G171), .A2(new_n680), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G5), .B2(new_n680), .ZN(new_n772));
  INV_X1    g347(.A(G1961), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AOI211_X1 g349(.A(new_n769), .B(new_n774), .C1(new_n773), .C2(new_n772), .ZN(new_n775));
  NOR2_X1   g350(.A1(G27), .A2(G29), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G164), .B2(G29), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n755), .A2(new_n756), .B1(G2078), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n556), .A2(G16), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G16), .B2(G19), .ZN(new_n780));
  INV_X1    g355(.A(G1341), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT31), .B(G11), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n775), .A2(new_n778), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n777), .A2(G2078), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n486), .A2(G140), .ZN(new_n786));
  INV_X1    g361(.A(G128), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n463), .A2(G116), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n490), .A2(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(new_n700), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n700), .A2(G26), .ZN(new_n793));
  OAI21_X1  g368(.A(KEYINPUT28), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(KEYINPUT28), .B2(new_n793), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n785), .B1(new_n795), .B2(G2067), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G2067), .B2(new_n795), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n780), .A2(new_n781), .ZN(new_n798));
  NOR4_X1   g373(.A1(new_n758), .A2(new_n784), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n718), .A2(new_n722), .A3(new_n727), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(G168), .A2(G16), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G16), .B2(G21), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT94), .B(G1966), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n800), .A2(new_n804), .ZN(G311));
  INV_X1    g380(.A(new_n799), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n717), .B2(new_n715), .ZN(new_n807));
  INV_X1    g382(.A(new_n804), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n807), .A2(new_n808), .A3(new_n722), .A4(new_n727), .ZN(G150));
  NAND2_X1  g384(.A1(new_n605), .A2(G559), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT38), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n513), .A2(G67), .ZN(new_n812));
  NAND2_X1  g387(.A1(G80), .A2(G543), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n506), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n523), .B2(G55), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n516), .A2(G93), .A3(new_n517), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n815), .A2(new_n816), .A3(KEYINPUT95), .ZN(new_n817));
  AOI21_X1  g392(.A(KEYINPUT95), .B1(new_n815), .B2(new_n816), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n555), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n815), .A2(new_n816), .ZN(new_n820));
  OAI21_X1  g395(.A(KEYINPUT96), .B1(new_n820), .B2(new_n555), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g397(.A(KEYINPUT96), .B(new_n555), .C1(new_n817), .C2(new_n818), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT39), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n811), .B(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT97), .Z(new_n828));
  NOR2_X1   g403(.A1(new_n817), .A2(new_n818), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n828), .A2(new_n831), .ZN(G145));
  NAND2_X1  g407(.A1(new_n486), .A2(G142), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT98), .Z(new_n834));
  OR2_X1    g409(.A1(G106), .A2(G2105), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n835), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n836));
  INV_X1    g411(.A(G130), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n490), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n628), .B(new_n482), .ZN(new_n841));
  INV_X1    g416(.A(G162), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n842), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n840), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n845), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n839), .B1(new_n847), .B2(new_n843), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n620), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n735), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n791), .B(G164), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n730), .A2(new_n620), .A3(new_n732), .A4(new_n734), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n852), .B1(new_n851), .B2(new_n853), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n849), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n854), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n846), .B(new_n848), .C1(new_n858), .C2(new_n855), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n753), .B(new_n706), .Z(new_n860));
  AND3_X1   g435(.A1(new_n857), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n860), .B1(new_n857), .B2(new_n859), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g441(.A1(new_n829), .A2(new_n608), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n614), .B(new_n824), .Z(new_n868));
  INV_X1    g443(.A(new_n603), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT10), .B1(new_n593), .B2(new_n595), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n871), .A2(new_n872), .A3(G299), .A4(new_n602), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n598), .A2(G299), .A3(new_n602), .A4(new_n603), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT99), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT100), .B1(new_n604), .B2(new_n742), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n604), .A2(KEYINPUT100), .A3(new_n742), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n868), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(KEYINPUT101), .Z(new_n882));
  AND4_X1   g457(.A1(KEYINPUT41), .A2(new_n876), .A3(new_n878), .A4(new_n879), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n604), .A2(KEYINPUT100), .A3(new_n742), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n884), .A2(new_n877), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT41), .B1(new_n885), .B2(new_n876), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n882), .B1(new_n887), .B2(new_n868), .ZN(new_n888));
  XNOR2_X1  g463(.A(G303), .B(G288), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(G305), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(G290), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT42), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n888), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n867), .B1(new_n893), .B2(new_n608), .ZN(G295));
  OAI21_X1  g469(.A(new_n867), .B1(new_n893), .B2(new_n608), .ZN(G331));
  NAND2_X1  g470(.A1(G286), .A2(G171), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n529), .A2(new_n531), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT75), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n532), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n900), .A2(G301), .A3(new_n527), .A4(new_n528), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n824), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n883), .B2(new_n886), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n906), .B2(new_n903), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n902), .A2(new_n824), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n896), .A2(new_n901), .B1(new_n822), .B2(new_n823), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(KEYINPUT103), .A3(new_n880), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n904), .A2(new_n891), .A3(new_n907), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n864), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n910), .A2(KEYINPUT103), .A3(new_n880), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT103), .B1(new_n910), .B2(new_n880), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n891), .B1(new_n916), .B2(new_n904), .ZN(new_n917));
  XNOR2_X1  g492(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n918));
  OR3_X1    g493(.A1(new_n913), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT104), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  INV_X1    g496(.A(new_n913), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n904), .B1(new_n906), .B2(new_n903), .ZN(new_n923));
  INV_X1    g498(.A(new_n891), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n921), .B1(new_n926), .B2(KEYINPUT43), .ZN(new_n927));
  OR4_X1    g502(.A1(KEYINPUT104), .A2(new_n913), .A3(new_n917), .A4(new_n918), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n920), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n918), .B1(new_n913), .B2(new_n917), .ZN(new_n930));
  INV_X1    g505(.A(new_n918), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n925), .A2(new_n864), .A3(new_n931), .A4(new_n912), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n921), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n934), .ZN(G397));
  INV_X1    g510(.A(G1384), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n497), .B2(new_n501), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n467), .A2(G40), .A3(new_n474), .A4(new_n481), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n939), .A2(G2067), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(KEYINPUT50), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n941), .B(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n944), .B(new_n936), .C1(new_n497), .C2(new_n501), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n945), .A2(KEYINPUT109), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(KEYINPUT109), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n938), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n940), .B1(new_n949), .B2(new_n726), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT60), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT60), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n725), .B1(new_n943), .B2(new_n948), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n952), .B1(new_n953), .B2(new_n940), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n605), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n950), .A2(KEYINPUT60), .A3(new_n604), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n937), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n938), .ZN(new_n960));
  OAI211_X1 g535(.A(KEYINPUT45), .B(new_n936), .C1(new_n497), .C2(new_n501), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  XOR2_X1   g538(.A(KEYINPUT121), .B(G1996), .Z(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT58), .B(G1341), .Z(new_n966));
  NAND2_X1  g541(.A1(new_n939), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n555), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n968), .B(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT61), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT116), .B1(new_n941), .B2(new_n960), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT116), .ZN(new_n973));
  AOI211_X1 g548(.A(new_n973), .B(new_n938), .C1(new_n937), .C2(KEYINPUT50), .ZN(new_n974));
  INV_X1    g549(.A(new_n945), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(KEYINPUT56), .B(G2072), .Z(new_n977));
  OAI22_X1  g552(.A1(new_n976), .A2(G1956), .B1(new_n962), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT57), .ZN(new_n979));
  NAND2_X1  g554(.A1(G299), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n564), .A2(KEYINPUT57), .A3(new_n567), .A4(new_n574), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT118), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT118), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n980), .A2(new_n984), .A3(new_n981), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT119), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n978), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n962), .A2(new_n977), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n941), .A2(new_n960), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n973), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n941), .A2(KEYINPUT116), .A3(new_n960), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n945), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n990), .B1(new_n994), .B2(new_n744), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT119), .B1(new_n995), .B2(new_n986), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n989), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n982), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n971), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n971), .ZN(new_n1000));
  INV_X1    g575(.A(new_n982), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n1001), .B2(new_n978), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n957), .B(new_n970), .C1(new_n999), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n950), .B2(new_n604), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT117), .B(new_n605), .C1(new_n953), .C2(new_n940), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n988), .B1(new_n978), .B2(new_n987), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n995), .A2(KEYINPUT119), .A3(new_n986), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1005), .B(new_n1006), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n998), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT120), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1009), .A2(KEYINPUT120), .A3(new_n998), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1003), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G303), .A2(G8), .ZN(new_n1015));
  NAND2_X1  g590(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g592(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n949), .A2(G2090), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT108), .B(G1971), .Z(new_n1021));
  NAND2_X1  g596(.A1(new_n962), .A2(KEYINPUT107), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT107), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n959), .A2(new_n1023), .A3(new_n960), .A4(new_n961), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1021), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(G8), .B(new_n1019), .C1(new_n1020), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1021), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(G2090), .B2(new_n949), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1032), .A2(KEYINPUT112), .A3(G8), .A4(new_n1019), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1028), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n939), .A2(G8), .ZN(new_n1035));
  INV_X1    g610(.A(G1976), .ZN(new_n1036));
  NOR2_X1   g611(.A1(G288), .A2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1035), .A2(KEYINPUT114), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT113), .B(G1976), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G288), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1039), .B1(new_n1035), .B2(new_n1041), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1044));
  XNOR2_X1  g619(.A(G305), .B(G1981), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1045), .B(KEYINPUT49), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1035), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1043), .A2(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n994), .A2(G2090), .ZN(new_n1049));
  OAI21_X1  g624(.A(G8), .B1(new_n1049), .B2(new_n1025), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1019), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1034), .A2(new_n1048), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G2078), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1022), .A2(new_n1054), .A3(new_n1024), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT124), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1057), .B(new_n1058), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n962), .A2(new_n1056), .A3(G2078), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n949), .B2(new_n773), .ZN(new_n1061));
  AOI21_X1  g636(.A(G301), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT124), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1064));
  OAI211_X1 g639(.A(G301), .B(new_n1061), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT54), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G171), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(new_n1065), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1053), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n943), .A2(new_n948), .A3(new_n764), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n963), .A2(G1966), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G8), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(G286), .A2(G8), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1076), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1083));
  OAI211_X1 g658(.A(G8), .B(new_n1079), .C1(new_n1075), .C2(G286), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1076), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G286), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1014), .A2(new_n1072), .A3(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1048), .B(new_n1086), .C1(new_n1019), .C2(new_n1032), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT63), .B1(new_n1090), .B2(G286), .ZN(new_n1091));
  AOI211_X1 g666(.A(G1976), .B(G288), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1092));
  NOR2_X1   g667(.A1(G305), .A2(G1981), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1093), .B(KEYINPUT115), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1047), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT63), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1052), .A2(new_n1097), .A3(G168), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1034), .B1(new_n1098), .B2(new_n1076), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1096), .B1(new_n1048), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1085), .A2(new_n1101), .A3(new_n1087), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1028), .A2(new_n1033), .B1(new_n1051), .B2(new_n1050), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1102), .A2(new_n1103), .A3(new_n1048), .A4(new_n1062), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1101), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT125), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1102), .A2(new_n1062), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1053), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1105), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1089), .A2(new_n1100), .A3(new_n1106), .A4(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n959), .A2(new_n938), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n589), .A2(new_n713), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1114), .B(KEYINPUT105), .Z(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n713), .B2(new_n589), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n706), .B(new_n708), .ZN(new_n1118));
  XOR2_X1   g693(.A(new_n1118), .B(KEYINPUT106), .Z(new_n1119));
  XNOR2_X1  g694(.A(new_n791), .B(G2067), .ZN(new_n1120));
  INV_X1    g695(.A(G1996), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n753), .B(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1113), .B1(new_n1117), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1112), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1120), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1113), .B1(new_n1126), .B2(new_n753), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1113), .A2(new_n1121), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT46), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT47), .ZN(new_n1131));
  AND4_X1   g706(.A1(new_n708), .A2(new_n1122), .A3(new_n706), .A4(new_n1120), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n786), .A2(G2067), .A3(new_n790), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1113), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1123), .A2(new_n1113), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT126), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1115), .A2(new_n1113), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT48), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1135), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1125), .A2(new_n1140), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g716(.A1(G401), .A2(G227), .ZN(new_n1143));
  AOI21_X1  g717(.A(new_n1143), .B1(new_n863), .B2(new_n864), .ZN(new_n1144));
  NAND4_X1  g718(.A1(new_n933), .A2(new_n461), .A3(new_n678), .A4(new_n1144), .ZN(G225));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n1146));
  NAND2_X1  g720(.A1(G225), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g721(.A(new_n461), .ZN(new_n1148));
  AOI21_X1  g722(.A(new_n1148), .B1(new_n930), .B2(new_n932), .ZN(new_n1149));
  NAND4_X1  g723(.A1(new_n1149), .A2(KEYINPUT127), .A3(new_n678), .A4(new_n1144), .ZN(new_n1150));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1150), .ZN(G308));
endmodule


