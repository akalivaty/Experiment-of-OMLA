//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n469), .B(KEYINPUT64), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n463), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n467), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n472), .A2(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n463), .A2(new_n468), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  OAI211_X1 g057(.A(G138), .B(new_n468), .C1(new_n461), .C2(new_n462), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  OR2_X1    g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n477), .A2(G126), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n484), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n485), .A2(new_n486), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G164));
  XNOR2_X1  g066(.A(KEYINPUT5), .B(G543), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G62), .ZN(new_n493));
  NAND2_X1  g068(.A1(G75), .A2(G543), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(KEYINPUT65), .B1(new_n495), .B2(G651), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT6), .B(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G50), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G88), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n498), .A2(new_n499), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n496), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n495), .A2(KEYINPUT65), .A3(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(G303));
  INV_X1    g084(.A(G303), .ZN(G166));
  INV_X1    g085(.A(new_n504), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G89), .ZN(new_n512));
  AND3_X1   g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  XOR2_X1   g088(.A(KEYINPUT67), .B(G51), .Z(new_n514));
  OAI221_X1 g089(.A(new_n512), .B1(KEYINPUT7), .B2(new_n513), .C1(new_n498), .C2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(KEYINPUT66), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n520), .B1(new_n501), .B2(new_n500), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G63), .ZN(new_n523));
  NAND3_X1  g098(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n516), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n515), .A2(new_n525), .ZN(G168));
  INV_X1    g101(.A(KEYINPUT69), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n492), .A2(new_n497), .A3(G90), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n529));
  OAI211_X1 g104(.A(G52), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n529), .B1(new_n528), .B2(new_n530), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n519), .A2(new_n521), .A3(G64), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n516), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n527), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n528), .A2(new_n530), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT68), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n536), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT69), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n537), .A2(new_n543), .ZN(G171));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT70), .B(G81), .Z(new_n546));
  OAI22_X1  g121(.A1(new_n498), .A2(new_n545), .B1(new_n504), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT71), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n519), .A2(new_n521), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G651), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g131(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n557));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND3_X1  g135(.A1(new_n497), .A2(G53), .A3(G543), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n504), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n492), .A2(new_n497), .A3(KEYINPUT73), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(G91), .A3(new_n565), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n492), .A2(G65), .ZN(new_n567));
  AND2_X1   g142(.A1(G78), .A2(G543), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND3_X1   g144(.A1(new_n562), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G299));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n537), .A2(new_n572), .A3(new_n543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n572), .B1(new_n537), .B2(new_n543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(G301));
  INV_X1    g150(.A(G168), .ZN(G286));
  AND2_X1   g151(.A1(new_n564), .A2(new_n565), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G87), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n578), .B(new_n579), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n522), .A2(G74), .ZN(new_n581));
  INV_X1    g156(.A(new_n498), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n581), .A2(G651), .B1(G49), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n580), .A2(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(new_n577), .A2(G86), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n492), .A2(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n516), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(G48), .B2(new_n582), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(G72), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G60), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n550), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n516), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI211_X1 g170(.A(KEYINPUT76), .B(new_n591), .C1(new_n550), .C2(new_n592), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n595), .A2(KEYINPUT77), .A3(new_n596), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n498), .A2(new_n602), .B1(new_n504), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT78), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n492), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G54), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n610), .A2(new_n516), .B1(new_n611), .B2(new_n498), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n564), .A2(G92), .A3(new_n565), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  AOI21_X1  g194(.A(KEYINPUT78), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n609), .B1(new_n607), .B2(new_n620), .ZN(G284));
  AOI21_X1  g196(.A(new_n609), .B1(new_n607), .B2(new_n620), .ZN(G321));
  NAND2_X1  g197(.A1(G299), .A2(new_n619), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G168), .B2(new_n619), .ZN(G280));
  XNOR2_X1  g199(.A(G280), .B(KEYINPUT80), .ZN(G297));
  INV_X1    g200(.A(new_n618), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g207(.A(new_n463), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n470), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT12), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G2100), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT81), .ZN(new_n638));
  AOI22_X1  g213(.A1(G123), .A2(new_n477), .B1(new_n472), .B2(G135), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n640));
  NOR3_X1   g215(.A1(new_n640), .A2(new_n468), .A3(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n468), .B2(G111), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n642), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n639), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  OAI211_X1 g220(.A(new_n638), .B(new_n645), .C1(G2100), .C2(new_n636), .ZN(G156));
  INV_X1    g221(.A(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(new_n650), .B2(new_n649), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n652), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n659), .A2(G14), .A3(new_n660), .ZN(G401));
  INV_X1    g236(.A(KEYINPUT18), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(KEYINPUT17), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2100), .ZN(new_n669));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n665), .B2(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2096), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n675), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n675), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1981), .B(G1986), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT83), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(G229));
  AOI21_X1  g266(.A(new_n604), .B1(new_n599), .B2(new_n600), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G16), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G16), .B2(G24), .ZN(new_n694));
  INV_X1    g269(.A(G1986), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT84), .B(G29), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n699), .A2(G25), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n472), .A2(G131), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n477), .A2(G119), .ZN(new_n702));
  OR2_X1    g277(.A1(G95), .A2(G2105), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n703), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n700), .B1(new_n706), .B2(new_n699), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT35), .B(G1991), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n696), .A2(new_n697), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G23), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n580), .A2(new_n583), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT33), .B(G1976), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n712), .A2(G22), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G166), .B2(new_n712), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1971), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n712), .A2(G6), .ZN(new_n721));
  INV_X1    g296(.A(G305), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n712), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT32), .B(G1981), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  AND3_X1   g301(.A1(new_n717), .A2(KEYINPUT34), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(KEYINPUT34), .B1(new_n717), .B2(new_n726), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n711), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(KEYINPUT36), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(KEYINPUT36), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(G32), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n472), .A2(G141), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G129), .B2(new_n477), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n470), .A2(G105), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT90), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n734), .B1(new_n743), .B2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT92), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT27), .B(G1996), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n712), .A2(G20), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT97), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT23), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G299), .B2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1956), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT94), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n712), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n712), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G1966), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n747), .B(new_n752), .C1(new_n753), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n733), .A2(G33), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n633), .A2(G127), .ZN(new_n759));
  NAND2_X1  g334(.A1(G115), .A2(G2104), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(G2105), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT25), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n472), .A2(G139), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n758), .B1(new_n769), .B2(new_n733), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G2072), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT89), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT24), .B(G34), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n698), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT88), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n474), .B2(new_n733), .ZN(new_n777));
  INV_X1    g352(.A(G2084), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n773), .B(new_n779), .C1(G2072), .C2(new_n770), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n745), .A2(new_n746), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT93), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n757), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(KEYINPUT93), .B1(new_n780), .B2(new_n781), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n698), .A2(G27), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT95), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G164), .B2(new_n698), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT96), .B(G2078), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT30), .B(G28), .ZN(new_n791));
  OR2_X1    g366(.A1(KEYINPUT31), .A2(G11), .ZN(new_n792));
  NAND2_X1  g367(.A1(KEYINPUT31), .A2(G11), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n791), .A2(new_n733), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n644), .B2(new_n698), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n778), .B2(new_n777), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n788), .A2(new_n789), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI211_X1 g373(.A(new_n790), .B(new_n798), .C1(new_n753), .C2(new_n756), .ZN(new_n799));
  NAND2_X1  g374(.A1(G162), .A2(new_n699), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n699), .A2(G35), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT29), .ZN(new_n803));
  INV_X1    g378(.A(G2090), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n712), .A2(G19), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n554), .B2(new_n712), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n803), .A2(new_n804), .B1(G1341), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n472), .A2(G140), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n477), .A2(G128), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n468), .A2(G116), .ZN(new_n810));
  OAI21_X1  g385(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n808), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G29), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT86), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n698), .A2(G26), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT87), .Z(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT28), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(G2067), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n803), .A2(new_n804), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n799), .A2(new_n807), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n806), .A2(G1341), .B1(G1966), .B2(new_n755), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G2067), .B2(new_n818), .ZN(new_n823));
  NOR2_X1   g398(.A1(G4), .A2(G16), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT85), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n618), .B2(new_n712), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1348), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(G5), .A2(G16), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G171), .B2(G16), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G1961), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n784), .A2(new_n785), .A3(new_n829), .A4(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(KEYINPUT98), .B1(new_n732), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n837));
  AOI211_X1 g412(.A(new_n837), .B(new_n834), .C1(new_n730), .C2(new_n731), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n836), .A2(new_n838), .ZN(G311));
  NAND2_X1  g414(.A1(new_n732), .A2(new_n835), .ZN(G150));
  NAND2_X1  g415(.A1(new_n522), .A2(G67), .ZN(new_n841));
  NAND2_X1  g416(.A1(G80), .A2(G543), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n516), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(G55), .ZN(new_n844));
  INV_X1    g419(.A(G93), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n498), .A2(new_n844), .B1(new_n504), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n847), .A2(new_n553), .A3(new_n548), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n548), .A2(new_n553), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n841), .A2(new_n842), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G651), .ZN(new_n851));
  INV_X1    g426(.A(new_n846), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n851), .A2(KEYINPUT99), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n843), .B2(new_n846), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n848), .B1(new_n849), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT38), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n627), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n861));
  AOI21_X1  g436(.A(G860), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n861), .B2(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n856), .A2(G860), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT37), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(G145));
  XNOR2_X1  g441(.A(new_n474), .B(new_n481), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n644), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n812), .B(new_n490), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n743), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n769), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n477), .A2(G130), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n468), .A2(G118), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(G142), .B2(new_n472), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n635), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n706), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT100), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n871), .A2(new_n878), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT101), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n868), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n882), .A2(new_n868), .ZN(new_n885));
  AOI21_X1  g460(.A(G37), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n884), .A2(KEYINPUT40), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT40), .B1(new_n884), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(G395));
  NAND2_X1  g464(.A1(new_n856), .A2(new_n619), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n692), .A2(KEYINPUT104), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n692), .A2(KEYINPUT104), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n714), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n895));
  NAND2_X1  g470(.A1(G290), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n692), .A2(KEYINPUT104), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(G288), .A3(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G303), .B(G305), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n893), .A2(new_n894), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n891), .A2(new_n892), .A3(new_n714), .ZN(new_n901));
  AOI21_X1  g476(.A(G288), .B1(new_n896), .B2(new_n897), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n899), .B(new_n894), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n629), .B(KEYINPUT102), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT99), .B1(new_n851), .B2(new_n852), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n843), .A2(new_n854), .A3(new_n846), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n849), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n554), .A2(new_n847), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n908), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n618), .A2(G299), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n614), .A2(new_n570), .A3(new_n617), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n614), .A2(new_n570), .A3(new_n617), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n570), .B1(new_n614), .B2(new_n617), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g496(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n922));
  OAI21_X1  g497(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n914), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n914), .B2(new_n921), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n907), .B(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n890), .B1(new_n927), .B2(new_n619), .ZN(G295));
  OAI21_X1  g503(.A(new_n890), .B1(new_n927), .B2(new_n619), .ZN(G331));
  XNOR2_X1  g504(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n915), .A2(new_n917), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n931), .A2(new_n922), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(new_n916), .B2(new_n931), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n533), .A2(new_n527), .A3(new_n536), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT69), .B1(new_n541), .B2(new_n542), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT74), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n537), .A2(new_n572), .A3(new_n543), .ZN(new_n937));
  AOI21_X1  g512(.A(G286), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(G171), .A2(G168), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n857), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(G168), .B1(new_n573), .B2(new_n574), .ZN(new_n941));
  INV_X1    g516(.A(new_n939), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n913), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n933), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n931), .B1(new_n940), .B2(new_n943), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n933), .A2(new_n940), .A3(new_n943), .A4(KEYINPUT111), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n905), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n940), .A2(new_n943), .A3(new_n923), .A4(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n940), .A2(new_n943), .A3(new_n923), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT109), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n953), .B1(new_n955), .B2(new_n947), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n899), .A2(new_n894), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n901), .A2(new_n902), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n904), .B1(new_n893), .B2(new_n898), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(G37), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n951), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n905), .B(new_n953), .C1(new_n947), .C2(new_n955), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n962), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n963), .B1(new_n965), .B2(KEYINPUT110), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n967));
  AOI211_X1 g542(.A(new_n967), .B(new_n962), .C1(new_n961), .C2(new_n964), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n930), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n961), .A2(new_n964), .A3(new_n962), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n951), .A2(new_n961), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT44), .B(new_n970), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(G397));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n490), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT45), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n977), .B2(new_n976), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n467), .A2(new_n471), .A3(G40), .A4(new_n473), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n706), .A2(new_n708), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n705), .A2(new_n709), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n812), .B(G2067), .Z(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1996), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n743), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n740), .A2(new_n742), .A3(G1996), .ZN(new_n989));
  AOI211_X1 g564(.A(new_n984), .B(new_n986), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n695), .B2(new_n692), .ZN(new_n991));
  NOR2_X1   g566(.A1(G290), .A2(G1986), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n981), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT125), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT118), .B(G86), .Z(new_n995));
  NAND2_X1  g570(.A1(new_n511), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n589), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(G1981), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT117), .B(G1981), .Z(new_n999));
  NAND3_X1  g574(.A1(new_n585), .A2(new_n589), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT119), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT49), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(KEYINPUT119), .A3(KEYINPUT49), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n976), .A2(KEYINPUT113), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n490), .A2(new_n1008), .A3(new_n975), .ZN(new_n1009));
  INV_X1    g584(.A(new_n980), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G8), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(KEYINPUT116), .A3(G8), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1006), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n714), .A2(G1976), .ZN(new_n1018));
  INV_X1    g593(.A(G1976), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(G288), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1015), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT116), .B1(new_n1011), .B2(G8), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1018), .B(new_n1020), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1017), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1010), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n804), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1971), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n976), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1010), .B1(new_n976), .B2(new_n1032), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1025), .B1(new_n1030), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G303), .A2(G8), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1037), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1024), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n490), .A2(new_n975), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n980), .B1(new_n1050), .B2(KEYINPUT45), .ZN(new_n1051));
  INV_X1    g626(.A(G2078), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(new_n1052), .A3(new_n1033), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1007), .A2(new_n1054), .A3(new_n1009), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n980), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1961), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1049), .A2(new_n1053), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n979), .A2(KEYINPUT53), .A3(new_n1052), .A4(new_n1051), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(G301), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT45), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(new_n1035), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1064), .A2(KEYINPUT53), .A3(new_n1052), .ZN(new_n1065));
  AOI21_X1  g640(.A(G301), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1048), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1036), .B1(new_n1057), .B2(G2090), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1068), .A2(new_n1043), .A3(G8), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT115), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1068), .A2(new_n1043), .A3(new_n1071), .A4(G8), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1053), .A2(new_n1049), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1057), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1074), .B(new_n1060), .C1(new_n1075), .C2(G1961), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1048), .B1(new_n1076), .B2(G171), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1059), .A2(G301), .A3(new_n1065), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1047), .A2(new_n1067), .A3(new_n1073), .A4(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT120), .B1(new_n1057), .B2(G2084), .ZN(new_n1081));
  INV_X1    g656(.A(G1966), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n1063), .B2(new_n1035), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1055), .A2(new_n1084), .A3(new_n778), .A4(new_n1056), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1081), .A2(G168), .A3(new_n1083), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G8), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1087), .A2(KEYINPUT51), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1081), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G286), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(G8), .A3(new_n1086), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1088), .B1(new_n1092), .B2(KEYINPUT51), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n994), .B1(new_n1080), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1028), .B1(new_n1026), .B2(KEYINPUT50), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT121), .B(G1956), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT56), .B(G2072), .Z(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n570), .B(KEYINPUT57), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1098), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n618), .ZN(new_n1105));
  OAI22_X1  g680(.A1(new_n1075), .A2(G1348), .B1(G2067), .B2(new_n1011), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1011), .A2(G2067), .ZN(new_n1109));
  INV_X1    g684(.A(G1348), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(new_n1057), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(KEYINPUT122), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1098), .A2(KEYINPUT123), .A3(new_n1102), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1102), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1103), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1105), .A2(new_n1113), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1114), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1115), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1121), .B2(new_n1103), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(KEYINPUT60), .B(new_n618), .C1(new_n1108), .C2(new_n1112), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1103), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1120), .B1(new_n1104), .B2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT58), .B(G1341), .Z(new_n1127));
  AOI22_X1  g702(.A1(new_n1099), .A2(new_n987), .B1(new_n1011), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(new_n849), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT59), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1129), .B(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .A4(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1108), .A2(new_n1112), .A3(KEYINPUT60), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1111), .A2(KEYINPUT122), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1134), .A2(new_n1138), .A3(new_n618), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1118), .B1(new_n1133), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1046), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1037), .A2(new_n1043), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1141), .A2(new_n1142), .A3(new_n1023), .A4(new_n1017), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1073), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1066), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1061), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1147), .A2(new_n1048), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1148));
  AOI21_X1  g723(.A(G168), .B1(new_n1089), .B2(new_n1081), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT51), .B1(new_n1087), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(KEYINPUT51), .B2(new_n1087), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1145), .A2(new_n1148), .A3(new_n1151), .A4(KEYINPUT125), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1094), .A2(new_n1140), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1090), .A2(G8), .ZN(new_n1154));
  NOR2_X1   g729(.A1(G286), .A2(KEYINPUT63), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1037), .B2(new_n1043), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1073), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1024), .A2(new_n1046), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1141), .A2(new_n1023), .A3(new_n1017), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1068), .A2(G8), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1043), .ZN(new_n1162));
  AOI21_X1  g737(.A(G286), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1163), .A2(G8), .A3(new_n1090), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT63), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1165));
  AOI211_X1 g740(.A(G1976), .B(G288), .C1(new_n1006), .C2(new_n1016), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1000), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1016), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1159), .A2(new_n1165), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1145), .B(new_n1066), .C1(new_n1093), .C2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1151), .A2(KEYINPUT62), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1169), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n993), .B1(new_n1153), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n981), .B1(new_n743), .B2(new_n986), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n981), .A2(new_n987), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1176), .A2(KEYINPUT46), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1176), .A2(KEYINPUT46), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1175), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT47), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n990), .A2(new_n980), .A3(new_n979), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n992), .A2(new_n981), .ZN(new_n1182));
  XNOR2_X1  g757(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1184), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1185));
  AOI211_X1 g760(.A(new_n982), .B(new_n986), .C1(new_n988), .C2(new_n989), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n812), .A2(G2067), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n981), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1180), .A2(new_n1185), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1174), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g765(.A1(new_n966), .A2(new_n968), .ZN(new_n1192));
  NOR4_X1   g766(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1193));
  INV_X1    g767(.A(new_n868), .ZN(new_n1194));
  INV_X1    g768(.A(new_n883), .ZN(new_n1195));
  AOI21_X1  g769(.A(new_n1194), .B1(new_n1195), .B2(new_n880), .ZN(new_n1196));
  INV_X1    g770(.A(new_n886), .ZN(new_n1197));
  OAI21_X1  g771(.A(new_n1193), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g772(.A1(new_n1192), .A2(new_n1198), .ZN(G308));
  OAI221_X1 g773(.A(new_n1193), .B1(new_n1196), .B2(new_n1197), .C1(new_n966), .C2(new_n968), .ZN(G225));
endmodule


