

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U322 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X2 U323 ( .A(n341), .B(n349), .Z(n385) );
  XNOR2_X1 U324 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U325 ( .A(KEYINPUT105), .B(KEYINPUT36), .ZN(n387) );
  XNOR2_X1 U326 ( .A(n352), .B(n351), .ZN(n356) );
  XNOR2_X1 U327 ( .A(n558), .B(n387), .ZN(n582) );
  XNOR2_X1 U328 ( .A(n455), .B(n454), .ZN(n456) );
  INV_X1 U329 ( .A(G190GAT), .ZN(n457) );
  XNOR2_X1 U330 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U331 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n291) );
  XNOR2_X1 U333 ( .A(G113GAT), .B(KEYINPUT83), .ZN(n290) );
  XNOR2_X1 U334 ( .A(n291), .B(n290), .ZN(n298) );
  XOR2_X1 U335 ( .A(KEYINPUT85), .B(G190GAT), .Z(n293) );
  XNOR2_X1 U336 ( .A(G43GAT), .B(G99GAT), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U338 ( .A(n294), .B(KEYINPUT82), .Z(n296) );
  XOR2_X1 U339 ( .A(G120GAT), .B(G71GAT), .Z(n340) );
  XNOR2_X1 U340 ( .A(G15GAT), .B(n340), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n309) );
  XOR2_X1 U343 ( .A(G183GAT), .B(G176GAT), .Z(n300) );
  NAND2_X1 U344 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U346 ( .A(n301), .B(KEYINPUT65), .Z(n307) );
  XOR2_X1 U347 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n303) );
  XNOR2_X1 U348 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n401) );
  XOR2_X1 U350 ( .A(G127GAT), .B(KEYINPUT0), .Z(n305) );
  XNOR2_X1 U351 ( .A(G134GAT), .B(KEYINPUT81), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n431) );
  XNOR2_X1 U353 ( .A(n401), .B(n431), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U355 ( .A(n309), .B(n308), .Z(n539) );
  INV_X1 U356 ( .A(n539), .ZN(n529) );
  XOR2_X1 U357 ( .A(G8GAT), .B(G15GAT), .Z(n311) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(G197GAT), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n326) );
  XOR2_X1 U360 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n313) );
  XNOR2_X1 U361 ( .A(KEYINPUT29), .B(KEYINPUT69), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U363 ( .A(G50GAT), .B(G36GAT), .Z(n315) );
  XOR2_X1 U364 ( .A(G141GAT), .B(G22GAT), .Z(n447) );
  XOR2_X1 U365 ( .A(G113GAT), .B(G1GAT), .Z(n424) );
  XNOR2_X1 U366 ( .A(n447), .B(n424), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U368 ( .A(n317), .B(n316), .Z(n319) );
  NAND2_X1 U369 ( .A1(G229GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U371 ( .A(n320), .B(KEYINPUT30), .Z(n324) );
  XOR2_X1 U372 ( .A(G29GAT), .B(G43GAT), .Z(n322) );
  XNOR2_X1 U373 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n348) );
  XNOR2_X1 U375 ( .A(n348), .B(KEYINPUT68), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n509) );
  INV_X1 U378 ( .A(n509), .ZN(n571) );
  XOR2_X1 U379 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n328) );
  NAND2_X1 U380 ( .A1(G230GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U382 ( .A(n329), .B(KEYINPUT73), .Z(n334) );
  XNOR2_X1 U383 ( .A(G106GAT), .B(G78GAT), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n330), .B(G148GAT), .ZN(n438) );
  XOR2_X1 U385 ( .A(G64GAT), .B(G92GAT), .Z(n332) );
  XNOR2_X1 U386 ( .A(G176GAT), .B(G204GAT), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n400) );
  XNOR2_X1 U388 ( .A(n438), .B(n400), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n336) );
  INV_X1 U390 ( .A(KEYINPUT33), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n338) );
  XOR2_X1 U392 ( .A(G57GAT), .B(KEYINPUT13), .Z(n365) );
  XNOR2_X1 U393 ( .A(n365), .B(KEYINPUT31), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U396 ( .A(G99GAT), .B(G85GAT), .ZN(n349) );
  XOR2_X1 U397 ( .A(KEYINPUT41), .B(n385), .Z(n508) );
  NAND2_X1 U398 ( .A1(n571), .A2(n508), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n342), .B(KEYINPUT46), .ZN(n381) );
  XOR2_X1 U400 ( .A(KEYINPUT74), .B(G92GAT), .Z(n344) );
  XNOR2_X1 U401 ( .A(G218GAT), .B(G106GAT), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U403 ( .A(n345), .B(KEYINPUT76), .Z(n347) );
  XOR2_X1 U404 ( .A(G50GAT), .B(G162GAT), .Z(n446) );
  XNOR2_X1 U405 ( .A(G134GAT), .B(n446), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n352) );
  XOR2_X1 U407 ( .A(G36GAT), .B(G190GAT), .Z(n395) );
  XNOR2_X1 U408 ( .A(n348), .B(n395), .ZN(n350) );
  XOR2_X1 U409 ( .A(KEYINPUT64), .B(KEYINPUT10), .Z(n354) );
  NAND2_X1 U410 ( .A1(G232GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U412 ( .A(n356), .B(n355), .Z(n361) );
  XOR2_X1 U413 ( .A(KEYINPUT11), .B(KEYINPUT77), .Z(n358) );
  XNOR2_X1 U414 ( .A(KEYINPUT66), .B(KEYINPUT9), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n359), .B(KEYINPUT75), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n558) );
  XOR2_X1 U418 ( .A(G78GAT), .B(G155GAT), .Z(n363) );
  XNOR2_X1 U419 ( .A(G22GAT), .B(G211GAT), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U421 ( .A(n365), .B(n364), .Z(n367) );
  NAND2_X1 U422 ( .A1(G231GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U424 ( .A(n368), .B(KEYINPUT14), .Z(n371) );
  XNOR2_X1 U425 ( .A(G8GAT), .B(G183GAT), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n369), .B(KEYINPUT78), .ZN(n398) );
  XNOR2_X1 U427 ( .A(n398), .B(KEYINPUT80), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n379) );
  XOR2_X1 U429 ( .A(G71GAT), .B(G127GAT), .Z(n373) );
  XNOR2_X1 U430 ( .A(G15GAT), .B(G1GAT), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U432 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n375) );
  XNOR2_X1 U433 ( .A(G64GAT), .B(KEYINPUT79), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U435 ( .A(n377), .B(n376), .Z(n378) );
  XOR2_X1 U436 ( .A(n379), .B(n378), .Z(n578) );
  NOR2_X1 U437 ( .A1(n558), .A2(n578), .ZN(n380) );
  AND2_X1 U438 ( .A1(n381), .A2(n380), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n382), .B(KEYINPUT115), .ZN(n384) );
  INV_X1 U440 ( .A(KEYINPUT47), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n393) );
  XNOR2_X1 U442 ( .A(KEYINPUT116), .B(KEYINPUT45), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n386), .B(KEYINPUT67), .ZN(n389) );
  INV_X1 U444 ( .A(n578), .ZN(n461) );
  NOR2_X1 U445 ( .A1(n582), .A2(n461), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n390) );
  NOR2_X1 U447 ( .A1(n385), .A2(n390), .ZN(n391) );
  NAND2_X1 U448 ( .A1(n391), .A2(n509), .ZN(n392) );
  NAND2_X1 U449 ( .A1(n393), .A2(n392), .ZN(n394) );
  XNOR2_X1 U450 ( .A(n394), .B(KEYINPUT48), .ZN(n537) );
  XOR2_X1 U451 ( .A(KEYINPUT96), .B(n395), .Z(n397) );
  NAND2_X1 U452 ( .A1(G226GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n399) );
  XOR2_X1 U454 ( .A(n399), .B(n398), .Z(n403) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U456 ( .A(n403), .B(n402), .ZN(n408) );
  XOR2_X1 U457 ( .A(KEYINPUT86), .B(G218GAT), .Z(n405) );
  XNOR2_X1 U458 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U460 ( .A(G197GAT), .B(n406), .ZN(n451) );
  INV_X1 U461 ( .A(n451), .ZN(n407) );
  XOR2_X1 U462 ( .A(n408), .B(n407), .Z(n466) );
  NAND2_X1 U463 ( .A1(n537), .A2(n466), .ZN(n410) );
  XOR2_X1 U464 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n434) );
  XOR2_X1 U466 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n412) );
  XNOR2_X1 U467 ( .A(KEYINPUT95), .B(KEYINPUT94), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U469 ( .A(KEYINPUT1), .B(G57GAT), .Z(n414) );
  XNOR2_X1 U470 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U472 ( .A(n416), .B(n415), .Z(n421) );
  XOR2_X1 U473 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n418) );
  NAND2_X1 U474 ( .A1(G225GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U476 ( .A(KEYINPUT91), .B(n419), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n429) );
  XOR2_X1 U478 ( .A(G85GAT), .B(G162GAT), .Z(n423) );
  XNOR2_X1 U479 ( .A(G120GAT), .B(G148GAT), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U481 ( .A(n425), .B(n424), .Z(n427) );
  XNOR2_X1 U482 ( .A(G29GAT), .B(G141GAT), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U484 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U485 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n430), .B(KEYINPUT2), .ZN(n439) );
  XNOR2_X1 U487 ( .A(n431), .B(n439), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n524) );
  NAND2_X1 U489 ( .A1(n434), .A2(n524), .ZN(n570) );
  XOR2_X1 U490 ( .A(KEYINPUT89), .B(KEYINPUT24), .Z(n436) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U493 ( .A(n437), .B(KEYINPUT23), .Z(n441) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U496 ( .A(G204GAT), .B(KEYINPUT88), .Z(n443) );
  XNOR2_X1 U497 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U499 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U502 ( .A(n451), .B(n450), .Z(n470) );
  NOR2_X1 U503 ( .A1(n570), .A2(n470), .ZN(n455) );
  XNOR2_X1 U504 ( .A(KEYINPUT122), .B(KEYINPUT55), .ZN(n453) );
  INV_X1 U505 ( .A(KEYINPUT121), .ZN(n452) );
  NOR2_X1 U506 ( .A1(n529), .A2(n456), .ZN(n567) );
  NAND2_X1 U507 ( .A1(n567), .A2(n558), .ZN(n460) );
  XOR2_X1 U508 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n458) );
  NOR2_X1 U509 ( .A1(n385), .A2(n509), .ZN(n497) );
  NOR2_X1 U510 ( .A1(n558), .A2(n461), .ZN(n462) );
  XNOR2_X1 U511 ( .A(KEYINPUT16), .B(n462), .ZN(n481) );
  INV_X1 U512 ( .A(n466), .ZN(n527) );
  XNOR2_X1 U513 ( .A(n527), .B(KEYINPUT97), .ZN(n463) );
  XOR2_X1 U514 ( .A(KEYINPUT27), .B(n463), .Z(n474) );
  NOR2_X1 U515 ( .A1(n524), .A2(n474), .ZN(n464) );
  XNOR2_X1 U516 ( .A(KEYINPUT98), .B(n464), .ZN(n536) );
  XOR2_X1 U517 ( .A(KEYINPUT28), .B(n470), .Z(n535) );
  AND2_X1 U518 ( .A1(n536), .A2(n535), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n529), .A2(n465), .ZN(n479) );
  NAND2_X1 U520 ( .A1(n466), .A2(n539), .ZN(n467) );
  XNOR2_X1 U521 ( .A(KEYINPUT101), .B(n467), .ZN(n468) );
  NOR2_X1 U522 ( .A1(n470), .A2(n468), .ZN(n469) );
  XNOR2_X1 U523 ( .A(n469), .B(KEYINPUT25), .ZN(n476) );
  XOR2_X1 U524 ( .A(KEYINPUT100), .B(KEYINPUT26), .Z(n472) );
  NAND2_X1 U525 ( .A1(n529), .A2(n470), .ZN(n471) );
  XNOR2_X1 U526 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U527 ( .A(KEYINPUT99), .B(n473), .ZN(n569) );
  OR2_X1 U528 ( .A1(n569), .A2(n474), .ZN(n475) );
  NAND2_X1 U529 ( .A1(n476), .A2(n475), .ZN(n477) );
  NAND2_X1 U530 ( .A1(n524), .A2(n477), .ZN(n478) );
  NAND2_X1 U531 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U532 ( .A(KEYINPUT102), .B(n480), .ZN(n495) );
  NAND2_X1 U533 ( .A1(n481), .A2(n495), .ZN(n510) );
  INV_X1 U534 ( .A(n510), .ZN(n482) );
  NAND2_X1 U535 ( .A1(n497), .A2(n482), .ZN(n489) );
  NOR2_X1 U536 ( .A1(n524), .A2(n489), .ZN(n483) );
  XOR2_X1 U537 ( .A(n483), .B(KEYINPUT34), .Z(n484) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(n484), .ZN(G1324GAT) );
  NOR2_X1 U539 ( .A1(n527), .A2(n489), .ZN(n485) );
  XOR2_X1 U540 ( .A(G8GAT), .B(n485), .Z(G1325GAT) );
  NOR2_X1 U541 ( .A1(n529), .A2(n489), .ZN(n487) );
  XNOR2_X1 U542 ( .A(KEYINPUT35), .B(KEYINPUT103), .ZN(n486) );
  XNOR2_X1 U543 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U544 ( .A(G15GAT), .B(n488), .Z(G1326GAT) );
  NOR2_X1 U545 ( .A1(n535), .A2(n489), .ZN(n490) );
  XOR2_X1 U546 ( .A(G22GAT), .B(n490), .Z(G1327GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n492) );
  XNOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U550 ( .A(KEYINPUT104), .B(n493), .ZN(n500) );
  NOR2_X1 U551 ( .A1(n578), .A2(n582), .ZN(n494) );
  NAND2_X1 U552 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U553 ( .A(KEYINPUT37), .B(n496), .ZN(n523) );
  NAND2_X1 U554 ( .A1(n497), .A2(n523), .ZN(n498) );
  XNOR2_X1 U555 ( .A(n498), .B(KEYINPUT38), .ZN(n506) );
  NOR2_X1 U556 ( .A1(n524), .A2(n506), .ZN(n499) );
  XNOR2_X1 U557 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NOR2_X1 U558 ( .A1(n506), .A2(n527), .ZN(n501) );
  XOR2_X1 U559 ( .A(G36GAT), .B(n501), .Z(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n503) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(KEYINPUT108), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n503), .B(n502), .ZN(n505) );
  NOR2_X1 U563 ( .A1(n529), .A2(n506), .ZN(n504) );
  XOR2_X1 U564 ( .A(n505), .B(n504), .Z(G1330GAT) );
  NOR2_X1 U565 ( .A1(n506), .A2(n535), .ZN(n507) );
  XOR2_X1 U566 ( .A(G50GAT), .B(n507), .Z(G1331GAT) );
  BUF_X1 U567 ( .A(n508), .Z(n562) );
  NAND2_X1 U568 ( .A1(n562), .A2(n509), .ZN(n521) );
  NOR2_X1 U569 ( .A1(n521), .A2(n510), .ZN(n511) );
  XOR2_X1 U570 ( .A(KEYINPUT110), .B(n511), .Z(n518) );
  NOR2_X1 U571 ( .A1(n524), .A2(n518), .ZN(n514) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(KEYINPUT111), .ZN(n512) );
  XNOR2_X1 U573 ( .A(n512), .B(KEYINPUT42), .ZN(n513) );
  XNOR2_X1 U574 ( .A(n514), .B(n513), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n518), .A2(n527), .ZN(n515) );
  XOR2_X1 U576 ( .A(KEYINPUT112), .B(n515), .Z(n516) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n516), .ZN(G1333GAT) );
  NOR2_X1 U578 ( .A1(n529), .A2(n518), .ZN(n517) );
  XOR2_X1 U579 ( .A(G71GAT), .B(n517), .Z(G1334GAT) );
  NOR2_X1 U580 ( .A1(n518), .A2(n535), .ZN(n520) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U582 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  INV_X1 U583 ( .A(n521), .ZN(n522) );
  NAND2_X1 U584 ( .A1(n523), .A2(n522), .ZN(n532) );
  NOR2_X1 U585 ( .A1(n524), .A2(n532), .ZN(n526) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(KEYINPUT113), .ZN(n525) );
  XNOR2_X1 U587 ( .A(n526), .B(n525), .ZN(G1336GAT) );
  NOR2_X1 U588 ( .A1(n527), .A2(n532), .ZN(n528) );
  XOR2_X1 U589 ( .A(G92GAT), .B(n528), .Z(G1337GAT) );
  NOR2_X1 U590 ( .A1(n529), .A2(n532), .ZN(n530) );
  XOR2_X1 U591 ( .A(KEYINPUT114), .B(n530), .Z(n531) );
  XNOR2_X1 U592 ( .A(G99GAT), .B(n531), .ZN(G1338GAT) );
  NOR2_X1 U593 ( .A1(n535), .A2(n532), .ZN(n533) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(n533), .Z(n534) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  INV_X1 U596 ( .A(n535), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n537), .A2(n536), .ZN(n551) );
  NOR2_X1 U598 ( .A1(n538), .A2(n551), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U600 ( .A(KEYINPUT117), .B(n541), .ZN(n548) );
  NAND2_X1 U601 ( .A1(n571), .A2(n548), .ZN(n542) );
  XNOR2_X1 U602 ( .A(G113GAT), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U604 ( .A1(n548), .A2(n562), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n546) );
  NAND2_X1 U607 ( .A1(n548), .A2(n578), .ZN(n545) );
  XNOR2_X1 U608 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U609 ( .A(G127GAT), .B(n547), .Z(G1342GAT) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U611 ( .A1(n548), .A2(n558), .ZN(n549) );
  XNOR2_X1 U612 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NOR2_X1 U613 ( .A1(n569), .A2(n551), .ZN(n559) );
  NAND2_X1 U614 ( .A1(n571), .A2(n559), .ZN(n552) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n554) );
  NAND2_X1 U617 ( .A1(n559), .A2(n562), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(n556) );
  XOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT52), .Z(n555) );
  XNOR2_X1 U620 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n559), .A2(n578), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n560), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n571), .A2(n567), .ZN(n561) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(n561), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n564) );
  NAND2_X1 U628 ( .A1(n567), .A2(n562), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(n566) );
  XOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT123), .Z(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n578), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT125), .Z(n573) );
  NOR2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n580) );
  NAND2_X1 U636 ( .A1(n580), .A2(n571), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n573), .B(n572), .ZN(n575) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n580), .A2(n385), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n580), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U645 ( .A(n580), .ZN(n581) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(G218GAT), .B(n585), .Z(G1355GAT) );
endmodule

