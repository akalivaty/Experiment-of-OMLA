//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1046, new_n1047;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT71), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n208), .A2(new_n202), .A3(new_n206), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n207), .A2(KEYINPUT71), .A3(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT73), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT66), .B(G190gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(G183gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  NOR4_X1   g024(.A1(new_n219), .A2(new_n222), .A3(new_n223), .A4(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G169gat), .ZN(new_n227));
  INV_X1    g026(.A(G176gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n228), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(KEYINPUT64), .ZN(new_n234));
  OAI211_X1 g033(.A(KEYINPUT25), .B(new_n232), .C1(new_n234), .C2(new_n230), .ZN(new_n235));
  INV_X1    g034(.A(new_n229), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(new_n230), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(KEYINPUT23), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n221), .A2(new_n223), .A3(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  OAI22_X1  g041(.A1(new_n226), .A2(new_n235), .B1(KEYINPUT25), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n231), .A2(new_n244), .A3(KEYINPUT26), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT26), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT68), .B1(new_n233), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n248), .B(new_n236), .C1(new_n234), .C2(KEYINPUT26), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT27), .B(G183gat), .Z(new_n250));
  OAI21_X1  g049(.A(KEYINPUT67), .B1(new_n250), .B2(new_n218), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT28), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(KEYINPUT67), .B(KEYINPUT28), .C1(new_n250), .C2(new_n218), .ZN(new_n254));
  NAND2_X1  g053(.A1(G183gat), .A2(G190gat), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n249), .A2(new_n253), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT29), .B1(new_n243), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G226gat), .A2(G233gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n217), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n258), .B1(new_n243), .B2(new_n256), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n256), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n261), .B1(new_n264), .B2(new_n258), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n216), .B(new_n260), .C1(new_n265), .C2(new_n217), .ZN(new_n266));
  XNOR2_X1  g065(.A(G8gat), .B(G36gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(G64gat), .ZN(new_n268));
  INV_X1    g067(.A(G92gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n215), .B(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n257), .A2(new_n259), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n272), .B1(new_n273), .B2(new_n261), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n266), .A2(new_n270), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT30), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n266), .A2(KEYINPUT30), .A3(new_n270), .A4(new_n274), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n266), .A2(new_n274), .ZN(new_n279));
  INV_X1    g078(.A(new_n270), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n277), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G85gat), .ZN(new_n284));
  INV_X1    g083(.A(G57gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(G1gat), .B(G29gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT0), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n287), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n285), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n292), .A2(G57gat), .A3(new_n288), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n284), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(G57gat), .B1(new_n292), .B2(new_n288), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n289), .A2(new_n285), .A3(new_n290), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(G85gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT78), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT78), .B1(new_n294), .B2(new_n297), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304));
  INV_X1    g103(.A(G155gat), .ZN(new_n305));
  INV_X1    g104(.A(G162gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n304), .B1(new_n307), .B2(KEYINPUT2), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n309));
  INV_X1    g108(.A(G141gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(G148gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n311), .B1(new_n310), .B2(G148gat), .ZN(new_n312));
  INV_X1    g111(.A(G148gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(G141gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(new_n309), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n308), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n307), .A2(new_n304), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n310), .A2(G148gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n319), .B2(KEYINPUT2), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G113gat), .ZN(new_n322));
  INV_X1    g121(.A(G120gat), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT1), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(new_n322), .B2(new_n323), .ZN(new_n325));
  XNOR2_X1  g124(.A(G127gat), .B(G134gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n326), .B(new_n324), .C1(new_n322), .C2(new_n323), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n321), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n316), .A2(new_n320), .A3(new_n328), .A4(new_n329), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT4), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n316), .A2(new_n320), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT3), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n316), .A2(new_n320), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n330), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n336), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT5), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(new_n330), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n334), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n346), .B1(new_n348), .B2(new_n338), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n343), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(new_n331), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n352), .A2(new_n341), .B1(new_n333), .B2(new_n335), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n338), .A2(KEYINPUT5), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n303), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n345), .A2(new_n349), .B1(new_n353), .B2(new_n354), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT79), .B1(new_n359), .B2(new_n302), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n298), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT6), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n359), .A2(new_n362), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT6), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT35), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n262), .A2(new_n330), .ZN(new_n368));
  INV_X1    g167(.A(G227gat), .ZN(new_n369));
  INV_X1    g168(.A(G233gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n243), .A2(new_n331), .A3(new_n256), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n368), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n374), .A2(KEYINPUT34), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(KEYINPUT34), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT69), .B(G71gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(G99gat), .ZN(new_n379));
  XOR2_X1   g178(.A(G15gat), .B(G43gat), .Z(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n372), .B1(new_n368), .B2(new_n373), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n382), .B2(KEYINPUT33), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n243), .A2(new_n331), .A3(new_n256), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n331), .B1(new_n243), .B2(new_n256), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n371), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n386), .A2(KEYINPUT32), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(KEYINPUT32), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT33), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n391), .A3(new_n381), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n377), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n377), .B1(new_n388), .B2(new_n392), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G22gat), .ZN(new_n396));
  INV_X1    g195(.A(G228gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(new_n370), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n342), .B1(new_n215), .B2(KEYINPUT29), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n340), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n215), .B(KEYINPUT72), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n343), .A2(new_n263), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n398), .B(new_n400), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n215), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT29), .B1(new_n210), .B2(new_n212), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n340), .B1(new_n406), .B2(KEYINPUT3), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n398), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n396), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n410), .A2(KEYINPUT76), .ZN(new_n411));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT31), .B(G50gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n404), .A2(new_n396), .A3(new_n409), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  OAI22_X1  g216(.A1(new_n411), .A2(new_n415), .B1(new_n417), .B2(new_n410), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n404), .A2(new_n409), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G22gat), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n420), .A2(KEYINPUT76), .A3(new_n416), .A4(new_n414), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n283), .A2(new_n367), .A3(new_n395), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT80), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT76), .ZN(new_n425));
  INV_X1    g224(.A(new_n398), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n272), .B2(new_n402), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n408), .B1(new_n427), .B2(new_n400), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n425), .B1(new_n428), .B2(new_n396), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n429), .A2(new_n414), .B1(new_n416), .B2(new_n420), .ZN(new_n430));
  INV_X1    g229(.A(new_n421), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n388), .A2(new_n392), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n375), .A2(new_n376), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n377), .A2(new_n388), .A3(new_n392), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT80), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n283), .A4(new_n367), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n424), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT81), .B1(new_n432), .B2(new_n437), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT81), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n395), .A2(new_n443), .A3(new_n422), .ZN(new_n444));
  INV_X1    g243(.A(new_n363), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n366), .B1(new_n445), .B2(new_n365), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT75), .B1(new_n282), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n270), .B1(new_n266), .B2(new_n274), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n276), .B2(new_n275), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT75), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n450), .A2(new_n451), .A3(new_n446), .A4(new_n278), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n442), .A2(new_n444), .A3(new_n448), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT35), .ZN(new_n454));
  INV_X1    g253(.A(new_n353), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT39), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n338), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n353), .A2(new_n337), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT39), .B1(new_n348), .B2(new_n338), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n457), .B(new_n302), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT40), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n282), .A2(new_n361), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT73), .B1(new_n273), .B2(new_n261), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n216), .B1(new_n463), .B2(new_n260), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n273), .A2(new_n261), .A3(new_n272), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT37), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT38), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n266), .A2(new_n468), .A3(new_n274), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n466), .A2(new_n467), .A3(new_n280), .A4(new_n469), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n361), .A2(new_n363), .B1(KEYINPUT6), .B2(new_n365), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n275), .A3(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n469), .A2(new_n280), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n279), .A2(KEYINPUT37), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n462), .B(new_n422), .C1(new_n472), .C2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT70), .B(KEYINPUT36), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n395), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n437), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n432), .B(KEYINPUT77), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n448), .A2(new_n452), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n441), .A2(new_n454), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n487));
  OR2_X1    g286(.A1(G43gat), .A2(G50gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(G43gat), .A2(G50gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT15), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT82), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT82), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n494), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n496));
  INV_X1    g295(.A(G36gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n493), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G29gat), .A2(G36gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT83), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(KEYINPUT83), .A2(G29gat), .A3(G36gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n491), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n488), .A2(KEYINPUT15), .A3(new_n489), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT15), .ZN(new_n509));
  AND2_X1   g308(.A1(G43gat), .A2(G50gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(G43gat), .A2(G50gat), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n492), .ZN(new_n514));
  AND4_X1   g313(.A1(KEYINPUT84), .A2(new_n513), .A3(new_n505), .A4(new_n514), .ZN(new_n515));
  OR2_X1    g314(.A1(G29gat), .A2(G36gat), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n516), .A2(KEYINPUT14), .B1(new_n496), .B2(new_n497), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(new_n504), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT84), .B1(new_n518), .B2(new_n513), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n507), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT16), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(G1gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT87), .ZN(new_n526));
  INV_X1    g325(.A(G8gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n521), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n527), .B1(new_n521), .B2(new_n526), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n525), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n530), .ZN(new_n532));
  AOI21_X1  g331(.A(G1gat), .B1(new_n521), .B2(new_n522), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n533), .A3(new_n528), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT84), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n508), .A2(new_n512), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n514), .A2(new_n503), .A3(new_n502), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n518), .A2(KEYINPUT84), .A3(new_n513), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n506), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n545));
  OAI21_X1  g344(.A(KEYINPUT86), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT86), .ZN(new_n547));
  INV_X1    g346(.A(new_n545), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n520), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n535), .B1(KEYINPUT17), .B2(new_n544), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n538), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n487), .B1(new_n552), .B2(KEYINPUT18), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n537), .B(KEYINPUT13), .Z(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n531), .A2(new_n534), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n544), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n555), .B1(new_n536), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n558), .B1(new_n552), .B2(KEYINPUT18), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n560));
  XOR2_X1   g359(.A(G113gat), .B(G141gat), .Z(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT11), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G169gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G197gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n563), .A2(G197gat), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n560), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n566), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n564), .A3(KEYINPUT12), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT18), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n556), .B1(new_n520), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(new_n546), .B2(new_n549), .ZN(new_n574));
  OAI211_X1 g373(.A(KEYINPUT88), .B(new_n571), .C1(new_n574), .C2(new_n538), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n553), .A2(new_n559), .A3(new_n570), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n567), .A2(new_n569), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n544), .A2(KEYINPUT86), .A3(new_n545), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n547), .B1(new_n520), .B2(new_n548), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n551), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n538), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(KEYINPUT18), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n558), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n552), .A2(KEYINPUT18), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n577), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n576), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n486), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G64gat), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT90), .B1(new_n590), .B2(G57gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT90), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n592), .A2(new_n285), .A3(G64gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(G57gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT91), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT91), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n591), .A2(new_n593), .A3(new_n597), .A4(new_n594), .ZN(new_n598));
  AND2_X1   g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(KEYINPUT9), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n596), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  OR3_X1    g402(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT89), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n285), .A2(G64gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n594), .ZN(new_n606));
  NAND2_X1  g405(.A1(G71gat), .A2(G78gat), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT9), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G71gat), .B(G78gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT89), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n604), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n603), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT93), .ZN(new_n617));
  XOR2_X1   g416(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n601), .B1(new_n595), .B2(KEYINPUT91), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n609), .A2(new_n606), .B1(new_n611), .B2(KEYINPUT89), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n620), .A2(new_n598), .B1(new_n621), .B2(new_n604), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n535), .B1(KEYINPUT21), .B2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n623), .B(G183gat), .Z(new_n624));
  OR2_X1    g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n619), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G127gat), .B(G155gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n204), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n625), .A2(new_n631), .A3(new_n626), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT96), .ZN(new_n636));
  AND2_X1   g435(.A1(G232gat), .A2(G233gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT41), .ZN(new_n638));
  NAND2_X1  g437(.A1(G99gat), .A2(G106gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT8), .ZN(new_n640));
  NAND2_X1  g439(.A1(G85gat), .A2(G92gat), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT7), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n284), .A2(new_n269), .ZN(new_n644));
  NAND3_X1  g443(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n640), .A2(new_n643), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G99gat), .B(G106gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT94), .ZN(new_n650));
  AOI22_X1  g449(.A1(KEYINPUT8), .A2(new_n639), .B1(new_n284), .B2(new_n269), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n651), .A2(new_n647), .A3(new_n643), .A4(new_n645), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n646), .A2(KEYINPUT94), .A3(new_n648), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n638), .B1(new_n544), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n657), .B1(new_n544), .B2(KEYINPUT17), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n656), .B1(new_n550), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G190gat), .B(G218gat), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n636), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n637), .A2(KEYINPUT41), .ZN(new_n663));
  XNOR2_X1  g462(.A(G134gat), .B(G162gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  AOI21_X1  g464(.A(new_n665), .B1(new_n659), .B2(new_n661), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n655), .B1(new_n520), .B2(new_n572), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n667), .B1(new_n546), .B2(new_n549), .ZN(new_n668));
  OAI211_X1 g467(.A(KEYINPUT96), .B(new_n660), .C1(new_n668), .C2(new_n656), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n662), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n659), .A2(new_n661), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n668), .A2(new_n660), .A3(new_n656), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n665), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT95), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n660), .B1(new_n668), .B2(new_n656), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n658), .B1(new_n578), .B2(new_n579), .ZN(new_n676));
  INV_X1    g475(.A(new_n656), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n661), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT95), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n665), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n670), .B1(new_n674), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n635), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(G230gat), .A2(G233gat), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n603), .A2(new_n613), .A3(new_n649), .A4(new_n652), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT10), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n686), .B(new_n687), .C1(new_n657), .C2(new_n622), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n603), .A2(KEYINPUT10), .A3(new_n613), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n657), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n685), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n655), .A2(new_n614), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n684), .B1(new_n692), .B2(new_n686), .ZN(new_n693));
  XNOR2_X1  g492(.A(G120gat), .B(G148gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G176gat), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(G204gat), .Z(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n691), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n691), .B2(new_n693), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n683), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n589), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n446), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT97), .B(G1gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1324gat));
  OAI21_X1  g505(.A(G8gat), .B1(new_n703), .B2(new_n283), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n708));
  INV_X1    g507(.A(new_n703), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT16), .B(G8gat), .Z(new_n710));
  NAND3_X1  g509(.A1(new_n709), .A2(new_n282), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT98), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n712), .A3(new_n708), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n712), .B1(new_n711), .B2(new_n708), .ZN(new_n715));
  OAI221_X1 g514(.A(new_n707), .B1(new_n708), .B2(new_n711), .C1(new_n714), .C2(new_n715), .ZN(G1325gat));
  INV_X1    g515(.A(G15gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n703), .B2(new_n437), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n718), .A2(KEYINPUT99), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(KEYINPUT99), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n481), .A2(new_n717), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT100), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n719), .A2(new_n720), .B1(new_n709), .B2(new_n722), .ZN(G1326gat));
  XNOR2_X1  g522(.A(new_n422), .B(KEYINPUT77), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n703), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT43), .B(G22gat), .Z(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1327gat));
  NOR2_X1   g526(.A1(new_n635), .A2(new_n701), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n662), .A2(new_n666), .A3(new_n669), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n680), .B1(new_n679), .B2(new_n665), .ZN(new_n730));
  INV_X1    g529(.A(new_n665), .ZN(new_n731));
  AOI211_X1 g530(.A(KEYINPUT95), .B(new_n731), .C1(new_n675), .C2(new_n678), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n729), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n728), .A2(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n734), .A2(G29gat), .A3(new_n446), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n589), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT101), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT45), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n448), .A2(new_n452), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n476), .B(new_n481), .C1(new_n739), .C2(new_n724), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT35), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n432), .A2(new_n437), .A3(KEYINPUT81), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n443), .B1(new_n395), .B2(new_n422), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n741), .B1(new_n744), .B2(new_n739), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n424), .A2(new_n440), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n740), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(KEYINPUT103), .A3(new_n733), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n747), .A2(KEYINPUT103), .A3(KEYINPUT44), .A4(new_n733), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n587), .A2(KEYINPUT102), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT102), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n576), .B2(new_n586), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n728), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n750), .A2(new_n751), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G29gat), .B1(new_n757), .B2(new_n446), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n738), .A2(new_n758), .ZN(G1328gat));
  OAI21_X1  g558(.A(G36gat), .B1(new_n757), .B2(new_n283), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n734), .A2(G36gat), .A3(new_n283), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n589), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT104), .ZN(G1329gat));
  OAI21_X1  g565(.A(G43gat), .B1(new_n757), .B2(new_n481), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n734), .A2(G43gat), .A3(new_n437), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n589), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1330gat));
  OAI21_X1  g571(.A(G50gat), .B1(new_n757), .B2(new_n422), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n734), .A2(new_n724), .A3(G50gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n589), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n773), .A2(KEYINPUT48), .A3(new_n775), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n757), .A2(new_n724), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n777), .A2(G50gat), .B1(new_n589), .B2(new_n774), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n778), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g578(.A(new_n701), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n683), .A2(new_n755), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n747), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(new_n446), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(new_n285), .ZN(G1332gat));
  INV_X1    g583(.A(new_n781), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT105), .B1(new_n486), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT105), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n747), .A2(new_n787), .A3(new_n781), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n283), .ZN(new_n790));
  NOR2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  AND2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n790), .B2(new_n791), .ZN(G1333gat));
  INV_X1    g593(.A(new_n481), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n786), .A2(new_n795), .A3(new_n788), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G71gat), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n437), .A2(G71gat), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT106), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT106), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n797), .A2(new_n803), .A3(new_n800), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT50), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n803), .B1(new_n797), .B2(new_n800), .ZN(new_n806));
  AOI211_X1 g605(.A(KEYINPUT106), .B(new_n799), .C1(new_n796), .C2(G71gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n805), .A2(new_n809), .ZN(G1334gat));
  NOR2_X1   g609(.A1(new_n789), .A2(new_n724), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(G78gat), .Z(G1335gat));
  INV_X1    g611(.A(new_n635), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n813), .B(new_n701), .C1(new_n754), .C2(new_n752), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n814), .B(KEYINPUT107), .Z(new_n815));
  NAND3_X1  g614(.A1(new_n750), .A2(new_n751), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(G85gat), .B1(new_n816), .B2(new_n446), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n755), .A2(new_n635), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n747), .A2(new_n733), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n747), .A2(KEYINPUT51), .A3(new_n733), .A4(new_n818), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n780), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n284), .A3(new_n447), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n817), .A2(new_n824), .ZN(G1336gat));
  OAI21_X1  g624(.A(G92gat), .B1(new_n816), .B2(new_n283), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n821), .A2(KEYINPUT108), .A3(new_n822), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n283), .A2(G92gat), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT108), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n819), .A2(new_n829), .A3(new_n820), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n827), .A2(new_n701), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT52), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(new_n823), .B2(new_n828), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n826), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(G1337gat));
  NAND4_X1  g635(.A1(new_n750), .A2(new_n795), .A3(new_n751), .A4(new_n815), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT109), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G99gat), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n837), .A2(KEYINPUT109), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n821), .A2(new_n822), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n437), .A2(G99gat), .A3(new_n780), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT110), .ZN(new_n843));
  OAI22_X1  g642(.A1(new_n839), .A2(new_n840), .B1(new_n841), .B2(new_n843), .ZN(G1338gat));
  NOR2_X1   g643(.A1(new_n422), .A2(G106gat), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT53), .B1(new_n823), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n750), .A2(new_n432), .A3(new_n751), .A4(new_n815), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT111), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G106gat), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n847), .A2(KEYINPUT111), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G106gat), .B1(new_n816), .B2(new_n724), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n827), .A2(new_n701), .A3(new_n830), .A4(new_n845), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT53), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n851), .A2(new_n855), .ZN(G1339gat));
  INV_X1    g655(.A(KEYINPUT55), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n688), .A2(new_n690), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n684), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n684), .B1(new_n689), .B2(new_n657), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(new_n688), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n857), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n696), .B1(new_n691), .B2(new_n860), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n698), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n858), .A2(new_n860), .A3(new_n684), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n861), .A2(new_n688), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT54), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n866), .B(new_n697), .C1(new_n868), .C2(new_n691), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n857), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n752), .A2(new_n754), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n536), .A2(new_n557), .A3(new_n555), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT112), .ZN(new_n874));
  INV_X1    g673(.A(new_n537), .ZN(new_n875));
  INV_X1    g674(.A(new_n536), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n574), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n565), .A2(new_n566), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n576), .A2(new_n881), .A3(new_n701), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n682), .B1(new_n872), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n865), .A2(new_n870), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n733), .A2(new_n576), .A3(new_n881), .A4(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n635), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n683), .A2(new_n755), .A3(new_n701), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n437), .A2(new_n282), .A3(new_n446), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n888), .A2(new_n587), .A3(new_n724), .A4(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT113), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n890), .A2(new_n891), .A3(G113gat), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n890), .B2(G113gat), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n888), .A2(new_n447), .A3(new_n744), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n283), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n755), .A2(new_n322), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n892), .A2(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT114), .ZN(G1340gat));
  AND2_X1   g697(.A1(new_n888), .A2(new_n724), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n889), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n900), .A2(new_n323), .A3(new_n780), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n894), .A2(new_n283), .A3(new_n701), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n323), .B2(new_n902), .ZN(G1341gat));
  OAI21_X1  g702(.A(G127gat), .B1(new_n900), .B2(new_n813), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n813), .A2(G127gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n895), .B2(new_n905), .ZN(G1342gat));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n907));
  INV_X1    g706(.A(G134gat), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n682), .A2(new_n282), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n894), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT115), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n910), .A2(KEYINPUT115), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n907), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n913), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(KEYINPUT56), .A3(new_n911), .ZN(new_n916));
  OAI21_X1  g715(.A(G134gat), .B1(new_n900), .B2(new_n682), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n914), .A2(new_n916), .A3(new_n917), .ZN(G1343gat));
  NOR2_X1   g717(.A1(new_n588), .A2(G141gat), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n888), .A2(new_n447), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n795), .A2(new_n422), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT118), .B1(new_n920), .B2(new_n921), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n283), .B(new_n919), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT57), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n888), .A2(new_n927), .A3(new_n432), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n282), .A2(new_n446), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n481), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n871), .B1(new_n586), .B2(new_n576), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n682), .B1(new_n882), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n635), .B1(new_n932), .B2(new_n885), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n483), .B1(new_n887), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n930), .B1(new_n934), .B2(KEYINPUT57), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n587), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT58), .B1(new_n937), .B2(G141gat), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n926), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n928), .A2(new_n755), .A3(new_n935), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(KEYINPUT116), .A3(G141gat), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n588), .A2(new_n282), .A3(G141gat), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n888), .A2(new_n447), .A3(new_n921), .A4(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT117), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT116), .B1(new_n940), .B2(G141gat), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n941), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT58), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n939), .B1(new_n947), .B2(new_n948), .ZN(G1344gat));
  XNOR2_X1  g748(.A(new_n922), .B(new_n923), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n283), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n701), .A2(new_n313), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT59), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n587), .A2(new_n884), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n576), .A2(new_n881), .A3(new_n701), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n733), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n884), .A2(new_n576), .A3(new_n881), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n682), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n954), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n932), .A2(new_n885), .A3(KEYINPUT119), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(new_n961), .A3(new_n813), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n683), .A2(new_n587), .A3(new_n701), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n724), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT120), .B1(new_n965), .B2(KEYINPUT57), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT120), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n932), .A2(new_n885), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n635), .B1(new_n968), .B2(new_n954), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n963), .B1(new_n969), .B2(new_n961), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n967), .B(new_n927), .C1(new_n970), .C2(new_n724), .ZN(new_n971));
  OAI211_X1 g770(.A(KEYINPUT57), .B(new_n432), .C1(new_n886), .C2(new_n887), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n966), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n973), .A2(new_n481), .A3(new_n701), .A4(new_n929), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n953), .B1(new_n974), .B2(G148gat), .ZN(new_n975));
  AOI211_X1 g774(.A(KEYINPUT59), .B(new_n313), .C1(new_n936), .C2(new_n701), .ZN(new_n976));
  OAI22_X1  g775(.A1(new_n951), .A2(new_n952), .B1(new_n975), .B2(new_n976), .ZN(G1345gat));
  NAND2_X1  g776(.A1(new_n635), .A2(new_n305), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n936), .A2(new_n635), .ZN(new_n979));
  OAI22_X1  g778(.A1(new_n951), .A2(new_n978), .B1(new_n305), .B2(new_n979), .ZN(G1346gat));
  NAND2_X1  g779(.A1(new_n936), .A2(new_n733), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n306), .B1(new_n981), .B2(KEYINPUT121), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n982), .B1(KEYINPUT121), .B2(new_n981), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n950), .A2(new_n306), .A3(new_n909), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1347gat));
  AND2_X1   g784(.A1(new_n888), .A2(new_n446), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(new_n282), .A3(new_n744), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n987), .A2(new_n227), .A3(new_n755), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n283), .A2(new_n437), .A3(new_n447), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n899), .A2(new_n587), .A3(new_n989), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n990), .A2(KEYINPUT122), .A3(G169gat), .ZN(new_n991));
  AOI21_X1  g790(.A(KEYINPUT122), .B1(new_n990), .B2(G169gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(G1348gat));
  NAND3_X1  g792(.A1(new_n987), .A2(new_n228), .A3(new_n701), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n899), .A2(new_n989), .ZN(new_n995));
  OAI21_X1  g794(.A(G176gat), .B1(new_n995), .B2(new_n780), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n994), .A2(new_n996), .ZN(G1349gat));
  NOR2_X1   g796(.A1(new_n813), .A2(new_n250), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n987), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g798(.A(G183gat), .B1(new_n995), .B2(new_n813), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT123), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(KEYINPUT60), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT60), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1003), .A2(new_n1005), .ZN(G1350gat));
  NAND3_X1  g805(.A1(new_n899), .A2(new_n733), .A3(new_n989), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(G190gat), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(KEYINPUT124), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT124), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1007), .A2(new_n1010), .A3(G190gat), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1009), .A2(KEYINPUT61), .A3(new_n1011), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n682), .A2(new_n218), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n987), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g813(.A(new_n1012), .B(new_n1014), .C1(KEYINPUT61), .C2(new_n1009), .ZN(G1351gat));
  INV_X1    g814(.A(KEYINPUT126), .ZN(new_n1016));
  NOR2_X1   g815(.A1(new_n283), .A2(new_n447), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n481), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g817(.A1(new_n1018), .A2(new_n588), .ZN(new_n1019));
  AND3_X1   g818(.A1(new_n973), .A2(KEYINPUT125), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g819(.A(KEYINPUT125), .B1(new_n973), .B2(new_n1019), .ZN(new_n1021));
  INV_X1    g820(.A(G197gat), .ZN(new_n1022));
  NOR3_X1   g821(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  AND4_X1   g822(.A1(new_n446), .A2(new_n888), .A3(new_n282), .A4(new_n921), .ZN(new_n1024));
  NAND3_X1  g823(.A1(new_n1024), .A2(new_n1022), .A3(new_n755), .ZN(new_n1025));
  INV_X1    g824(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g825(.A(new_n1016), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  AND2_X1   g826(.A1(new_n973), .A2(new_n1019), .ZN(new_n1028));
  OAI21_X1  g827(.A(G197gat), .B1(new_n1028), .B2(KEYINPUT125), .ZN(new_n1029));
  OAI211_X1 g828(.A(KEYINPUT126), .B(new_n1025), .C1(new_n1029), .C2(new_n1020), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1027), .A2(new_n1030), .ZN(G1352gat));
  XNOR2_X1  g830(.A(KEYINPUT127), .B(G204gat), .ZN(new_n1032));
  NOR2_X1   g831(.A1(new_n780), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g832(.A1(new_n1024), .A2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g833(.A(new_n1034), .B(KEYINPUT62), .Z(new_n1035));
  INV_X1    g834(.A(new_n1018), .ZN(new_n1036));
  NAND3_X1  g835(.A1(new_n973), .A2(new_n701), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n1037), .A2(new_n1032), .ZN(new_n1038));
  NAND2_X1  g837(.A1(new_n1035), .A2(new_n1038), .ZN(G1353gat));
  NAND3_X1  g838(.A1(new_n1024), .A2(new_n204), .A3(new_n635), .ZN(new_n1040));
  AND2_X1   g839(.A1(new_n973), .A2(new_n1036), .ZN(new_n1041));
  NAND2_X1  g840(.A1(new_n1041), .A2(new_n635), .ZN(new_n1042));
  AND3_X1   g841(.A1(new_n1042), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1043));
  AOI21_X1  g842(.A(KEYINPUT63), .B1(new_n1042), .B2(G211gat), .ZN(new_n1044));
  OAI21_X1  g843(.A(new_n1040), .B1(new_n1043), .B2(new_n1044), .ZN(G1354gat));
  AOI21_X1  g844(.A(G218gat), .B1(new_n1024), .B2(new_n733), .ZN(new_n1046));
  NOR2_X1   g845(.A1(new_n682), .A2(new_n205), .ZN(new_n1047));
  AOI21_X1  g846(.A(new_n1046), .B1(new_n1041), .B2(new_n1047), .ZN(G1355gat));
endmodule


