

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U550 ( .A1(n642), .A2(n795), .ZN(n644) );
  NOR2_X4 U551 ( .A1(G543), .A2(G651), .ZN(n824) );
  NAND2_X1 U552 ( .A1(n641), .A2(n640), .ZN(n795) );
  NOR2_X4 U553 ( .A1(n605), .A2(n555), .ZN(n631) );
  XOR2_X2 U554 ( .A(KEYINPUT0), .B(G543), .Z(n605) );
  XNOR2_X1 U555 ( .A(n689), .B(KEYINPUT97), .ZN(n690) );
  OR2_X1 U556 ( .A1(n662), .A2(n533), .ZN(n530) );
  OR2_X1 U557 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U558 ( .A1(n537), .A2(n536), .ZN(n535) );
  INV_X1 U559 ( .A(n584), .ZN(n536) );
  NOR2_X1 U560 ( .A1(n583), .A2(n518), .ZN(n537) );
  NOR2_X1 U561 ( .A1(n579), .A2(G2105), .ZN(n727) );
  NAND2_X1 U562 ( .A1(n715), .A2(n998), .ZN(n548) );
  XNOR2_X1 U563 ( .A(n580), .B(KEYINPUT65), .ZN(n732) );
  INV_X1 U564 ( .A(KEYINPUT17), .ZN(n577) );
  NOR2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n578) );
  NOR2_X1 U566 ( .A1(n625), .A2(n935), .ZN(n627) );
  NAND2_X1 U567 ( .A1(n519), .A2(n530), .ZN(n529) );
  NAND2_X1 U568 ( .A1(G171), .A2(n685), .ZN(n678) );
  INV_X1 U569 ( .A(n994), .ZN(n706) );
  INV_X1 U570 ( .A(n696), .ZN(n544) );
  INV_X1 U571 ( .A(G2104), .ZN(n579) );
  XNOR2_X1 U572 ( .A(n558), .B(n557), .ZN(n648) );
  XNOR2_X1 U573 ( .A(n556), .B(KEYINPUT1), .ZN(n557) );
  INV_X1 U574 ( .A(KEYINPUT66), .ZN(n556) );
  XNOR2_X1 U575 ( .A(n546), .B(KEYINPUT103), .ZN(n762) );
  NAND2_X1 U576 ( .A1(n547), .A2(n524), .ZN(n546) );
  NAND2_X1 U577 ( .A1(n548), .A2(n521), .ZN(n547) );
  XOR2_X1 U578 ( .A(KEYINPUT15), .B(n654), .Z(n983) );
  NOR2_X1 U579 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U580 ( .A1(n517), .A2(n534), .ZN(n539) );
  XNOR2_X1 U581 ( .A(n585), .B(KEYINPUT80), .ZN(n534) );
  NAND2_X1 U582 ( .A1(n732), .A2(G126), .ZN(n585) );
  XNOR2_X1 U583 ( .A(n574), .B(n573), .ZN(n576) );
  INV_X1 U584 ( .A(KEYINPUT23), .ZN(n573) );
  NAND2_X2 U585 ( .A1(n535), .A2(n539), .ZN(n625) );
  AND2_X1 U586 ( .A1(n659), .A2(KEYINPUT93), .ZN(n516) );
  INV_X1 U587 ( .A(n539), .ZN(G164) );
  AND2_X1 U588 ( .A1(n589), .A2(n588), .ZN(n517) );
  NAND2_X1 U589 ( .A1(n538), .A2(G40), .ZN(n518) );
  XOR2_X1 U590 ( .A(n667), .B(KEYINPUT94), .Z(n519) );
  AND2_X1 U591 ( .A1(n662), .A2(n533), .ZN(n520) );
  AND2_X1 U592 ( .A1(n724), .A2(n723), .ZN(n521) );
  AND2_X1 U593 ( .A1(n697), .A2(n695), .ZN(n522) );
  AND2_X1 U594 ( .A1(n707), .A2(n706), .ZN(n523) );
  AND2_X1 U595 ( .A1(n771), .A2(n759), .ZN(n524) );
  AND2_X1 U596 ( .A1(n550), .A2(n990), .ZN(n525) );
  NAND2_X1 U597 ( .A1(n712), .A2(KEYINPUT33), .ZN(n526) );
  INV_X1 U598 ( .A(KEYINPUT93), .ZN(n533) );
  NAND2_X1 U599 ( .A1(n527), .A2(n532), .ZN(n531) );
  NAND2_X1 U600 ( .A1(n528), .A2(n520), .ZN(n527) );
  NAND2_X1 U601 ( .A1(n660), .A2(n659), .ZN(n528) );
  NAND2_X1 U602 ( .A1(n660), .A2(n516), .ZN(n532) );
  NOR2_X2 U603 ( .A1(n531), .A2(n529), .ZN(n668) );
  NOR2_X1 U604 ( .A1(n584), .A2(n583), .ZN(G160) );
  NAND2_X1 U605 ( .A1(G160), .A2(G40), .ZN(n726) );
  NOR2_X1 U606 ( .A1(G164), .A2(G1384), .ZN(n725) );
  INV_X1 U607 ( .A(G1384), .ZN(n538) );
  NAND2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n522), .A2(n544), .ZN(n540) );
  XNOR2_X1 U610 ( .A(n705), .B(n545), .ZN(n541) );
  NAND2_X1 U611 ( .A1(n542), .A2(n525), .ZN(n713) );
  NAND2_X1 U612 ( .A1(n543), .A2(n523), .ZN(n542) );
  INV_X1 U613 ( .A(KEYINPUT32), .ZN(n545) );
  XNOR2_X1 U614 ( .A(KEYINPUT28), .B(n670), .ZN(n549) );
  NOR2_X1 U615 ( .A1(n721), .A2(n711), .ZN(n550) );
  INV_X1 U616 ( .A(KEYINPUT26), .ZN(n626) );
  INV_X1 U617 ( .A(KEYINPUT64), .ZN(n643) );
  INV_X1 U618 ( .A(KEYINPUT92), .ZN(n655) );
  NAND2_X1 U619 ( .A1(n661), .A2(n983), .ZN(n662) );
  INV_X1 U620 ( .A(KEYINPUT29), .ZN(n672) );
  INV_X1 U621 ( .A(KEYINPUT13), .ZN(n635) );
  XNOR2_X1 U622 ( .A(n649), .B(KEYINPUT71), .ZN(n650) );
  AND2_X2 U623 ( .A1(G2104), .A2(G2105), .ZN(n906) );
  NAND2_X1 U624 ( .A1(n824), .A2(G89), .ZN(n551) );
  XNOR2_X1 U625 ( .A(n551), .B(KEYINPUT4), .ZN(n553) );
  INV_X1 U626 ( .A(G651), .ZN(n555) );
  NAND2_X1 U627 ( .A1(G76), .A2(n631), .ZN(n552) );
  NAND2_X1 U628 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U629 ( .A(n554), .B(KEYINPUT5), .ZN(n563) );
  NOR2_X2 U630 ( .A1(n605), .A2(G651), .ZN(n820) );
  NAND2_X1 U631 ( .A1(n820), .A2(G51), .ZN(n560) );
  NOR2_X1 U632 ( .A1(G543), .A2(n555), .ZN(n558) );
  BUF_X1 U633 ( .A(n648), .Z(n821) );
  NAND2_X1 U634 ( .A1(G63), .A2(n821), .ZN(n559) );
  NAND2_X1 U635 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U636 ( .A(KEYINPUT6), .B(n561), .Z(n562) );
  NAND2_X1 U637 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U638 ( .A(n564), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U639 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U640 ( .A1(n820), .A2(G52), .ZN(n566) );
  NAND2_X1 U641 ( .A1(G64), .A2(n821), .ZN(n565) );
  NAND2_X1 U642 ( .A1(n566), .A2(n565), .ZN(n572) );
  NAND2_X1 U643 ( .A1(G90), .A2(n824), .ZN(n568) );
  NAND2_X1 U644 ( .A1(G77), .A2(n631), .ZN(n567) );
  NAND2_X1 U645 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U646 ( .A(KEYINPUT67), .B(n569), .ZN(n570) );
  XNOR2_X1 U647 ( .A(KEYINPUT9), .B(n570), .ZN(n571) );
  NOR2_X1 U648 ( .A1(n572), .A2(n571), .ZN(G171) );
  NAND2_X1 U649 ( .A1(n727), .A2(G101), .ZN(n574) );
  NAND2_X1 U650 ( .A1(n906), .A2(G113), .ZN(n575) );
  NAND2_X1 U651 ( .A1(n576), .A2(n575), .ZN(n584) );
  XNOR2_X2 U652 ( .A(n578), .B(n577), .ZN(n728) );
  NAND2_X1 U653 ( .A1(n728), .A2(G137), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n579), .A2(G2105), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n732), .A2(G125), .ZN(n581) );
  NAND2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U657 ( .A1(G102), .A2(n727), .ZN(n587) );
  NAND2_X1 U658 ( .A1(G114), .A2(n906), .ZN(n586) );
  AND2_X1 U659 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U660 ( .A1(n728), .A2(G138), .ZN(n588) );
  NAND2_X1 U661 ( .A1(G91), .A2(n824), .ZN(n591) );
  NAND2_X1 U662 ( .A1(G78), .A2(n631), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U664 ( .A1(n820), .A2(G53), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G65), .A2(n821), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n594) );
  OR2_X1 U667 ( .A1(n595), .A2(n594), .ZN(G299) );
  NAND2_X1 U668 ( .A1(G88), .A2(n824), .ZN(n597) );
  NAND2_X1 U669 ( .A1(G75), .A2(n631), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n820), .A2(G50), .ZN(n599) );
  NAND2_X1 U672 ( .A1(G62), .A2(n821), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U674 ( .A1(n601), .A2(n600), .ZN(G166) );
  INV_X1 U675 ( .A(G166), .ZN(G303) );
  NAND2_X1 U676 ( .A1(G49), .A2(n820), .ZN(n603) );
  NAND2_X1 U677 ( .A1(G74), .A2(G651), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U679 ( .A1(n821), .A2(n604), .ZN(n608) );
  NAND2_X1 U680 ( .A1(G87), .A2(n605), .ZN(n606) );
  XOR2_X1 U681 ( .A(KEYINPUT75), .B(n606), .Z(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(G288) );
  NAND2_X1 U683 ( .A1(G73), .A2(n631), .ZN(n609) );
  XNOR2_X1 U684 ( .A(n609), .B(KEYINPUT2), .ZN(n616) );
  NAND2_X1 U685 ( .A1(G86), .A2(n824), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G48), .A2(n820), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n821), .A2(G61), .ZN(n612) );
  XOR2_X1 U689 ( .A(KEYINPUT76), .B(n612), .Z(n613) );
  NOR2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(G305) );
  NAND2_X1 U692 ( .A1(G85), .A2(n824), .ZN(n618) );
  NAND2_X1 U693 ( .A1(G60), .A2(n821), .ZN(n617) );
  NAND2_X1 U694 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U695 ( .A1(G72), .A2(n631), .ZN(n620) );
  NAND2_X1 U696 ( .A1(G47), .A2(n820), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n621) );
  OR2_X1 U698 ( .A1(n622), .A2(n621), .ZN(G290) );
  NAND2_X1 U699 ( .A1(G8), .A2(n625), .ZN(n721) );
  NOR2_X1 U700 ( .A1(G1966), .A2(n721), .ZN(n696) );
  INV_X1 U701 ( .A(G1996), .ZN(n935) );
  XNOR2_X1 U702 ( .A(n627), .B(n626), .ZN(n629) );
  NAND2_X1 U703 ( .A1(n625), .A2(G1341), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n642) );
  NAND2_X1 U705 ( .A1(G56), .A2(n648), .ZN(n630) );
  XOR2_X1 U706 ( .A(KEYINPUT14), .B(n630), .Z(n638) );
  NAND2_X1 U707 ( .A1(G68), .A2(n631), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n824), .A2(G81), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(KEYINPUT12), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U712 ( .A(n639), .B(KEYINPUT70), .ZN(n641) );
  NAND2_X1 U713 ( .A1(G43), .A2(n820), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(n661) );
  NAND2_X1 U715 ( .A1(G92), .A2(n824), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n645), .B(KEYINPUT72), .ZN(n653) );
  NAND2_X1 U717 ( .A1(G79), .A2(n631), .ZN(n647) );
  NAND2_X1 U718 ( .A1(G54), .A2(n820), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U720 ( .A1(G66), .A2(n648), .ZN(n649) );
  NOR2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U722 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U723 ( .A1(n661), .A2(n983), .ZN(n656) );
  XNOR2_X1 U724 ( .A(n656), .B(n655), .ZN(n660) );
  NOR2_X1 U725 ( .A1(G2067), .A2(n625), .ZN(n658) );
  INV_X1 U726 ( .A(n625), .ZN(n675) );
  NOR2_X1 U727 ( .A1(n675), .A2(G1348), .ZN(n657) );
  NOR2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n659) );
  INV_X1 U729 ( .A(G2072), .ZN(n1021) );
  NOR2_X1 U730 ( .A1(n625), .A2(n1021), .ZN(n664) );
  XNOR2_X1 U731 ( .A(KEYINPUT27), .B(KEYINPUT90), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n664), .B(n663), .ZN(n666) );
  XOR2_X1 U733 ( .A(G1956), .B(KEYINPUT91), .Z(n958) );
  NAND2_X1 U734 ( .A1(n625), .A2(n958), .ZN(n665) );
  NAND2_X1 U735 ( .A1(n666), .A2(n665), .ZN(n669) );
  NOR2_X1 U736 ( .A1(G299), .A2(n669), .ZN(n667) );
  XNOR2_X1 U737 ( .A(n668), .B(KEYINPUT95), .ZN(n671) );
  NAND2_X1 U738 ( .A1(G299), .A2(n669), .ZN(n670) );
  NAND2_X1 U739 ( .A1(n671), .A2(n549), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n673), .B(n672), .ZN(n679) );
  XOR2_X1 U741 ( .A(G2078), .B(KEYINPUT25), .Z(n674) );
  XNOR2_X1 U742 ( .A(KEYINPUT89), .B(n674), .ZN(n936) );
  NOR2_X1 U743 ( .A1(n625), .A2(n936), .ZN(n677) );
  XOR2_X1 U744 ( .A(G1961), .B(KEYINPUT88), .Z(n956) );
  NOR2_X1 U745 ( .A1(n675), .A2(n956), .ZN(n676) );
  NOR2_X1 U746 ( .A1(n677), .A2(n676), .ZN(n685) );
  NAND2_X1 U747 ( .A1(n679), .A2(n678), .ZN(n691) );
  NOR2_X1 U748 ( .A1(n625), .A2(G2084), .ZN(n680) );
  XNOR2_X1 U749 ( .A(n680), .B(KEYINPUT87), .ZN(n693) );
  NAND2_X1 U750 ( .A1(G8), .A2(n693), .ZN(n681) );
  NOR2_X1 U751 ( .A1(n696), .A2(n681), .ZN(n683) );
  XOR2_X1 U752 ( .A(KEYINPUT96), .B(KEYINPUT30), .Z(n682) );
  XNOR2_X1 U753 ( .A(n683), .B(n682), .ZN(n684) );
  NOR2_X1 U754 ( .A1(G168), .A2(n684), .ZN(n687) );
  NOR2_X1 U755 ( .A1(G171), .A2(n685), .ZN(n686) );
  NOR2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U757 ( .A(n688), .B(KEYINPUT31), .ZN(n689) );
  NAND2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U759 ( .A(n692), .B(KEYINPUT98), .ZN(n697) );
  INV_X1 U760 ( .A(n693), .ZN(n694) );
  NAND2_X1 U761 ( .A1(G8), .A2(n694), .ZN(n695) );
  NAND2_X1 U762 ( .A1(n697), .A2(G286), .ZN(n704) );
  INV_X1 U763 ( .A(G8), .ZN(n702) );
  NOR2_X1 U764 ( .A1(G1971), .A2(n721), .ZN(n699) );
  NOR2_X1 U765 ( .A1(G2090), .A2(n625), .ZN(n698) );
  NOR2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U767 ( .A1(n700), .A2(G303), .ZN(n701) );
  NAND2_X1 U768 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U769 ( .A1(G1971), .A2(G303), .ZN(n993) );
  XNOR2_X1 U770 ( .A(n993), .B(KEYINPUT99), .ZN(n707) );
  NOR2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n994) );
  NAND2_X1 U772 ( .A1(KEYINPUT33), .A2(n994), .ZN(n708) );
  NOR2_X1 U773 ( .A1(n721), .A2(n708), .ZN(n709) );
  XOR2_X1 U774 ( .A(KEYINPUT101), .B(n709), .Z(n711) );
  NAND2_X1 U775 ( .A1(G288), .A2(G1976), .ZN(n710) );
  XNOR2_X1 U776 ( .A(n710), .B(KEYINPUT100), .ZN(n990) );
  INV_X1 U777 ( .A(n711), .ZN(n712) );
  NAND2_X1 U778 ( .A1(n713), .A2(n526), .ZN(n714) );
  XNOR2_X1 U779 ( .A(n714), .B(KEYINPUT102), .ZN(n715) );
  XOR2_X1 U780 ( .A(G1981), .B(G305), .Z(n998) );
  NOR2_X1 U781 ( .A1(G2090), .A2(G303), .ZN(n716) );
  NAND2_X1 U782 ( .A1(G8), .A2(n716), .ZN(n717) );
  NAND2_X1 U783 ( .A1(n543), .A2(n717), .ZN(n718) );
  NAND2_X1 U784 ( .A1(n721), .A2(n718), .ZN(n724) );
  NOR2_X1 U785 ( .A1(G1981), .A2(G305), .ZN(n719) );
  XOR2_X1 U786 ( .A(n719), .B(KEYINPUT24), .Z(n720) );
  NOR2_X1 U787 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U788 ( .A(n722), .B(KEYINPUT86), .Z(n723) );
  NOR2_X1 U789 ( .A1(n725), .A2(n726), .ZN(n775) );
  BUF_X1 U790 ( .A(n727), .Z(n910) );
  NAND2_X1 U791 ( .A1(G104), .A2(n910), .ZN(n730) );
  NAND2_X1 U792 ( .A1(G140), .A2(n728), .ZN(n729) );
  NAND2_X1 U793 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U794 ( .A(KEYINPUT34), .B(n731), .ZN(n739) );
  NAND2_X1 U795 ( .A1(G116), .A2(n906), .ZN(n735) );
  BUF_X1 U796 ( .A(n732), .Z(n733) );
  NAND2_X1 U797 ( .A1(G128), .A2(n733), .ZN(n734) );
  NAND2_X1 U798 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U799 ( .A(KEYINPUT35), .B(n736), .Z(n737) );
  XNOR2_X1 U800 ( .A(KEYINPUT82), .B(n737), .ZN(n738) );
  NOR2_X1 U801 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U802 ( .A(KEYINPUT36), .B(n740), .ZN(n920) );
  XNOR2_X1 U803 ( .A(G2067), .B(KEYINPUT37), .ZN(n773) );
  NOR2_X1 U804 ( .A1(n920), .A2(n773), .ZN(n1015) );
  NAND2_X1 U805 ( .A1(n775), .A2(n1015), .ZN(n771) );
  NAND2_X1 U806 ( .A1(G117), .A2(n906), .ZN(n742) );
  NAND2_X1 U807 ( .A1(G129), .A2(n733), .ZN(n741) );
  NAND2_X1 U808 ( .A1(n742), .A2(n741), .ZN(n746) );
  NAND2_X1 U809 ( .A1(G105), .A2(n910), .ZN(n743) );
  XNOR2_X1 U810 ( .A(n743), .B(KEYINPUT85), .ZN(n744) );
  XNOR2_X1 U811 ( .A(n744), .B(KEYINPUT38), .ZN(n745) );
  NOR2_X1 U812 ( .A1(n746), .A2(n745), .ZN(n748) );
  NAND2_X1 U813 ( .A1(n728), .A2(G141), .ZN(n747) );
  NAND2_X1 U814 ( .A1(n748), .A2(n747), .ZN(n892) );
  NAND2_X1 U815 ( .A1(G1996), .A2(n892), .ZN(n758) );
  NAND2_X1 U816 ( .A1(G131), .A2(n728), .ZN(n749) );
  XNOR2_X1 U817 ( .A(n749), .B(KEYINPUT84), .ZN(n756) );
  NAND2_X1 U818 ( .A1(G107), .A2(n906), .ZN(n751) );
  NAND2_X1 U819 ( .A1(G119), .A2(n733), .ZN(n750) );
  NAND2_X1 U820 ( .A1(n751), .A2(n750), .ZN(n754) );
  NAND2_X1 U821 ( .A1(G95), .A2(n910), .ZN(n752) );
  XNOR2_X1 U822 ( .A(KEYINPUT83), .B(n752), .ZN(n753) );
  NOR2_X1 U823 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U824 ( .A1(n756), .A2(n755), .ZN(n889) );
  NAND2_X1 U825 ( .A1(G1991), .A2(n889), .ZN(n757) );
  NAND2_X1 U826 ( .A1(n758), .A2(n757), .ZN(n1016) );
  NAND2_X1 U827 ( .A1(n775), .A2(n1016), .ZN(n759) );
  XOR2_X1 U828 ( .A(KEYINPUT81), .B(G1986), .Z(n760) );
  XNOR2_X1 U829 ( .A(G290), .B(n760), .ZN(n992) );
  NAND2_X1 U830 ( .A1(n992), .A2(n775), .ZN(n761) );
  NAND2_X1 U831 ( .A1(n762), .A2(n761), .ZN(n778) );
  XOR2_X1 U832 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n770) );
  NOR2_X1 U833 ( .A1(G1996), .A2(n892), .ZN(n1026) );
  NOR2_X1 U834 ( .A1(G1991), .A2(n889), .ZN(n1011) );
  NOR2_X1 U835 ( .A1(G1986), .A2(G290), .ZN(n763) );
  XNOR2_X1 U836 ( .A(KEYINPUT104), .B(n763), .ZN(n764) );
  NOR2_X1 U837 ( .A1(n1011), .A2(n764), .ZN(n765) );
  XOR2_X1 U838 ( .A(KEYINPUT105), .B(n765), .Z(n766) );
  NOR2_X1 U839 ( .A1(n1016), .A2(n766), .ZN(n767) );
  XNOR2_X1 U840 ( .A(n767), .B(KEYINPUT106), .ZN(n768) );
  NOR2_X1 U841 ( .A1(n1026), .A2(n768), .ZN(n769) );
  XNOR2_X1 U842 ( .A(n770), .B(n769), .ZN(n772) );
  NAND2_X1 U843 ( .A1(n772), .A2(n771), .ZN(n774) );
  NAND2_X1 U844 ( .A1(n920), .A2(n773), .ZN(n1030) );
  NAND2_X1 U845 ( .A1(n774), .A2(n1030), .ZN(n776) );
  NAND2_X1 U846 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U847 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U848 ( .A(n779), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U849 ( .A(G2451), .B(G2446), .ZN(n789) );
  XOR2_X1 U850 ( .A(G2430), .B(KEYINPUT109), .Z(n781) );
  XNOR2_X1 U851 ( .A(G2454), .B(G2435), .ZN(n780) );
  XNOR2_X1 U852 ( .A(n781), .B(n780), .ZN(n785) );
  XOR2_X1 U853 ( .A(G2438), .B(KEYINPUT108), .Z(n783) );
  XNOR2_X1 U854 ( .A(G1341), .B(G1348), .ZN(n782) );
  XNOR2_X1 U855 ( .A(n783), .B(n782), .ZN(n784) );
  XOR2_X1 U856 ( .A(n785), .B(n784), .Z(n787) );
  XNOR2_X1 U857 ( .A(G2443), .B(G2427), .ZN(n786) );
  XNOR2_X1 U858 ( .A(n787), .B(n786), .ZN(n788) );
  XNOR2_X1 U859 ( .A(n789), .B(n788), .ZN(n790) );
  AND2_X1 U860 ( .A1(n790), .A2(G14), .ZN(G401) );
  AND2_X1 U861 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U862 ( .A(G57), .ZN(G237) );
  XOR2_X1 U863 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n792) );
  NAND2_X1 U864 ( .A1(G7), .A2(G661), .ZN(n791) );
  XNOR2_X1 U865 ( .A(n792), .B(n791), .ZN(n793) );
  XNOR2_X1 U866 ( .A(KEYINPUT68), .B(n793), .ZN(G223) );
  INV_X1 U867 ( .A(G223), .ZN(n856) );
  NAND2_X1 U868 ( .A1(n856), .A2(G567), .ZN(n794) );
  XOR2_X1 U869 ( .A(KEYINPUT11), .B(n794), .Z(G234) );
  INV_X1 U870 ( .A(G860), .ZN(n800) );
  OR2_X1 U871 ( .A1(n795), .A2(n800), .ZN(G153) );
  INV_X1 U872 ( .A(G171), .ZN(G301) );
  NAND2_X1 U873 ( .A1(G868), .A2(G301), .ZN(n797) );
  INV_X1 U874 ( .A(G868), .ZN(n803) );
  NAND2_X1 U875 ( .A1(n983), .A2(n803), .ZN(n796) );
  NAND2_X1 U876 ( .A1(n797), .A2(n796), .ZN(G284) );
  NOR2_X1 U877 ( .A1(G286), .A2(n803), .ZN(n799) );
  NOR2_X1 U878 ( .A1(G868), .A2(G299), .ZN(n798) );
  NOR2_X1 U879 ( .A1(n799), .A2(n798), .ZN(G297) );
  NAND2_X1 U880 ( .A1(n800), .A2(G559), .ZN(n801) );
  INV_X1 U881 ( .A(n983), .ZN(n818) );
  NAND2_X1 U882 ( .A1(n801), .A2(n818), .ZN(n802) );
  XNOR2_X1 U883 ( .A(n802), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U884 ( .A1(n983), .A2(n803), .ZN(n804) );
  XNOR2_X1 U885 ( .A(n804), .B(KEYINPUT73), .ZN(n805) );
  NOR2_X1 U886 ( .A1(G559), .A2(n805), .ZN(n807) );
  NOR2_X1 U887 ( .A1(G868), .A2(n795), .ZN(n806) );
  NOR2_X1 U888 ( .A1(n807), .A2(n806), .ZN(G282) );
  NAND2_X1 U889 ( .A1(G99), .A2(n910), .ZN(n809) );
  NAND2_X1 U890 ( .A1(G111), .A2(n906), .ZN(n808) );
  NAND2_X1 U891 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U892 ( .A(KEYINPUT74), .B(n810), .ZN(n815) );
  NAND2_X1 U893 ( .A1(n733), .A2(G123), .ZN(n811) );
  XNOR2_X1 U894 ( .A(n811), .B(KEYINPUT18), .ZN(n813) );
  NAND2_X1 U895 ( .A1(G135), .A2(n728), .ZN(n812) );
  NAND2_X1 U896 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U897 ( .A1(n815), .A2(n814), .ZN(n1010) );
  XNOR2_X1 U898 ( .A(n1010), .B(G2096), .ZN(n817) );
  INV_X1 U899 ( .A(G2100), .ZN(n816) );
  NAND2_X1 U900 ( .A1(n817), .A2(n816), .ZN(G156) );
  NAND2_X1 U901 ( .A1(n818), .A2(G559), .ZN(n838) );
  XNOR2_X1 U902 ( .A(n795), .B(n838), .ZN(n819) );
  NOR2_X1 U903 ( .A1(n819), .A2(G860), .ZN(n829) );
  NAND2_X1 U904 ( .A1(n820), .A2(G55), .ZN(n823) );
  NAND2_X1 U905 ( .A1(G67), .A2(n821), .ZN(n822) );
  NAND2_X1 U906 ( .A1(n823), .A2(n822), .ZN(n828) );
  NAND2_X1 U907 ( .A1(G93), .A2(n824), .ZN(n826) );
  NAND2_X1 U908 ( .A1(G80), .A2(n631), .ZN(n825) );
  NAND2_X1 U909 ( .A1(n826), .A2(n825), .ZN(n827) );
  NOR2_X1 U910 ( .A1(n828), .A2(n827), .ZN(n831) );
  XNOR2_X1 U911 ( .A(n829), .B(n831), .ZN(G145) );
  NOR2_X1 U912 ( .A1(G868), .A2(n831), .ZN(n830) );
  XOR2_X1 U913 ( .A(KEYINPUT78), .B(n830), .Z(n842) );
  XNOR2_X1 U914 ( .A(n831), .B(G290), .ZN(n832) );
  XNOR2_X1 U915 ( .A(n832), .B(n795), .ZN(n833) );
  XNOR2_X1 U916 ( .A(KEYINPUT19), .B(n833), .ZN(n835) );
  XNOR2_X1 U917 ( .A(G305), .B(G166), .ZN(n834) );
  XNOR2_X1 U918 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U919 ( .A(n836), .B(G288), .Z(n837) );
  XNOR2_X1 U920 ( .A(G299), .B(n837), .ZN(n923) );
  XNOR2_X1 U921 ( .A(n923), .B(n838), .ZN(n839) );
  NAND2_X1 U922 ( .A1(n839), .A2(G868), .ZN(n840) );
  XOR2_X1 U923 ( .A(KEYINPUT77), .B(n840), .Z(n841) );
  NAND2_X1 U924 ( .A1(n842), .A2(n841), .ZN(G295) );
  NAND2_X1 U925 ( .A1(G2078), .A2(G2084), .ZN(n843) );
  XOR2_X1 U926 ( .A(KEYINPUT20), .B(n843), .Z(n844) );
  NAND2_X1 U927 ( .A1(G2090), .A2(n844), .ZN(n845) );
  XNOR2_X1 U928 ( .A(KEYINPUT21), .B(n845), .ZN(n846) );
  NAND2_X1 U929 ( .A1(n846), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U930 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U931 ( .A(KEYINPUT22), .B(KEYINPUT79), .Z(n848) );
  NAND2_X1 U932 ( .A1(G132), .A2(G82), .ZN(n847) );
  XNOR2_X1 U933 ( .A(n848), .B(n847), .ZN(n849) );
  NOR2_X1 U934 ( .A1(n849), .A2(G218), .ZN(n850) );
  NAND2_X1 U935 ( .A1(G96), .A2(n850), .ZN(n861) );
  NAND2_X1 U936 ( .A1(n861), .A2(G2106), .ZN(n854) );
  NAND2_X1 U937 ( .A1(G69), .A2(G120), .ZN(n851) );
  NOR2_X1 U938 ( .A1(G237), .A2(n851), .ZN(n852) );
  NAND2_X1 U939 ( .A1(G108), .A2(n852), .ZN(n862) );
  NAND2_X1 U940 ( .A1(n862), .A2(G567), .ZN(n853) );
  NAND2_X1 U941 ( .A1(n854), .A2(n853), .ZN(n863) );
  NAND2_X1 U942 ( .A1(G661), .A2(G483), .ZN(n855) );
  NOR2_X1 U943 ( .A1(n863), .A2(n855), .ZN(n858) );
  NAND2_X1 U944 ( .A1(n858), .A2(G36), .ZN(G176) );
  NAND2_X1 U945 ( .A1(G2106), .A2(n856), .ZN(G217) );
  AND2_X1 U946 ( .A1(G15), .A2(G2), .ZN(n857) );
  NAND2_X1 U947 ( .A1(G661), .A2(n857), .ZN(G259) );
  NAND2_X1 U948 ( .A1(G1), .A2(G3), .ZN(n859) );
  NAND2_X1 U949 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U950 ( .A(n860), .B(KEYINPUT110), .ZN(G188) );
  INV_X1 U952 ( .A(G132), .ZN(G219) );
  INV_X1 U953 ( .A(G120), .ZN(G236) );
  INV_X1 U954 ( .A(G96), .ZN(G221) );
  INV_X1 U955 ( .A(G82), .ZN(G220) );
  INV_X1 U956 ( .A(G69), .ZN(G235) );
  NOR2_X1 U957 ( .A1(n862), .A2(n861), .ZN(G325) );
  INV_X1 U958 ( .A(G325), .ZN(G261) );
  INV_X1 U959 ( .A(n863), .ZN(G319) );
  XOR2_X1 U960 ( .A(G2100), .B(G2096), .Z(n865) );
  XNOR2_X1 U961 ( .A(KEYINPUT42), .B(G2678), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U963 ( .A(KEYINPUT43), .B(G2090), .Z(n867) );
  XNOR2_X1 U964 ( .A(G2067), .B(G2072), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U966 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U967 ( .A(G2078), .B(G2084), .ZN(n870) );
  XNOR2_X1 U968 ( .A(n871), .B(n870), .ZN(G227) );
  XOR2_X1 U969 ( .A(G1996), .B(G1961), .Z(n873) );
  XNOR2_X1 U970 ( .A(G1981), .B(G1966), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n873), .B(n872), .ZN(n877) );
  XOR2_X1 U972 ( .A(G1971), .B(G1956), .Z(n875) );
  XNOR2_X1 U973 ( .A(G1986), .B(G1976), .ZN(n874) );
  XNOR2_X1 U974 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U975 ( .A(n877), .B(n876), .Z(n879) );
  XNOR2_X1 U976 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n879), .B(n878), .ZN(n881) );
  XOR2_X1 U978 ( .A(G1991), .B(G2474), .Z(n880) );
  XNOR2_X1 U979 ( .A(n881), .B(n880), .ZN(G229) );
  NAND2_X1 U980 ( .A1(G100), .A2(n910), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G112), .A2(n906), .ZN(n882) );
  NAND2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n888) );
  NAND2_X1 U983 ( .A1(G124), .A2(n733), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n884), .B(KEYINPUT44), .ZN(n886) );
  NAND2_X1 U985 ( .A1(n728), .A2(G136), .ZN(n885) );
  NAND2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n887) );
  NOR2_X1 U987 ( .A1(n888), .A2(n887), .ZN(G162) );
  XNOR2_X1 U988 ( .A(n889), .B(G162), .ZN(n891) );
  XNOR2_X1 U989 ( .A(G160), .B(G164), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n891), .B(n890), .ZN(n896) );
  XNOR2_X1 U991 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n892), .B(n1010), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U994 ( .A(n896), .B(n895), .Z(n919) );
  NAND2_X1 U995 ( .A1(G103), .A2(n910), .ZN(n898) );
  NAND2_X1 U996 ( .A1(G139), .A2(n728), .ZN(n897) );
  NAND2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n905) );
  NAND2_X1 U998 ( .A1(n906), .A2(G115), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n899), .B(KEYINPUT114), .ZN(n901) );
  NAND2_X1 U1000 ( .A1(G127), .A2(n733), .ZN(n900) );
  NAND2_X1 U1001 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(KEYINPUT47), .B(n902), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(KEYINPUT115), .B(n903), .ZN(n904) );
  NOR2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(n1020) );
  NAND2_X1 U1005 ( .A1(G118), .A2(n906), .ZN(n908) );
  NAND2_X1 U1006 ( .A1(G130), .A2(n733), .ZN(n907) );
  NAND2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(KEYINPUT112), .B(n909), .ZN(n916) );
  NAND2_X1 U1009 ( .A1(G106), .A2(n910), .ZN(n912) );
  NAND2_X1 U1010 ( .A1(G142), .A2(n728), .ZN(n911) );
  NAND2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(KEYINPUT45), .B(n913), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(KEYINPUT113), .B(n914), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(n1020), .B(n917), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n919), .B(n918), .ZN(n921) );
  XOR2_X1 U1017 ( .A(n921), .B(n920), .Z(n922) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n922), .ZN(G395) );
  XNOR2_X1 U1019 ( .A(G286), .B(n983), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(n924), .B(n923), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(n925), .B(G171), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(G37), .A2(n926), .ZN(G397) );
  NOR2_X1 U1023 ( .A1(G227), .A2(G229), .ZN(n927) );
  XOR2_X1 U1024 ( .A(KEYINPUT49), .B(n927), .Z(n928) );
  NAND2_X1 U1025 ( .A1(G319), .A2(n928), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(G401), .A2(n929), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(KEYINPUT116), .B(n930), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(G395), .A2(G397), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(G225) );
  INV_X1 U1030 ( .A(G225), .ZN(G308) );
  INV_X1 U1031 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1032 ( .A(G2084), .B(G34), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(n933), .B(KEYINPUT54), .ZN(n951) );
  XNOR2_X1 U1034 ( .A(G2090), .B(G35), .ZN(n948) );
  XOR2_X1 U1035 ( .A(G1991), .B(G25), .Z(n934) );
  NAND2_X1 U1036 ( .A1(n934), .A2(G28), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(n935), .B(G32), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(n936), .B(G27), .ZN(n937) );
  NAND2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1040 ( .A(KEYINPUT121), .B(n939), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(G2067), .B(G26), .ZN(n941) );
  XNOR2_X1 U1042 ( .A(G2072), .B(G33), .ZN(n940) );
  NOR2_X1 U1043 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1046 ( .A(KEYINPUT53), .B(n946), .ZN(n947) );
  NOR2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1048 ( .A(KEYINPUT122), .B(n949), .Z(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1050 ( .A(KEYINPUT123), .B(n952), .Z(n953) );
  NOR2_X1 U1051 ( .A1(G29), .A2(n953), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(KEYINPUT55), .B(n954), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(n955), .B(KEYINPUT120), .ZN(n1042) );
  XNOR2_X1 U1054 ( .A(n956), .B(G5), .ZN(n970) );
  XNOR2_X1 U1055 ( .A(G1348), .B(KEYINPUT59), .ZN(n957) );
  XNOR2_X1 U1056 ( .A(n957), .B(G4), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(G1341), .B(G19), .ZN(n960) );
  XNOR2_X1 U1058 ( .A(n958), .B(G20), .ZN(n959) );
  NOR2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(KEYINPUT126), .B(G1981), .ZN(n963) );
  XNOR2_X1 U1062 ( .A(G6), .B(n963), .ZN(n964) );
  NOR2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1064 ( .A(KEYINPUT60), .B(n966), .Z(n968) );
  XNOR2_X1 U1065 ( .A(G1966), .B(G21), .ZN(n967) );
  NOR2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(G1986), .B(G24), .ZN(n972) );
  XNOR2_X1 U1069 ( .A(G22), .B(G1971), .ZN(n971) );
  NOR2_X1 U1070 ( .A1(n972), .A2(n971), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(G1976), .B(KEYINPUT127), .ZN(n973) );
  XNOR2_X1 U1072 ( .A(n973), .B(G23), .ZN(n974) );
  NAND2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1074 ( .A(KEYINPUT58), .B(n976), .ZN(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1076 ( .A(KEYINPUT61), .B(n979), .ZN(n981) );
  INV_X1 U1077 ( .A(G16), .ZN(n980) );
  NAND2_X1 U1078 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1079 ( .A1(n982), .A2(G11), .ZN(n1040) );
  XNOR2_X1 U1080 ( .A(G301), .B(G1961), .ZN(n985) );
  XNOR2_X1 U1081 ( .A(n983), .B(G1348), .ZN(n984) );
  NOR2_X1 U1082 ( .A1(n985), .A2(n984), .ZN(n1004) );
  XNOR2_X1 U1083 ( .A(G299), .B(G1956), .ZN(n988) );
  INV_X1 U1084 ( .A(G1971), .ZN(n986) );
  NOR2_X1 U1085 ( .A1(n986), .A2(G166), .ZN(n987) );
  NOR2_X1 U1086 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1087 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1088 ( .A1(n992), .A2(n991), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1091 ( .A(KEYINPUT124), .B(n997), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G168), .ZN(n999) );
  NAND2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1094 ( .A(KEYINPUT57), .B(n1000), .Z(n1001) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(G1341), .B(n795), .ZN(n1005) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XOR2_X1 U1099 ( .A(G16), .B(KEYINPUT56), .Z(n1007) );
  NOR2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1101 ( .A(KEYINPUT125), .B(n1009), .ZN(n1038) );
  XNOR2_X1 U1102 ( .A(KEYINPUT119), .B(KEYINPUT52), .ZN(n1035) );
  XOR2_X1 U1103 ( .A(G160), .B(G2084), .Z(n1014) );
  NOR2_X1 U1104 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1105 ( .A(KEYINPUT117), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1106 ( .A1(n1014), .A2(n1013), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1109 ( .A(KEYINPUT118), .B(n1019), .ZN(n1033) );
  XOR2_X1 U1110 ( .A(G164), .B(G2078), .Z(n1023) );
  XNOR2_X1 U1111 ( .A(n1021), .B(n1020), .ZN(n1022) );
  NOR2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1113 ( .A(KEYINPUT50), .B(n1024), .Z(n1029) );
  XOR2_X1 U1114 ( .A(G2090), .B(G162), .Z(n1025) );
  NOR2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1116 ( .A(KEYINPUT51), .B(n1027), .ZN(n1028) );
  NOR2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1120 ( .A(n1035), .B(n1034), .ZN(n1036) );
  NAND2_X1 U1121 ( .A1(n1036), .A2(G29), .ZN(n1037) );
  NAND2_X1 U1122 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NOR2_X1 U1123 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NAND2_X1 U1124 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  XOR2_X1 U1125 ( .A(KEYINPUT62), .B(n1043), .Z(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

