//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT29), .ZN(new_n203));
  AND2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  INV_X1    g004(.A(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n204), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(G169gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(new_n206), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(KEYINPUT25), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(KEYINPUT24), .A3(new_n216), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n216), .A2(KEYINPUT24), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n222));
  OR2_X1    g021(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(new_n227), .B2(KEYINPUT23), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n221), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n217), .A2(new_n218), .ZN(new_n230));
  AND2_X1   g029(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n210), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n209), .A2(new_n233), .A3(KEYINPUT66), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n229), .A2(new_n230), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n220), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT27), .B(G183gat), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT67), .B1(new_n238), .B2(new_n214), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT69), .B1(new_n207), .B2(KEYINPUT26), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n207), .A2(KEYINPUT26), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT26), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n243), .A2(new_n226), .A3(new_n244), .A4(new_n247), .ZN(new_n248));
  OR2_X1    g047(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n250));
  AOI21_X1  g049(.A(G190gat), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n240), .B1(new_n251), .B2(KEYINPUT67), .ZN(new_n252));
  AND4_X1   g051(.A1(new_n216), .A2(new_n242), .A3(new_n248), .A4(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n203), .B1(new_n237), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G226gat), .ZN(new_n255));
  INV_X1    g054(.A(G233gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G211gat), .B(G218gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT74), .ZN(new_n261));
  XNOR2_X1  g060(.A(G197gat), .B(G204gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT22), .ZN(new_n263));
  INV_X1    g062(.A(G211gat), .ZN(new_n264));
  INV_X1    g063(.A(G218gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n260), .A2(KEYINPUT74), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n260), .A2(KEYINPUT74), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n269), .A2(new_n266), .A3(new_n262), .A4(new_n270), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n268), .A2(KEYINPUT75), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT75), .B1(new_n268), .B2(new_n271), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n257), .B1(new_n237), .B2(new_n253), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT85), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n259), .A2(KEYINPUT85), .A3(new_n274), .A4(new_n275), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n275), .A2(KEYINPUT76), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT76), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n282), .B(new_n257), .C1(new_n237), .C2(new_n253), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n281), .A2(new_n283), .B1(new_n258), .B2(new_n254), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(new_n274), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT37), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G8gat), .B(G36gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(G64gat), .B(G92gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n274), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n259), .A2(new_n291), .A3(new_n275), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n284), .B2(new_n291), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT37), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n290), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n286), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT87), .ZN(new_n299));
  OR2_X1    g098(.A1(KEYINPUT77), .A2(G155gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(KEYINPUT77), .A2(G155gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(G162gat), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT2), .ZN(new_n303));
  XNOR2_X1  g102(.A(G141gat), .B(G148gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G155gat), .B(G162gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n306), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(KEYINPUT2), .B2(new_n304), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n311));
  INV_X1    g110(.A(G113gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G120gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT72), .B(G120gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(new_n312), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316));
  XNOR2_X1  g115(.A(G127gat), .B(G134gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G120gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G113gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n313), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n321), .B1(new_n313), .B2(new_n320), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT1), .ZN(new_n324));
  NOR2_X1   g123(.A1(G127gat), .A2(G134gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT70), .B(G127gat), .ZN(new_n327));
  INV_X1    g126(.A(G134gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n318), .B1(new_n324), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n307), .A2(new_n331), .A3(new_n309), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n311), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n329), .ZN(new_n334));
  OR2_X1    g133(.A1(new_n322), .A2(new_n323), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(KEYINPUT1), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT2), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n306), .B1(new_n305), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n304), .B1(new_n302), .B2(KEYINPUT2), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n338), .B1(new_n306), .B2(new_n339), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n336), .A2(new_n340), .A3(KEYINPUT4), .A4(new_n318), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT4), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(new_n330), .B2(new_n310), .ZN(new_n343));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n333), .A2(new_n341), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n336), .A2(new_n340), .A3(new_n318), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n310), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n344), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT5), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n345), .B(new_n346), .C1(new_n351), .C2(new_n350), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n355));
  XNOR2_X1  g154(.A(G57gat), .B(G85gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n357), .B(new_n358), .Z(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n353), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(KEYINPUT84), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT84), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n353), .A2(new_n365), .A3(new_n354), .A4(new_n360), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n353), .A2(new_n354), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT6), .B1(new_n368), .B2(new_n359), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n363), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n293), .A2(new_n290), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT87), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n286), .A2(new_n295), .A3(new_n373), .A4(new_n297), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n299), .A2(new_n370), .A3(new_n372), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT88), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n295), .B1(new_n294), .B2(new_n293), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n296), .ZN(new_n378));
  AOI211_X1 g177(.A(new_n363), .B(new_n371), .C1(new_n367), .C2(new_n369), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT88), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n379), .A2(new_n380), .A3(new_n299), .A4(new_n374), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n376), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT89), .ZN(new_n383));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT31), .B(G50gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G22gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n268), .A2(new_n271), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n203), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n340), .B1(new_n390), .B2(new_n331), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G228gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(new_n256), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n332), .A2(new_n203), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n392), .B(new_n394), .C1(new_n274), .C2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n274), .A2(new_n395), .ZN(new_n397));
  OAI22_X1  g196(.A1(new_n397), .A2(new_n391), .B1(new_n393), .B2(new_n256), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n388), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OR2_X1    g198(.A1(new_n399), .A2(KEYINPUT82), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n396), .A2(new_n398), .A3(new_n388), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n387), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n401), .A2(KEYINPUT82), .ZN(new_n403));
  INV_X1    g202(.A(new_n401), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n387), .B1(new_n404), .B2(new_n399), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT81), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g206(.A(KEYINPUT81), .B(new_n387), .C1(new_n404), .C2(new_n399), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n402), .A2(new_n403), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT30), .B1(new_n293), .B2(new_n290), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n371), .B(new_n410), .Z(new_n411));
  NAND3_X1  g210(.A1(new_n333), .A2(new_n343), .A3(new_n341), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(KEYINPUT39), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n413), .A2(new_n344), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n348), .A2(new_n349), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(KEYINPUT39), .A3(new_n344), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n359), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(KEYINPUT40), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(KEYINPUT40), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n414), .A2(new_n359), .A3(new_n420), .A4(new_n416), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n419), .A2(new_n421), .B1(new_n364), .B2(new_n366), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n409), .B1(new_n411), .B2(new_n422), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n382), .A2(new_n383), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n383), .B1(new_n382), .B2(new_n423), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT73), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT36), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n237), .A2(new_n253), .ZN(new_n430));
  INV_X1    g229(.A(new_n330), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433));
  OR3_X1    g232(.A1(new_n432), .A2(KEYINPUT34), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n433), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT32), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT34), .B1(new_n432), .B2(new_n433), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n436), .B1(new_n434), .B2(new_n437), .ZN(new_n440));
  XNOR2_X1  g239(.A(G15gat), .B(G43gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(G71gat), .ZN(new_n442));
  INV_X1    g241(.A(G99gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n435), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(KEYINPUT33), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n439), .A2(new_n440), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n446), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n434), .A2(new_n437), .ZN(new_n449));
  INV_X1    g248(.A(new_n436), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n448), .B1(new_n451), .B2(new_n438), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n428), .B(new_n429), .C1(new_n447), .C2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n446), .B1(new_n439), .B2(new_n440), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n448), .A3(new_n438), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n454), .A2(new_n455), .A3(new_n426), .A4(new_n427), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n369), .A2(new_n361), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n458), .B(KEYINPUT80), .Z(new_n459));
  INV_X1    g258(.A(new_n363), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n411), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n409), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n457), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n424), .A2(new_n425), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT35), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n447), .A2(new_n452), .ZN(new_n466));
  INV_X1    g265(.A(new_n411), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n462), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n465), .B1(new_n468), .B2(new_n370), .ZN(new_n469));
  INV_X1    g268(.A(new_n466), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(new_n409), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(KEYINPUT35), .A3(new_n461), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n202), .B1(new_n464), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n382), .A2(new_n423), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT89), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n461), .A2(new_n462), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n453), .A2(new_n456), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n382), .A2(new_n383), .A3(new_n423), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n476), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n469), .A2(new_n472), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(KEYINPUT90), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n474), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT16), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n485), .B1(new_n486), .B2(G1gat), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(G1gat), .B2(new_n485), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(G8gat), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT14), .ZN(new_n490));
  INV_X1    g289(.A(G29gat), .ZN(new_n491));
  INV_X1    g290(.A(G36gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n493), .A2(new_n494), .B1(G29gat), .B2(G36gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(G43gat), .B(G50gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(KEYINPUT15), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(KEYINPUT15), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n497), .B(new_n498), .Z(new_n499));
  INV_X1    g298(.A(KEYINPUT91), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT17), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n497), .B(new_n498), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT91), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n503), .A2(new_n502), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n489), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n501), .A2(new_n504), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n509), .A2(new_n489), .ZN(new_n510));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n508), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT92), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT18), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT18), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n509), .A2(new_n489), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n503), .B(new_n500), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n506), .B1(new_n518), .B2(new_n502), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n517), .B1(new_n519), .B2(new_n489), .ZN(new_n520));
  OAI211_X1 g319(.A(KEYINPUT92), .B(new_n516), .C1(new_n520), .C2(new_n512), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n509), .B(new_n489), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n511), .B(KEYINPUT13), .Z(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n515), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  INV_X1    g325(.A(G197gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT11), .B(G169gat), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n528), .B(new_n529), .Z(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT12), .Z(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n515), .A2(new_n521), .A3(new_n531), .A4(new_n524), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(KEYINPUT93), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT93), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n525), .A2(new_n536), .A3(new_n532), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT98), .ZN(new_n539));
  NAND2_X1  g338(.A1(G85gat), .A2(G92gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  INV_X1    g340(.A(G106gat), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT8), .B1(new_n443), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n541), .B(new_n543), .C1(G85gat), .C2(G92gat), .ZN(new_n544));
  XOR2_X1   g343(.A(G99gat), .B(G106gat), .Z(new_n545));
  OR2_X1    g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n545), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n519), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n509), .A2(new_n549), .ZN(new_n551));
  NAND3_X1  g350(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(G190gat), .B(G218gat), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n551), .B(new_n552), .C1(new_n519), .C2(new_n549), .ZN(new_n555));
  INV_X1    g354(.A(new_n553), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT97), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n539), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n554), .A2(KEYINPUT98), .A3(new_n557), .ZN(new_n561));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n564), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n539), .B(new_n566), .C1(new_n558), .C2(new_n559), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT94), .ZN(new_n570));
  INV_X1    g369(.A(G64gat), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n570), .B1(new_n571), .B2(G57gat), .ZN(new_n572));
  INV_X1    g371(.A(G57gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(KEYINPUT94), .A3(G64gat), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n572), .B(new_n574), .C1(new_n573), .C2(G64gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(G71gat), .B(G78gat), .ZN(new_n576));
  AND2_X1   g375(.A1(G71gat), .A2(G78gat), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n575), .B(new_n576), .C1(KEYINPUT9), .C2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT95), .ZN(new_n579));
  INV_X1    g378(.A(new_n576), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581));
  XNOR2_X1  g380(.A(G57gat), .B(G64gat), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT21), .ZN(new_n585));
  XOR2_X1   g384(.A(KEYINPUT96), .B(G211gat), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n587), .A2(new_n588), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n489), .B1(new_n584), .B2(KEYINPUT21), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(new_n213), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(G127gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n592), .B(G183gat), .ZN(new_n595));
  INV_X1    g394(.A(G127gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n594), .B(new_n597), .C1(new_n589), .C2(new_n590), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G155gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n599), .A2(new_n600), .A3(new_n603), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n569), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(G230gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(new_n256), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT100), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n546), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n547), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n544), .A2(new_n612), .A3(new_n545), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n584), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n584), .A2(KEYINPUT99), .A3(new_n549), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT99), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n579), .A2(new_n583), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n618), .B1(new_n619), .B2(new_n548), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n611), .B(new_n616), .C1(new_n617), .C2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n584), .A2(KEYINPUT10), .A3(new_n549), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n610), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n616), .B1(new_n617), .B2(new_n620), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n610), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n484), .A2(new_n538), .A3(new_n608), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n459), .A2(new_n460), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT101), .B(G1gat), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(G1324gat));
  NOR2_X1   g438(.A1(new_n635), .A2(new_n467), .ZN(new_n640));
  INV_X1    g439(.A(G8gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n486), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n486), .A2(new_n641), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n640), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n647), .B(new_n648), .C1(new_n641), .C2(new_n640), .ZN(G1325gat));
  INV_X1    g448(.A(new_n635), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n478), .B(KEYINPUT102), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n650), .A2(G15gat), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(G15gat), .B1(new_n650), .B2(new_n466), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(G1326gat));
  NAND3_X1  g454(.A1(new_n650), .A2(new_n388), .A3(new_n409), .ZN(new_n656));
  OAI21_X1  g455(.A(G22gat), .B1(new_n635), .B2(new_n462), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  NAND2_X1  g459(.A1(new_n481), .A2(new_n482), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n568), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n565), .A2(KEYINPUT104), .A3(new_n567), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n661), .A2(new_n662), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n568), .B1(new_n474), .B2(new_n483), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n668), .B1(new_n669), .B2(new_n662), .ZN(new_n670));
  INV_X1    g469(.A(new_n636), .ZN(new_n671));
  INV_X1    g470(.A(new_n606), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n603), .B1(new_n599), .B2(new_n600), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n535), .A2(new_n537), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n674), .A2(new_n675), .A3(new_n633), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n670), .A2(new_n671), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(G29gat), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n669), .A2(new_n676), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n491), .A3(new_n671), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT45), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(new_n685), .ZN(G1328gat));
  NAND3_X1  g485(.A1(new_n683), .A2(new_n492), .A3(new_n411), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n687), .A2(KEYINPUT46), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(KEYINPUT46), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n662), .B1(new_n484), .B2(new_n569), .ZN(new_n690));
  INV_X1    g489(.A(new_n668), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n676), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n692), .A2(new_n467), .A3(new_n693), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n688), .B(new_n689), .C1(new_n492), .C2(new_n694), .ZN(G1329gat));
  NOR2_X1   g494(.A1(new_n682), .A2(G43gat), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n466), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n692), .A2(new_n457), .A3(new_n693), .ZN(new_n698));
  INV_X1    g497(.A(G43gat), .ZN(new_n699));
  OAI211_X1 g498(.A(KEYINPUT47), .B(new_n697), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n670), .A2(new_n652), .A3(new_n676), .ZN(new_n701));
  AOI22_X1  g500(.A1(new_n701), .A2(G43gat), .B1(new_n696), .B2(new_n466), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(KEYINPUT47), .B2(new_n702), .ZN(G1330gat));
  NAND4_X1  g502(.A1(new_n670), .A2(G50gat), .A3(new_n409), .A4(new_n676), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n682), .A2(new_n462), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(G50gat), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g506(.A1(new_n661), .A2(new_n675), .A3(new_n608), .A4(new_n633), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n636), .B(KEYINPUT106), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(new_n573), .ZN(G1332gat));
  NOR2_X1   g510(.A1(new_n708), .A2(new_n467), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT49), .B(G64gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n712), .B2(new_n715), .ZN(G1333gat));
  OAI21_X1  g515(.A(G71gat), .B1(new_n708), .B2(new_n651), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n708), .A2(G71gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(new_n470), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g519(.A1(new_n708), .A2(new_n462), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g521(.A1(new_n607), .A2(new_n675), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n481), .B2(new_n482), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n569), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(KEYINPUT51), .A3(new_n569), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n634), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(G85gat), .B1(new_n729), .B2(new_n671), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n723), .A2(new_n634), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n481), .A2(KEYINPUT90), .A3(new_n482), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT90), .B1(new_n481), .B2(new_n482), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n569), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT44), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n732), .B1(new_n736), .B2(new_n668), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n671), .A2(G85gat), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n730), .B1(new_n737), .B2(new_n738), .ZN(G1336gat));
  OAI211_X1 g538(.A(new_n411), .B(new_n731), .C1(new_n690), .C2(new_n691), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n670), .A2(KEYINPUT108), .A3(new_n411), .A4(new_n731), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(G92gat), .A3(new_n743), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n724), .A2(KEYINPUT51), .A3(new_n569), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT51), .B1(new_n724), .B2(new_n569), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n634), .A2(G92gat), .A3(new_n467), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT52), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n744), .A2(new_n750), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n740), .A2(G92gat), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n749), .B(KEYINPUT107), .Z(new_n753));
  NOR2_X1   g552(.A1(new_n747), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT52), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n751), .A2(new_n755), .ZN(G1337gat));
  AOI21_X1  g555(.A(G99gat), .B1(new_n729), .B2(new_n466), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n651), .A2(new_n443), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n757), .B1(new_n737), .B2(new_n758), .ZN(G1338gat));
  OAI211_X1 g558(.A(new_n409), .B(new_n731), .C1(new_n690), .C2(new_n691), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT111), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT109), .B(G106gat), .Z(new_n762));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n670), .A2(new_n763), .A3(new_n409), .A4(new_n731), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n542), .B(new_n633), .C1(new_n745), .C2(new_n746), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n462), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(KEYINPUT53), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT110), .B1(new_n766), .B2(new_n462), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n729), .A2(new_n771), .A3(new_n542), .A4(new_n409), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n762), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n737), .B2(new_n409), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT53), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n769), .A2(new_n776), .ZN(G1339gat));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n778));
  INV_X1    g577(.A(new_n530), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n520), .A2(new_n512), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n522), .A2(new_n523), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n782), .A2(KEYINPUT114), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(KEYINPUT114), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n783), .A2(new_n534), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n633), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n621), .A2(new_n610), .A3(new_n622), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n624), .A2(KEYINPUT54), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n623), .A2(new_n789), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n790), .A2(KEYINPUT113), .A3(new_n630), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT113), .B1(new_n790), .B2(new_n630), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n788), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(KEYINPUT55), .B(new_n788), .C1(new_n791), .C2(new_n792), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n631), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n786), .B1(new_n797), .B2(new_n675), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n666), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n785), .A2(new_n795), .A3(new_n631), .A4(new_n796), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n666), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n674), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n674), .A2(new_n634), .A3(new_n568), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT112), .B1(new_n803), .B2(new_n538), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n608), .A2(new_n805), .A3(new_n675), .A4(new_n634), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n778), .B1(new_n808), .B2(new_n409), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n636), .A2(new_n411), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n804), .A2(new_n806), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n666), .A2(new_n800), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n666), .B2(new_n798), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n813), .B2(new_n674), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(KEYINPUT115), .A3(new_n462), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n809), .A2(new_n466), .A3(new_n810), .A4(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(G113gat), .B1(new_n816), .B2(new_n675), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n808), .A2(new_n468), .A3(new_n709), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n312), .A3(new_n538), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(G1340gat));
  OAI21_X1  g619(.A(G120gat), .B1(new_n816), .B2(new_n634), .ZN(new_n821));
  INV_X1    g620(.A(new_n314), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n818), .A2(new_n822), .A3(new_n633), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1341gat));
  NOR3_X1   g623(.A1(new_n816), .A2(new_n327), .A3(new_n607), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n818), .A2(new_n674), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n327), .B2(new_n826), .ZN(G1342gat));
  NAND3_X1  g626(.A1(new_n818), .A2(new_n328), .A3(new_n569), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n828), .A2(KEYINPUT56), .ZN(new_n829));
  OAI21_X1  g628(.A(G134gat), .B1(new_n816), .B2(new_n568), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(KEYINPUT56), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(G1343gat));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n833), .B(new_n409), .C1(new_n802), .C2(new_n807), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n478), .A2(new_n636), .A3(new_n411), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n538), .A2(new_n631), .A3(new_n796), .A4(new_n795), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n569), .B1(new_n836), .B2(new_n786), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n607), .B1(new_n837), .B2(new_n812), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n462), .B1(new_n838), .B2(new_n811), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n834), .B(new_n835), .C1(new_n833), .C2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G141gat), .B1(new_n840), .B2(new_n675), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT58), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n651), .A2(new_n409), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n808), .A2(new_n709), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(G141gat), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n846), .A2(new_n847), .A3(new_n467), .A4(new_n538), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n841), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n841), .B2(new_n848), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n844), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n841), .A2(new_n848), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT117), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n841), .B2(new_n842), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n848), .A3(new_n849), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n852), .A2(new_n858), .ZN(G1344gat));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT57), .B1(new_n808), .B2(new_n462), .ZN(new_n861));
  INV_X1    g660(.A(new_n837), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n800), .A2(new_n568), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n674), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n803), .A2(new_n538), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n833), .B(new_n409), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n861), .A2(new_n633), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n835), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n860), .B1(new_n869), .B2(G148gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n860), .B1(new_n840), .B2(new_n634), .ZN(new_n871));
  INV_X1    g670(.A(G148gat), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n846), .A2(new_n467), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n633), .A2(new_n872), .ZN(new_n875));
  OAI22_X1  g674(.A1(new_n870), .A2(new_n873), .B1(new_n874), .B2(new_n875), .ZN(G1345gat));
  NAND2_X1  g675(.A1(new_n300), .A2(new_n301), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n840), .A2(new_n877), .A3(new_n607), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n846), .A2(new_n467), .A3(new_n674), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n877), .B2(new_n879), .ZN(G1346gat));
  OAI21_X1  g679(.A(G162gat), .B1(new_n840), .B2(new_n666), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n874), .A2(G162gat), .A3(new_n568), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(G1347gat));
  NAND4_X1  g685(.A1(new_n814), .A2(new_n636), .A3(new_n471), .A4(new_n411), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n205), .B1(new_n887), .B2(new_n675), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889));
  INV_X1    g688(.A(new_n709), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n467), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n709), .A2(KEYINPUT119), .A3(new_n411), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n809), .A2(new_n466), .A3(new_n815), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n538), .A2(G169gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n888), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT120), .ZN(G1348gat));
  INV_X1    g696(.A(new_n887), .ZN(new_n898));
  AOI21_X1  g697(.A(G176gat), .B1(new_n898), .B2(new_n633), .ZN(new_n899));
  INV_X1    g698(.A(new_n894), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n634), .A2(new_n232), .A3(new_n231), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(G1349gat));
  OAI21_X1  g701(.A(G183gat), .B1(new_n894), .B2(new_n607), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n898), .A2(new_n238), .A3(new_n674), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g705(.A(G190gat), .B1(new_n894), .B2(new_n568), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n898), .A2(new_n214), .A3(new_n667), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT121), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n907), .A2(new_n908), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n909), .A2(new_n911), .A3(new_n912), .ZN(G1351gat));
  NOR2_X1   g712(.A1(new_n845), .A2(new_n467), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n814), .A2(new_n916), .A3(new_n636), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n914), .A2(new_n915), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT123), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n921), .B1(new_n917), .B2(new_n918), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n920), .A2(new_n922), .A3(new_n527), .A4(new_n538), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n891), .A2(new_n651), .A3(new_n892), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n924), .B(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n861), .A3(new_n866), .ZN(new_n927));
  OAI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n675), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n923), .A2(new_n928), .A3(KEYINPUT125), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1352gat));
  NAND2_X1  g732(.A1(new_n868), .A2(new_n926), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT126), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n868), .A2(new_n936), .A3(new_n926), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(G204gat), .A3(new_n937), .ZN(new_n938));
  NOR4_X1   g737(.A1(new_n917), .A2(G204gat), .A3(new_n634), .A4(new_n918), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT62), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1353gat));
  NAND4_X1  g740(.A1(new_n926), .A2(new_n674), .A3(new_n861), .A4(new_n866), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(G211gat), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT63), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n920), .A2(new_n922), .A3(new_n264), .A4(new_n674), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n944), .A2(KEYINPUT63), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n944), .A2(KEYINPUT63), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n942), .A2(G211gat), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(G1354gat));
  NOR3_X1   g749(.A1(new_n927), .A2(new_n265), .A3(new_n568), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n920), .A2(new_n922), .A3(new_n667), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n951), .B1(new_n265), .B2(new_n952), .ZN(G1355gat));
endmodule


