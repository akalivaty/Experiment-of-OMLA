

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U319 ( .A(n295), .B(n373), .ZN(n296) );
  INV_X1 U320 ( .A(KEYINPUT77), .ZN(n301) );
  XNOR2_X1 U321 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n443) );
  AND2_X1 U322 ( .A1(G232GAT), .A2(G233GAT), .ZN(n287) );
  XOR2_X1 U323 ( .A(n404), .B(n403), .Z(n288) );
  XNOR2_X1 U324 ( .A(n405), .B(n287), .ZN(n295) );
  XNOR2_X1 U325 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n403) );
  XNOR2_X1 U326 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U327 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U328 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U329 ( .A(KEYINPUT93), .B(n457), .ZN(n509) );
  XNOR2_X1 U330 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n446) );
  XNOR2_X1 U331 ( .A(n447), .B(n446), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n290) );
  XNOR2_X1 U333 ( .A(G162GAT), .B(KEYINPUT9), .ZN(n289) );
  XNOR2_X1 U334 ( .A(n290), .B(n289), .ZN(n306) );
  XOR2_X1 U335 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n292) );
  XOR2_X1 U336 ( .A(G50GAT), .B(KEYINPUT74), .Z(n433) );
  XOR2_X1 U337 ( .A(G36GAT), .B(G190GAT), .Z(n390) );
  XNOR2_X1 U338 ( .A(n433), .B(n390), .ZN(n291) );
  XNOR2_X1 U339 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U340 ( .A(n293), .B(KEYINPUT10), .Z(n298) );
  XOR2_X1 U341 ( .A(G29GAT), .B(G134GAT), .Z(n405) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n294), .B(KEYINPUT8), .ZN(n373) );
  XNOR2_X1 U344 ( .A(G218GAT), .B(n296), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n304) );
  XOR2_X1 U346 ( .A(KEYINPUT71), .B(G92GAT), .Z(n300) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G85GAT), .ZN(n299) );
  XNOR2_X1 U348 ( .A(n300), .B(n299), .ZN(n347) );
  XNOR2_X1 U349 ( .A(G106GAT), .B(n347), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n534) );
  XOR2_X1 U351 ( .A(KEYINPUT64), .B(KEYINPUT84), .Z(n308) );
  XNOR2_X1 U352 ( .A(KEYINPUT20), .B(KEYINPUT82), .ZN(n307) );
  XNOR2_X1 U353 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U354 ( .A(G176GAT), .B(G190GAT), .Z(n310) );
  XNOR2_X1 U355 ( .A(G43GAT), .B(G15GAT), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U357 ( .A(n312), .B(n311), .ZN(n327) );
  XOR2_X1 U358 ( .A(G127GAT), .B(KEYINPUT81), .Z(n314) );
  XNOR2_X1 U359 ( .A(KEYINPUT0), .B(KEYINPUT80), .ZN(n313) );
  XNOR2_X1 U360 ( .A(n314), .B(n313), .ZN(n407) );
  XOR2_X1 U361 ( .A(G134GAT), .B(n407), .Z(n316) );
  NAND2_X1 U362 ( .A1(G227GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U364 ( .A(n317), .B(G99GAT), .Z(n325) );
  XOR2_X1 U365 ( .A(KEYINPUT83), .B(KEYINPUT17), .Z(n319) );
  XNOR2_X1 U366 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U368 ( .A(G169GAT), .B(n320), .Z(n400) );
  XOR2_X1 U369 ( .A(G71GAT), .B(G120GAT), .Z(n322) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(G183GAT), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n400), .B(n323), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U374 ( .A(n327), .B(n326), .ZN(n525) );
  XNOR2_X1 U375 ( .A(KEYINPUT36), .B(KEYINPUT102), .ZN(n328) );
  XNOR2_X1 U376 ( .A(n534), .B(n328), .ZN(n478) );
  XOR2_X1 U377 ( .A(G57GAT), .B(G78GAT), .Z(n330) );
  XNOR2_X1 U378 ( .A(G1GAT), .B(G127GAT), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n330), .B(n329), .ZN(n344) );
  XOR2_X1 U380 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n332) );
  XNOR2_X1 U381 ( .A(G64GAT), .B(KEYINPUT79), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U383 ( .A(G8GAT), .B(G183GAT), .Z(n387) );
  XOR2_X1 U384 ( .A(n387), .B(G211GAT), .Z(n334) );
  XOR2_X1 U385 ( .A(G22GAT), .B(G15GAT), .Z(n371) );
  XNOR2_X1 U386 ( .A(n371), .B(G155GAT), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U388 ( .A(n336), .B(n335), .Z(n338) );
  NAND2_X1 U389 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U390 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U391 ( .A(n339), .B(KEYINPUT78), .Z(n342) );
  XNOR2_X1 U392 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n340), .B(KEYINPUT70), .ZN(n348) );
  XNOR2_X1 U394 ( .A(n348), .B(KEYINPUT12), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U396 ( .A(n344), .B(n343), .Z(n559) );
  NAND2_X1 U397 ( .A1(n478), .A2(n559), .ZN(n346) );
  XNOR2_X1 U398 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n346), .B(n345), .ZN(n377) );
  XOR2_X1 U400 ( .A(n348), .B(n347), .Z(n352) );
  XNOR2_X1 U401 ( .A(G106GAT), .B(G78GAT), .ZN(n349) );
  XNOR2_X1 U402 ( .A(n349), .B(G204GAT), .ZN(n432) );
  XNOR2_X1 U403 ( .A(G120GAT), .B(G148GAT), .ZN(n350) );
  XNOR2_X1 U404 ( .A(n350), .B(G57GAT), .ZN(n406) );
  XNOR2_X1 U405 ( .A(n432), .B(n406), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n359) );
  XOR2_X1 U407 ( .A(G176GAT), .B(G64GAT), .Z(n386) );
  XOR2_X1 U408 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n354) );
  XNOR2_X1 U409 ( .A(KEYINPUT32), .B(KEYINPUT72), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U411 ( .A(n386), .B(n355), .Z(n357) );
  NAND2_X1 U412 ( .A1(G230GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n359), .B(n358), .ZN(n448) );
  XOR2_X1 U415 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n361) );
  NAND2_X1 U416 ( .A1(G229GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U418 ( .A(n362), .B(KEYINPUT29), .Z(n370) );
  XOR2_X1 U419 ( .A(G141GAT), .B(G36GAT), .Z(n364) );
  XNOR2_X1 U420 ( .A(G29GAT), .B(G50GAT), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U422 ( .A(KEYINPUT30), .B(G8GAT), .Z(n366) );
  XNOR2_X1 U423 ( .A(G169GAT), .B(G197GAT), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n372) );
  XOR2_X1 U427 ( .A(n372), .B(n371), .Z(n375) );
  XOR2_X1 U428 ( .A(G113GAT), .B(G1GAT), .Z(n411) );
  XNOR2_X1 U429 ( .A(n373), .B(n411), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n566) );
  INV_X1 U431 ( .A(n566), .ZN(n552) );
  NOR2_X1 U432 ( .A1(n448), .A2(n552), .ZN(n376) );
  NAND2_X1 U433 ( .A1(n377), .A2(n376), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n378), .B(KEYINPUT112), .ZN(n384) );
  INV_X1 U435 ( .A(n534), .ZN(n550) );
  INV_X1 U436 ( .A(n559), .ZN(n575) );
  NAND2_X1 U437 ( .A1(n550), .A2(n575), .ZN(n381) );
  XOR2_X1 U438 ( .A(KEYINPUT41), .B(n448), .Z(n554) );
  INV_X1 U439 ( .A(n554), .ZN(n544) );
  NOR2_X1 U440 ( .A1(n566), .A2(n544), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n379), .B(KEYINPUT46), .ZN(n380) );
  NOR2_X1 U442 ( .A1(n381), .A2(n380), .ZN(n382) );
  XNOR2_X1 U443 ( .A(KEYINPUT47), .B(n382), .ZN(n383) );
  NAND2_X1 U444 ( .A1(n384), .A2(n383), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n385), .B(KEYINPUT48), .ZN(n520) );
  XOR2_X1 U446 ( .A(n387), .B(n386), .Z(n389) );
  NAND2_X1 U447 ( .A1(G226GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n391) );
  XOR2_X1 U449 ( .A(n391), .B(n390), .Z(n399) );
  XOR2_X1 U450 ( .A(KEYINPUT87), .B(G218GAT), .Z(n393) );
  XNOR2_X1 U451 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U453 ( .A(G197GAT), .B(n394), .Z(n437) );
  XOR2_X1 U454 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n396) );
  XNOR2_X1 U455 ( .A(G204GAT), .B(G92GAT), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n437), .B(n397), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n402) );
  INV_X1 U459 ( .A(n400), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n511) );
  NAND2_X1 U461 ( .A1(n520), .A2(n511), .ZN(n404) );
  XOR2_X1 U462 ( .A(n406), .B(n405), .Z(n413) );
  XOR2_X1 U463 ( .A(n407), .B(KEYINPUT4), .Z(n409) );
  NAND2_X1 U464 ( .A1(G225GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U468 ( .A(KEYINPUT89), .B(KEYINPUT6), .Z(n415) );
  XNOR2_X1 U469 ( .A(G85GAT), .B(KEYINPUT92), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U471 ( .A(n417), .B(n416), .Z(n425) );
  XOR2_X1 U472 ( .A(KEYINPUT3), .B(G162GAT), .Z(n419) );
  XNOR2_X1 U473 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U475 ( .A(G141GAT), .B(n420), .Z(n441) );
  XOR2_X1 U476 ( .A(KEYINPUT1), .B(KEYINPUT90), .Z(n422) );
  XNOR2_X1 U477 ( .A(KEYINPUT5), .B(KEYINPUT91), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n441), .B(n423), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n457) );
  INV_X1 U481 ( .A(n509), .ZN(n563) );
  XOR2_X1 U482 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n427) );
  XNOR2_X1 U483 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U485 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n429) );
  XNOR2_X1 U486 ( .A(G22GAT), .B(G148GAT), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U488 ( .A(n431), .B(n430), .Z(n439) );
  XOR2_X1 U489 ( .A(n433), .B(n432), .Z(n435) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n460) );
  AND2_X1 U495 ( .A1(n563), .A2(n460), .ZN(n442) );
  NAND2_X1 U496 ( .A1(n288), .A2(n442), .ZN(n444) );
  NOR2_X1 U497 ( .A1(n525), .A2(n445), .ZN(n560) );
  NAND2_X1 U498 ( .A1(n534), .A2(n560), .ZN(n447) );
  INV_X1 U499 ( .A(n448), .ZN(n570) );
  NAND2_X1 U500 ( .A1(n552), .A2(n570), .ZN(n449) );
  XOR2_X1 U501 ( .A(n449), .B(KEYINPUT73), .Z(n483) );
  NOR2_X1 U502 ( .A1(n534), .A2(n575), .ZN(n450) );
  XNOR2_X1 U503 ( .A(n450), .B(KEYINPUT16), .ZN(n465) );
  INV_X1 U504 ( .A(n525), .ZN(n514) );
  NAND2_X1 U505 ( .A1(n511), .A2(n514), .ZN(n451) );
  NAND2_X1 U506 ( .A1(n460), .A2(n451), .ZN(n452) );
  XOR2_X1 U507 ( .A(KEYINPUT25), .B(n452), .Z(n455) );
  NOR2_X1 U508 ( .A1(n460), .A2(n514), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n453), .B(KEYINPUT26), .ZN(n564) );
  XNOR2_X1 U510 ( .A(n511), .B(KEYINPUT27), .ZN(n461) );
  NAND2_X1 U511 ( .A1(n564), .A2(n461), .ZN(n454) );
  NAND2_X1 U512 ( .A1(n455), .A2(n454), .ZN(n456) );
  XNOR2_X1 U513 ( .A(KEYINPUT96), .B(n456), .ZN(n458) );
  NAND2_X1 U514 ( .A1(n458), .A2(n457), .ZN(n464) );
  XOR2_X1 U515 ( .A(KEYINPUT28), .B(KEYINPUT67), .Z(n459) );
  XNOR2_X1 U516 ( .A(n460), .B(n459), .ZN(n523) );
  NAND2_X1 U517 ( .A1(n509), .A2(n461), .ZN(n521) );
  NOR2_X1 U518 ( .A1(n514), .A2(n521), .ZN(n462) );
  NAND2_X1 U519 ( .A1(n523), .A2(n462), .ZN(n463) );
  NAND2_X1 U520 ( .A1(n464), .A2(n463), .ZN(n479) );
  NAND2_X1 U521 ( .A1(n465), .A2(n479), .ZN(n495) );
  NOR2_X1 U522 ( .A1(n483), .A2(n495), .ZN(n475) );
  NAND2_X1 U523 ( .A1(n509), .A2(n475), .ZN(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT98), .B(KEYINPUT34), .Z(n467) );
  XNOR2_X1 U525 ( .A(G1GAT), .B(KEYINPUT97), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(G1324GAT) );
  XOR2_X1 U528 ( .A(G8GAT), .B(KEYINPUT99), .Z(n471) );
  NAND2_X1 U529 ( .A1(n475), .A2(n511), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n471), .B(n470), .ZN(G1325GAT) );
  XOR2_X1 U531 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n473) );
  NAND2_X1 U532 ( .A1(n475), .A2(n514), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U534 ( .A(G15GAT), .B(n474), .ZN(G1326GAT) );
  XOR2_X1 U535 ( .A(G22GAT), .B(KEYINPUT101), .Z(n477) );
  INV_X1 U536 ( .A(n523), .ZN(n517) );
  NAND2_X1 U537 ( .A1(n475), .A2(n517), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(G1327GAT) );
  XOR2_X1 U539 ( .A(G29GAT), .B(KEYINPUT39), .Z(n486) );
  NAND2_X1 U540 ( .A1(n478), .A2(n479), .ZN(n480) );
  NOR2_X1 U541 ( .A1(n559), .A2(n480), .ZN(n482) );
  XNOR2_X1 U542 ( .A(KEYINPUT37), .B(KEYINPUT103), .ZN(n481) );
  XOR2_X1 U543 ( .A(n482), .B(n481), .Z(n508) );
  OR2_X1 U544 ( .A1(n483), .A2(n508), .ZN(n484) );
  XOR2_X1 U545 ( .A(KEYINPUT38), .B(n484), .Z(n493) );
  NAND2_X1 U546 ( .A1(n493), .A2(n509), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(G1328GAT) );
  NAND2_X1 U548 ( .A1(n493), .A2(n511), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n487), .B(KEYINPUT104), .ZN(n488) );
  XNOR2_X1 U550 ( .A(G36GAT), .B(n488), .ZN(G1329GAT) );
  XNOR2_X1 U551 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n492) );
  XOR2_X1 U552 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n490) );
  NAND2_X1 U553 ( .A1(n493), .A2(n514), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(G1330GAT) );
  NAND2_X1 U556 ( .A1(n517), .A2(n493), .ZN(n494) );
  XNOR2_X1 U557 ( .A(G50GAT), .B(n494), .ZN(G1331GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n497) );
  NAND2_X1 U559 ( .A1(n554), .A2(n566), .ZN(n507) );
  NOR2_X1 U560 ( .A1(n507), .A2(n495), .ZN(n504) );
  NAND2_X1 U561 ( .A1(n504), .A2(n509), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(n498), .ZN(G1332GAT) );
  NAND2_X1 U564 ( .A1(n504), .A2(n511), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n499), .B(KEYINPUT108), .ZN(n500) );
  XNOR2_X1 U566 ( .A(G64GAT), .B(n500), .ZN(G1333GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n502) );
  NAND2_X1 U568 ( .A1(n504), .A2(n514), .ZN(n501) );
  XNOR2_X1 U569 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(n503), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .Z(n506) );
  NAND2_X1 U572 ( .A1(n504), .A2(n517), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(G1335GAT) );
  NOR2_X1 U574 ( .A1(n508), .A2(n507), .ZN(n516) );
  NAND2_X1 U575 ( .A1(n516), .A2(n509), .ZN(n510) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(n510), .ZN(G1336GAT) );
  XOR2_X1 U577 ( .A(G92GAT), .B(KEYINPUT111), .Z(n513) );
  NAND2_X1 U578 ( .A1(n516), .A2(n511), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(G1337GAT) );
  NAND2_X1 U580 ( .A1(n514), .A2(n516), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n515), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n518), .B(KEYINPUT44), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  INV_X1 U585 ( .A(n520), .ZN(n522) );
  NOR2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n539) );
  NAND2_X1 U587 ( .A1(n523), .A2(n539), .ZN(n524) );
  NOR2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n535), .A2(n552), .ZN(n526) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U592 ( .A1(n535), .A2(n554), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n530) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(KEYINPUT114), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U597 ( .A(KEYINPUT113), .B(n531), .Z(n533) );
  NAND2_X1 U598 ( .A1(n535), .A2(n559), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n537) );
  NAND2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n539), .A2(n564), .ZN(n549) );
  NOR2_X1 U605 ( .A1(n566), .A2(n549), .ZN(n541) );
  XNOR2_X1 U606 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n543) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n546) );
  NOR2_X1 U611 ( .A1(n544), .A2(n549), .ZN(n545) );
  XOR2_X1 U612 ( .A(n546), .B(n545), .Z(G1345GAT) );
  NOR2_X1 U613 ( .A1(n575), .A2(n549), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1346GAT) );
  NOR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U617 ( .A(G162GAT), .B(n551), .Z(G1347GAT) );
  NAND2_X1 U618 ( .A1(n560), .A2(n552), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G169GAT), .B(n553), .ZN(G1348GAT) );
  XNOR2_X1 U620 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n558) );
  NAND2_X1 U621 ( .A1(n560), .A2(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT56), .Z(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1349GAT) );
  XOR2_X1 U625 ( .A(G183GAT), .B(KEYINPUT123), .Z(n562) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1350GAT) );
  AND2_X1 U628 ( .A1(n563), .A2(n288), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n565), .A2(n564), .ZN(n577) );
  NOR2_X1 U630 ( .A1(n566), .A2(n577), .ZN(n568) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U634 ( .A1(n577), .A2(n570), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U639 ( .A1(n575), .A2(n577), .ZN(n576) );
  XOR2_X1 U640 ( .A(G211GAT), .B(n576), .Z(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n580) );
  INV_X1 U642 ( .A(n577), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n578), .A2(n478), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(G218GAT), .B(n581), .Z(G1355GAT) );
endmodule

