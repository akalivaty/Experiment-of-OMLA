

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U551 ( .A1(n525), .A2(G2105), .ZN(n887) );
  AND2_X2 U552 ( .A1(G138), .A2(n549), .ZN(n518) );
  AND2_X2 U553 ( .A1(G2104), .A2(G2105), .ZN(n547) );
  NAND2_X2 U554 ( .A1(G8), .A2(n709), .ZN(n778) );
  OR2_X1 U555 ( .A1(n700), .A2(n699), .ZN(n723) );
  AND2_X1 U556 ( .A1(n725), .A2(G2072), .ZN(n693) );
  NAND2_X1 U557 ( .A1(n690), .A2(n781), .ZN(n709) );
  AND2_X1 U558 ( .A1(n781), .A2(n690), .ZN(n725) );
  NOR2_X1 U559 ( .A1(G1384), .A2(G164), .ZN(n689) );
  XNOR2_X1 U560 ( .A(n552), .B(KEYINPUT91), .ZN(G164) );
  NOR2_X1 U561 ( .A1(n550), .A2(n518), .ZN(n551) );
  NOR2_X2 U562 ( .A1(G2105), .A2(n525), .ZN(n891) );
  XOR2_X2 U563 ( .A(KEYINPUT0), .B(G543), .Z(n538) );
  NOR2_X1 U564 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  OR2_X2 U565 ( .A1(n771), .A2(n770), .ZN(n522) );
  BUF_X1 U566 ( .A(n549), .Z(n517) );
  NOR2_X1 U567 ( .A1(n698), .A2(n979), .ZN(n697) );
  XNOR2_X1 U568 ( .A(n693), .B(n692), .ZN(n694) );
  NAND2_X1 U569 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U570 ( .A(n708), .B(n707), .ZN(n713) );
  AND2_X1 U571 ( .A1(n978), .A2(n716), .ZN(n706) );
  INV_X1 U572 ( .A(KEYINPUT105), .ZN(n739) );
  XNOR2_X1 U573 ( .A(n724), .B(KEYINPUT29), .ZN(n749) );
  NAND2_X1 U574 ( .A1(n723), .A2(n722), .ZN(n724) );
  AND2_X1 U575 ( .A1(n546), .A2(n545), .ZN(n519) );
  AND2_X1 U576 ( .A1(n780), .A2(n779), .ZN(n520) );
  OR2_X1 U577 ( .A1(n769), .A2(n778), .ZN(n521) );
  AND2_X1 U578 ( .A1(n988), .A2(n829), .ZN(n523) );
  INV_X1 U579 ( .A(n781), .ZN(n702) );
  NOR2_X1 U580 ( .A1(n703), .A2(n702), .ZN(n705) );
  INV_X1 U581 ( .A(KEYINPUT103), .ZN(n707) );
  NOR2_X1 U582 ( .A1(n757), .A2(n753), .ZN(n730) );
  NAND2_X1 U583 ( .A1(n974), .A2(n521), .ZN(n770) );
  NOR2_X1 U584 ( .A1(n816), .A2(n523), .ZN(n817) );
  NOR2_X1 U585 ( .A1(n599), .A2(n598), .ZN(n601) );
  BUF_X1 U586 ( .A(n547), .Z(n888) );
  XNOR2_X1 U587 ( .A(n601), .B(n600), .ZN(n978) );
  NOR2_X1 U588 ( .A1(n533), .A2(n532), .ZN(G160) );
  INV_X1 U589 ( .A(G2104), .ZN(n525) );
  NAND2_X1 U590 ( .A1(G101), .A2(n891), .ZN(n524) );
  XOR2_X1 U591 ( .A(KEYINPUT23), .B(n524), .Z(n528) );
  NAND2_X1 U592 ( .A1(G125), .A2(n887), .ZN(n526) );
  XOR2_X1 U593 ( .A(KEYINPUT65), .B(n526), .Z(n527) );
  NAND2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n533) );
  NAND2_X1 U595 ( .A1(n888), .A2(G113), .ZN(n531) );
  XOR2_X1 U596 ( .A(KEYINPUT17), .B(n529), .Z(n549) );
  NAND2_X1 U597 ( .A1(n517), .A2(G137), .ZN(n530) );
  NAND2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n532) );
  INV_X1 U599 ( .A(G651), .ZN(n539) );
  NOR2_X1 U600 ( .A1(G543), .A2(n539), .ZN(n535) );
  XNOR2_X1 U601 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n655) );
  NAND2_X1 U603 ( .A1(G62), .A2(n655), .ZN(n537) );
  NOR2_X4 U604 ( .A1(G651), .A2(n538), .ZN(n656) );
  NAND2_X1 U605 ( .A1(G50), .A2(n656), .ZN(n536) );
  NAND2_X1 U606 ( .A1(n537), .A2(n536), .ZN(n543) );
  NOR2_X1 U607 ( .A1(G651), .A2(G543), .ZN(n650) );
  NAND2_X1 U608 ( .A1(G88), .A2(n650), .ZN(n541) );
  NOR2_X2 U609 ( .A1(n538), .A2(n539), .ZN(n651) );
  NAND2_X1 U610 ( .A1(G75), .A2(n651), .ZN(n540) );
  NAND2_X1 U611 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U612 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n544), .B(KEYINPUT86), .ZN(G166) );
  INV_X1 U614 ( .A(G166), .ZN(G303) );
  NAND2_X1 U615 ( .A1(G126), .A2(n887), .ZN(n546) );
  NAND2_X1 U616 ( .A1(G102), .A2(n891), .ZN(n545) );
  NAND2_X1 U617 ( .A1(n547), .A2(G114), .ZN(n548) );
  XOR2_X1 U618 ( .A(KEYINPUT90), .B(n548), .Z(n550) );
  NAND2_X1 U619 ( .A1(n519), .A2(n551), .ZN(n552) );
  NAND2_X1 U620 ( .A1(G64), .A2(n655), .ZN(n554) );
  NAND2_X1 U621 ( .A1(G52), .A2(n656), .ZN(n553) );
  NAND2_X1 U622 ( .A1(n554), .A2(n553), .ZN(n559) );
  NAND2_X1 U623 ( .A1(G90), .A2(n650), .ZN(n556) );
  NAND2_X1 U624 ( .A1(G77), .A2(n651), .ZN(n555) );
  NAND2_X1 U625 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U626 ( .A(KEYINPUT9), .B(n557), .Z(n558) );
  NOR2_X1 U627 ( .A1(n559), .A2(n558), .ZN(G171) );
  AND2_X1 U628 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U629 ( .A1(G65), .A2(n655), .ZN(n561) );
  NAND2_X1 U630 ( .A1(G53), .A2(n656), .ZN(n560) );
  NAND2_X1 U631 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U632 ( .A1(G91), .A2(n650), .ZN(n563) );
  NAND2_X1 U633 ( .A1(G78), .A2(n651), .ZN(n562) );
  NAND2_X1 U634 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U635 ( .A1(n565), .A2(n564), .ZN(n979) );
  INV_X1 U636 ( .A(n979), .ZN(G299) );
  INV_X1 U637 ( .A(G82), .ZN(G220) );
  INV_X1 U638 ( .A(G57), .ZN(G237) );
  NAND2_X1 U639 ( .A1(n650), .A2(G89), .ZN(n566) );
  XNOR2_X1 U640 ( .A(n566), .B(KEYINPUT4), .ZN(n568) );
  NAND2_X1 U641 ( .A1(G76), .A2(n651), .ZN(n567) );
  NAND2_X1 U642 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U643 ( .A(KEYINPUT5), .B(n569), .ZN(n576) );
  XNOR2_X1 U644 ( .A(KEYINPUT76), .B(KEYINPUT6), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n655), .A2(G63), .ZN(n572) );
  NAND2_X1 U646 ( .A1(n656), .A2(G51), .ZN(n570) );
  XOR2_X1 U647 ( .A(KEYINPUT75), .B(n570), .Z(n571) );
  NAND2_X1 U648 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U649 ( .A(n574), .B(n573), .Z(n575) );
  NAND2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U651 ( .A(KEYINPUT7), .B(n577), .ZN(G168) );
  XOR2_X1 U652 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U653 ( .A1(G7), .A2(G661), .ZN(n578) );
  XNOR2_X1 U654 ( .A(n578), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U655 ( .A(G223), .ZN(n843) );
  NAND2_X1 U656 ( .A1(n843), .A2(G567), .ZN(n579) );
  XOR2_X1 U657 ( .A(KEYINPUT11), .B(n579), .Z(G234) );
  NAND2_X1 U658 ( .A1(n650), .A2(G81), .ZN(n580) );
  XNOR2_X1 U659 ( .A(n580), .B(KEYINPUT12), .ZN(n582) );
  NAND2_X1 U660 ( .A1(G68), .A2(n651), .ZN(n581) );
  NAND2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U662 ( .A(KEYINPUT13), .B(n583), .Z(n587) );
  NAND2_X1 U663 ( .A1(G56), .A2(n655), .ZN(n584) );
  XNOR2_X1 U664 ( .A(n584), .B(KEYINPUT69), .ZN(n585) );
  XNOR2_X1 U665 ( .A(n585), .B(KEYINPUT14), .ZN(n586) );
  NOR2_X1 U666 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U667 ( .A1(n656), .A2(G43), .ZN(n588) );
  NAND2_X1 U668 ( .A1(n589), .A2(n588), .ZN(n977) );
  INV_X1 U669 ( .A(n977), .ZN(n590) );
  NAND2_X1 U670 ( .A1(n590), .A2(G860), .ZN(G153) );
  XOR2_X1 U671 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  INV_X1 U672 ( .A(G868), .ZN(n670) );
  NOR2_X1 U673 ( .A1(G301), .A2(n670), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n656), .A2(G54), .ZN(n591) );
  XNOR2_X1 U675 ( .A(n591), .B(KEYINPUT72), .ZN(n593) );
  NAND2_X1 U676 ( .A1(G79), .A2(n651), .ZN(n592) );
  NAND2_X1 U677 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U678 ( .A(n594), .B(KEYINPUT73), .ZN(n596) );
  NAND2_X1 U679 ( .A1(G66), .A2(n655), .ZN(n595) );
  NAND2_X1 U680 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U681 ( .A1(G92), .A2(n650), .ZN(n597) );
  XNOR2_X1 U682 ( .A(KEYINPUT71), .B(n597), .ZN(n598) );
  XOR2_X1 U683 ( .A(KEYINPUT74), .B(KEYINPUT15), .Z(n600) );
  INV_X1 U684 ( .A(n978), .ZN(n912) );
  NOR2_X1 U685 ( .A1(n912), .A2(G868), .ZN(n602) );
  NOR2_X1 U686 ( .A1(n603), .A2(n602), .ZN(G284) );
  NOR2_X1 U687 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U688 ( .A1(G286), .A2(n670), .ZN(n604) );
  NOR2_X1 U689 ( .A1(n605), .A2(n604), .ZN(G297) );
  INV_X1 U690 ( .A(G559), .ZN(n606) );
  NOR2_X1 U691 ( .A1(G860), .A2(n606), .ZN(n607) );
  XNOR2_X1 U692 ( .A(KEYINPUT77), .B(n607), .ZN(n608) );
  NAND2_X1 U693 ( .A1(n608), .A2(n978), .ZN(n609) );
  XNOR2_X1 U694 ( .A(n609), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U695 ( .A1(G868), .A2(n978), .ZN(n610) );
  NOR2_X1 U696 ( .A1(G559), .A2(n610), .ZN(n611) );
  XNOR2_X1 U697 ( .A(n611), .B(KEYINPUT78), .ZN(n613) );
  NOR2_X1 U698 ( .A1(n977), .A2(G868), .ZN(n612) );
  NOR2_X1 U699 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U700 ( .A1(n887), .A2(G123), .ZN(n614) );
  XNOR2_X1 U701 ( .A(n614), .B(KEYINPUT18), .ZN(n616) );
  NAND2_X1 U702 ( .A1(G111), .A2(n888), .ZN(n615) );
  NAND2_X1 U703 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U704 ( .A1(G99), .A2(n891), .ZN(n618) );
  NAND2_X1 U705 ( .A1(G135), .A2(n517), .ZN(n617) );
  NAND2_X1 U706 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U707 ( .A1(n620), .A2(n619), .ZN(n925) );
  XNOR2_X1 U708 ( .A(n925), .B(G2096), .ZN(n622) );
  INV_X1 U709 ( .A(G2100), .ZN(n621) );
  NAND2_X1 U710 ( .A1(n622), .A2(n621), .ZN(G156) );
  NAND2_X1 U711 ( .A1(G559), .A2(n978), .ZN(n667) );
  XNOR2_X1 U712 ( .A(n977), .B(n667), .ZN(n623) );
  NOR2_X1 U713 ( .A1(n623), .A2(G860), .ZN(n632) );
  NAND2_X1 U714 ( .A1(G67), .A2(n655), .ZN(n625) );
  NAND2_X1 U715 ( .A1(G55), .A2(n656), .ZN(n624) );
  NAND2_X1 U716 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U717 ( .A(KEYINPUT80), .B(n626), .ZN(n631) );
  NAND2_X1 U718 ( .A1(G93), .A2(n650), .ZN(n628) );
  NAND2_X1 U719 ( .A1(G80), .A2(n651), .ZN(n627) );
  NAND2_X1 U720 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U721 ( .A(KEYINPUT79), .B(n629), .Z(n630) );
  OR2_X1 U722 ( .A1(n631), .A2(n630), .ZN(n669) );
  XOR2_X1 U723 ( .A(n632), .B(n669), .Z(G145) );
  NAND2_X1 U724 ( .A1(G86), .A2(n650), .ZN(n634) );
  NAND2_X1 U725 ( .A1(G61), .A2(n655), .ZN(n633) );
  NAND2_X1 U726 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U727 ( .A(KEYINPUT83), .B(n635), .Z(n638) );
  NAND2_X1 U728 ( .A1(n651), .A2(G73), .ZN(n636) );
  XOR2_X1 U729 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U730 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U731 ( .A(n639), .B(KEYINPUT84), .ZN(n641) );
  NAND2_X1 U732 ( .A1(G48), .A2(n656), .ZN(n640) );
  NAND2_X1 U733 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U734 ( .A(KEYINPUT85), .B(n642), .Z(G305) );
  NAND2_X1 U735 ( .A1(n656), .A2(G49), .ZN(n643) );
  XOR2_X1 U736 ( .A(KEYINPUT81), .B(n643), .Z(n645) );
  NAND2_X1 U737 ( .A1(G651), .A2(G74), .ZN(n644) );
  NAND2_X1 U738 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U739 ( .A1(n655), .A2(n646), .ZN(n647) );
  XNOR2_X1 U740 ( .A(n647), .B(KEYINPUT82), .ZN(n649) );
  NAND2_X1 U741 ( .A1(G87), .A2(n538), .ZN(n648) );
  NAND2_X1 U742 ( .A1(n649), .A2(n648), .ZN(G288) );
  NAND2_X1 U743 ( .A1(G85), .A2(n650), .ZN(n653) );
  NAND2_X1 U744 ( .A1(G72), .A2(n651), .ZN(n652) );
  NAND2_X1 U745 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U746 ( .A(KEYINPUT66), .B(n654), .Z(n660) );
  NAND2_X1 U747 ( .A1(G60), .A2(n655), .ZN(n658) );
  NAND2_X1 U748 ( .A1(G47), .A2(n656), .ZN(n657) );
  AND2_X1 U749 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U750 ( .A1(n660), .A2(n659), .ZN(G290) );
  XNOR2_X1 U751 ( .A(KEYINPUT19), .B(G299), .ZN(n661) );
  XNOR2_X1 U752 ( .A(n661), .B(n977), .ZN(n664) );
  XOR2_X1 U753 ( .A(n669), .B(G305), .Z(n662) );
  XNOR2_X1 U754 ( .A(n662), .B(G288), .ZN(n663) );
  XNOR2_X1 U755 ( .A(n664), .B(n663), .ZN(n666) );
  XNOR2_X1 U756 ( .A(G290), .B(G303), .ZN(n665) );
  XNOR2_X1 U757 ( .A(n666), .B(n665), .ZN(n913) );
  XNOR2_X1 U758 ( .A(n667), .B(n913), .ZN(n668) );
  NAND2_X1 U759 ( .A1(n668), .A2(G868), .ZN(n672) );
  NAND2_X1 U760 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U761 ( .A1(n672), .A2(n671), .ZN(G295) );
  XOR2_X1 U762 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n676) );
  NAND2_X1 U763 ( .A1(G2078), .A2(G2084), .ZN(n673) );
  XOR2_X1 U764 ( .A(KEYINPUT20), .B(n673), .Z(n674) );
  NAND2_X1 U765 ( .A1(n674), .A2(G2090), .ZN(n675) );
  XNOR2_X1 U766 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U767 ( .A1(G2072), .A2(n677), .ZN(G158) );
  XNOR2_X1 U768 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U769 ( .A(KEYINPUT68), .B(G132), .Z(G219) );
  NAND2_X1 U770 ( .A1(G69), .A2(G120), .ZN(n678) );
  NOR2_X1 U771 ( .A1(G237), .A2(n678), .ZN(n679) );
  NAND2_X1 U772 ( .A1(G108), .A2(n679), .ZN(n849) );
  NAND2_X1 U773 ( .A1(n849), .A2(G567), .ZN(n685) );
  NOR2_X1 U774 ( .A1(G219), .A2(G220), .ZN(n680) );
  XOR2_X1 U775 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U776 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U777 ( .A1(G96), .A2(n682), .ZN(n848) );
  NAND2_X1 U778 ( .A1(G2106), .A2(n848), .ZN(n683) );
  XNOR2_X1 U779 ( .A(KEYINPUT88), .B(n683), .ZN(n684) );
  NAND2_X1 U780 ( .A1(n685), .A2(n684), .ZN(n850) );
  NAND2_X1 U781 ( .A1(G661), .A2(G483), .ZN(n686) );
  XOR2_X1 U782 ( .A(KEYINPUT89), .B(n686), .Z(n687) );
  NOR2_X1 U783 ( .A1(n850), .A2(n687), .ZN(n846) );
  NAND2_X1 U784 ( .A1(n846), .A2(G36), .ZN(G176) );
  NAND2_X1 U785 ( .A1(G160), .A2(G40), .ZN(n782) );
  INV_X1 U786 ( .A(n782), .ZN(n690) );
  XNOR2_X2 U787 ( .A(n689), .B(KEYINPUT64), .ZN(n781) );
  NAND2_X1 U788 ( .A1(G1956), .A2(n709), .ZN(n691) );
  XNOR2_X1 U789 ( .A(KEYINPUT101), .B(n691), .ZN(n695) );
  XOR2_X1 U790 ( .A(KEYINPUT100), .B(KEYINPUT27), .Z(n692) );
  NOR2_X1 U791 ( .A1(n695), .A2(n694), .ZN(n698) );
  XOR2_X1 U792 ( .A(KEYINPUT102), .B(KEYINPUT28), .Z(n696) );
  XNOR2_X1 U793 ( .A(n697), .B(n696), .ZN(n718) );
  INV_X1 U794 ( .A(n718), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n698), .A2(n979), .ZN(n699) );
  AND2_X1 U796 ( .A1(n709), .A2(G1341), .ZN(n701) );
  NOR2_X1 U797 ( .A1(n701), .A2(n977), .ZN(n715) );
  INV_X1 U798 ( .A(G1996), .ZN(n954) );
  OR2_X1 U799 ( .A1(n782), .A2(n954), .ZN(n703) );
  INV_X1 U800 ( .A(KEYINPUT26), .ZN(n704) );
  XNOR2_X1 U801 ( .A(n705), .B(n704), .ZN(n716) );
  NAND2_X1 U802 ( .A1(n715), .A2(n706), .ZN(n708) );
  NOR2_X1 U803 ( .A1(n725), .A2(G1348), .ZN(n711) );
  NOR2_X1 U804 ( .A1(G2067), .A2(n709), .ZN(n710) );
  NOR2_X1 U805 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U806 ( .A(n714), .B(KEYINPUT104), .ZN(n721) );
  AND2_X1 U807 ( .A1(n716), .A2(n715), .ZN(n717) );
  OR2_X1 U808 ( .A1(n978), .A2(n717), .ZN(n719) );
  AND2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U810 ( .A1(n721), .A2(n720), .ZN(n722) );
  OR2_X1 U811 ( .A1(n725), .A2(G1961), .ZN(n727) );
  XNOR2_X1 U812 ( .A(G2078), .B(KEYINPUT25), .ZN(n953) );
  NAND2_X1 U813 ( .A1(n725), .A2(n953), .ZN(n726) );
  NAND2_X1 U814 ( .A1(n727), .A2(n726), .ZN(n729) );
  NAND2_X1 U815 ( .A1(n729), .A2(G171), .ZN(n750) );
  AND2_X1 U816 ( .A1(n750), .A2(G286), .ZN(n728) );
  NAND2_X1 U817 ( .A1(n749), .A2(n728), .ZN(n738) );
  INV_X1 U818 ( .A(G286), .ZN(n736) );
  NOR2_X1 U819 ( .A1(G171), .A2(n729), .ZN(n734) );
  NOR2_X1 U820 ( .A1(G1966), .A2(n778), .ZN(n757) );
  NOR2_X1 U821 ( .A1(G2084), .A2(n709), .ZN(n753) );
  NAND2_X1 U822 ( .A1(n730), .A2(G8), .ZN(n731) );
  XNOR2_X1 U823 ( .A(n731), .B(KEYINPUT30), .ZN(n732) );
  NOR2_X1 U824 ( .A1(G168), .A2(n732), .ZN(n733) );
  NOR2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U826 ( .A(n735), .B(KEYINPUT31), .Z(n751) );
  OR2_X1 U827 ( .A1(n736), .A2(n751), .ZN(n737) );
  AND2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n740) );
  XNOR2_X1 U829 ( .A(n740), .B(n739), .ZN(n745) );
  NOR2_X1 U830 ( .A1(G1971), .A2(n778), .ZN(n742) );
  NOR2_X1 U831 ( .A1(G2090), .A2(n709), .ZN(n741) );
  NOR2_X1 U832 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U833 ( .A1(n743), .A2(G303), .ZN(n744) );
  NAND2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n746), .A2(G8), .ZN(n748) );
  XOR2_X1 U836 ( .A(KEYINPUT106), .B(KEYINPUT32), .Z(n747) );
  XNOR2_X1 U837 ( .A(n748), .B(n747), .ZN(n759) );
  NAND2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n752) );
  NAND2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n755) );
  NAND2_X1 U840 ( .A1(G8), .A2(n753), .ZN(n754) );
  NAND2_X1 U841 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U842 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U843 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U844 ( .A(n760), .B(KEYINPUT107), .ZN(n772) );
  NOR2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n983) );
  NOR2_X1 U846 ( .A1(G303), .A2(G1971), .ZN(n761) );
  XNOR2_X1 U847 ( .A(KEYINPUT108), .B(n761), .ZN(n762) );
  NOR2_X1 U848 ( .A1(n983), .A2(n762), .ZN(n763) );
  XOR2_X1 U849 ( .A(KEYINPUT109), .B(n763), .Z(n764) );
  NAND2_X1 U850 ( .A1(n772), .A2(n764), .ZN(n766) );
  NAND2_X1 U851 ( .A1(G288), .A2(G1976), .ZN(n765) );
  XNOR2_X1 U852 ( .A(n765), .B(KEYINPUT110), .ZN(n984) );
  NAND2_X1 U853 ( .A1(n766), .A2(n984), .ZN(n767) );
  NOR2_X1 U854 ( .A1(n778), .A2(n767), .ZN(n768) );
  NOR2_X1 U855 ( .A1(KEYINPUT33), .A2(n768), .ZN(n771) );
  XOR2_X1 U856 ( .A(G1981), .B(G305), .Z(n974) );
  NAND2_X1 U857 ( .A1(n983), .A2(KEYINPUT33), .ZN(n769) );
  NOR2_X1 U858 ( .A1(G2090), .A2(G303), .ZN(n773) );
  NAND2_X1 U859 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n772), .A2(n774), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n775), .A2(n778), .ZN(n780) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U863 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  OR2_X1 U864 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n522), .A2(n520), .ZN(n818) );
  NOR2_X1 U866 ( .A1(n782), .A2(n781), .ZN(n829) );
  XNOR2_X1 U867 ( .A(G2067), .B(KEYINPUT37), .ZN(n827) );
  NAND2_X1 U868 ( .A1(n887), .A2(G128), .ZN(n783) );
  XOR2_X1 U869 ( .A(KEYINPUT93), .B(n783), .Z(n785) );
  NAND2_X1 U870 ( .A1(n888), .A2(G116), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n787) );
  XNOR2_X1 U872 ( .A(KEYINPUT94), .B(KEYINPUT35), .ZN(n786) );
  XNOR2_X1 U873 ( .A(n787), .B(n786), .ZN(n793) );
  NAND2_X1 U874 ( .A1(n891), .A2(G104), .ZN(n788) );
  XNOR2_X1 U875 ( .A(n788), .B(KEYINPUT92), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G140), .A2(n517), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U878 ( .A(KEYINPUT34), .B(n791), .Z(n792) );
  NAND2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U880 ( .A(KEYINPUT36), .B(n794), .Z(n906) );
  OR2_X1 U881 ( .A1(n827), .A2(n906), .ZN(n795) );
  XNOR2_X1 U882 ( .A(n795), .B(KEYINPUT95), .ZN(n944) );
  NAND2_X1 U883 ( .A1(n829), .A2(n944), .ZN(n825) );
  NAND2_X1 U884 ( .A1(G129), .A2(n887), .ZN(n797) );
  NAND2_X1 U885 ( .A1(G117), .A2(n888), .ZN(n796) );
  NAND2_X1 U886 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U887 ( .A(KEYINPUT98), .B(n798), .ZN(n801) );
  NAND2_X1 U888 ( .A1(n891), .A2(G105), .ZN(n799) );
  XOR2_X1 U889 ( .A(KEYINPUT38), .B(n799), .Z(n800) );
  NOR2_X1 U890 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U891 ( .A1(n517), .A2(G141), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n803), .A2(n802), .ZN(n884) );
  NAND2_X1 U893 ( .A1(n884), .A2(G1996), .ZN(n813) );
  NAND2_X1 U894 ( .A1(G119), .A2(n887), .ZN(n805) );
  NAND2_X1 U895 ( .A1(G131), .A2(n517), .ZN(n804) );
  NAND2_X1 U896 ( .A1(n805), .A2(n804), .ZN(n808) );
  NAND2_X1 U897 ( .A1(n891), .A2(G95), .ZN(n806) );
  XOR2_X1 U898 ( .A(KEYINPUT96), .B(n806), .Z(n807) );
  NOR2_X1 U899 ( .A1(n808), .A2(n807), .ZN(n810) );
  NAND2_X1 U900 ( .A1(n888), .A2(G107), .ZN(n809) );
  NAND2_X1 U901 ( .A1(n810), .A2(n809), .ZN(n885) );
  NAND2_X1 U902 ( .A1(G1991), .A2(n885), .ZN(n811) );
  XOR2_X1 U903 ( .A(KEYINPUT97), .B(n811), .Z(n812) );
  NAND2_X1 U904 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U905 ( .A(n814), .B(KEYINPUT99), .ZN(n934) );
  INV_X1 U906 ( .A(n934), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n815), .A2(n829), .ZN(n819) );
  NAND2_X1 U908 ( .A1(n825), .A2(n819), .ZN(n816) );
  XNOR2_X1 U909 ( .A(G1986), .B(G290), .ZN(n988) );
  NAND2_X1 U910 ( .A1(n818), .A2(n817), .ZN(n832) );
  NOR2_X1 U911 ( .A1(G1996), .A2(n884), .ZN(n931) );
  INV_X1 U912 ( .A(n819), .ZN(n822) );
  NOR2_X1 U913 ( .A1(G1991), .A2(n885), .ZN(n929) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U915 ( .A1(n929), .A2(n820), .ZN(n821) );
  NOR2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U917 ( .A1(n931), .A2(n823), .ZN(n824) );
  XNOR2_X1 U918 ( .A(n824), .B(KEYINPUT39), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n826), .A2(n825), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n906), .A2(n827), .ZN(n926) );
  NAND2_X1 U921 ( .A1(n828), .A2(n926), .ZN(n830) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U924 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U925 ( .A(G1348), .B(G2454), .ZN(n834) );
  XNOR2_X1 U926 ( .A(n834), .B(G2430), .ZN(n835) );
  XNOR2_X1 U927 ( .A(n835), .B(G1341), .ZN(n841) );
  XOR2_X1 U928 ( .A(G2443), .B(G2427), .Z(n837) );
  XNOR2_X1 U929 ( .A(G2438), .B(G2446), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n837), .B(n836), .ZN(n839) );
  XOR2_X1 U931 ( .A(G2451), .B(G2435), .Z(n838) );
  XNOR2_X1 U932 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U933 ( .A(n841), .B(n840), .ZN(n842) );
  NAND2_X1 U934 ( .A1(n842), .A2(G14), .ZN(n917) );
  XNOR2_X1 U935 ( .A(KEYINPUT111), .B(n917), .ZN(G401) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U938 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n845) );
  XNOR2_X1 U940 ( .A(KEYINPUT112), .B(n845), .ZN(n847) );
  NAND2_X1 U941 ( .A1(n847), .A2(n846), .ZN(G188) );
  INV_X1 U943 ( .A(G120), .ZN(G236) );
  INV_X1 U944 ( .A(G96), .ZN(G221) );
  INV_X1 U945 ( .A(G69), .ZN(G235) );
  NOR2_X1 U946 ( .A1(n849), .A2(n848), .ZN(G325) );
  INV_X1 U947 ( .A(G325), .ZN(G261) );
  INV_X1 U948 ( .A(n850), .ZN(G319) );
  XOR2_X1 U949 ( .A(KEYINPUT42), .B(G2084), .Z(n852) );
  XNOR2_X1 U950 ( .A(G2090), .B(G2072), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U952 ( .A(n853), .B(G2100), .Z(n855) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2078), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U955 ( .A(G2096), .B(KEYINPUT43), .Z(n857) );
  XNOR2_X1 U956 ( .A(KEYINPUT113), .B(G2678), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U958 ( .A(n859), .B(n858), .Z(G227) );
  XOR2_X1 U959 ( .A(G1976), .B(G1961), .Z(n861) );
  XNOR2_X1 U960 ( .A(G1986), .B(G1971), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U962 ( .A(n862), .B(KEYINPUT41), .Z(n864) );
  XNOR2_X1 U963 ( .A(G1996), .B(G1991), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U965 ( .A(G2474), .B(G1981), .Z(n866) );
  XNOR2_X1 U966 ( .A(G1956), .B(G1966), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(G229) );
  NAND2_X1 U969 ( .A1(G100), .A2(n891), .ZN(n870) );
  NAND2_X1 U970 ( .A1(G112), .A2(n888), .ZN(n869) );
  NAND2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U972 ( .A(KEYINPUT114), .B(n871), .ZN(n876) );
  NAND2_X1 U973 ( .A1(n887), .A2(G124), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n872), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G136), .A2(n517), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U977 ( .A1(n876), .A2(n875), .ZN(G162) );
  NAND2_X1 U978 ( .A1(G103), .A2(n891), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G139), .A2(n517), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G127), .A2(n887), .ZN(n880) );
  NAND2_X1 U982 ( .A1(G115), .A2(n888), .ZN(n879) );
  NAND2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n935) );
  XNOR2_X1 U986 ( .A(n935), .B(n884), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n886), .B(n885), .ZN(n905) );
  XOR2_X1 U988 ( .A(KEYINPUT46), .B(KEYINPUT116), .Z(n900) );
  NAND2_X1 U989 ( .A1(G130), .A2(n887), .ZN(n890) );
  NAND2_X1 U990 ( .A1(G118), .A2(n888), .ZN(n889) );
  NAND2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n897) );
  NAND2_X1 U992 ( .A1(G106), .A2(n891), .ZN(n893) );
  NAND2_X1 U993 ( .A1(G142), .A2(n517), .ZN(n892) );
  NAND2_X1 U994 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U995 ( .A(KEYINPUT45), .B(n894), .ZN(n895) );
  XNOR2_X1 U996 ( .A(KEYINPUT115), .B(n895), .ZN(n896) );
  NOR2_X1 U997 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n898), .B(KEYINPUT48), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U1000 ( .A(n901), .B(KEYINPUT117), .Z(n903) );
  XNOR2_X1 U1001 ( .A(n925), .B(KEYINPUT118), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1003 ( .A(n905), .B(n904), .Z(n908) );
  XOR2_X1 U1004 ( .A(G160), .B(n906), .Z(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n910) );
  XOR2_X1 U1006 ( .A(G162), .B(G164), .Z(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n911), .ZN(G395) );
  XNOR2_X1 U1009 ( .A(G171), .B(n912), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n915), .B(G286), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n916), .ZN(G397) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n917), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n918) );
  XOR2_X1 U1015 ( .A(KEYINPUT49), .B(n918), .Z(n919) );
  XNOR2_X1 U1016 ( .A(n919), .B(KEYINPUT119), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n923) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1022 ( .A(G2084), .B(G160), .Z(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n942) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1028 ( .A(KEYINPUT51), .B(n932), .Z(n933) );
  NAND2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n940) );
  XOR2_X1 U1030 ( .A(G2072), .B(n935), .Z(n937) );
  XOR2_X1 U1031 ( .A(G164), .B(G2078), .Z(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1033 ( .A(KEYINPUT50), .B(n938), .Z(n939) );
  NOR2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n945), .ZN(n946) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n969) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n969), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n947), .A2(G29), .ZN(n1029) );
  XOR2_X1 U1041 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n962) );
  XOR2_X1 U1042 ( .A(G1991), .B(G25), .Z(n952) );
  XNOR2_X1 U1043 ( .A(G2067), .B(G26), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(G2072), .B(G33), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(n950), .B(KEYINPUT120), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n959) );
  XOR2_X1 U1048 ( .A(n953), .B(G27), .Z(n956) );
  XOR2_X1 U1049 ( .A(n954), .B(G32), .Z(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n957), .B(KEYINPUT121), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n960), .A2(G28), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(n962), .B(n961), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(G35), .B(G2090), .ZN(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n967) );
  XOR2_X1 U1057 ( .A(G2084), .B(G34), .Z(n965) );
  XNOR2_X1 U1058 ( .A(KEYINPUT54), .B(n965), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(n969), .B(n968), .ZN(n971) );
  INV_X1 U1061 ( .A(G29), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n972), .ZN(n1027) );
  XNOR2_X1 U1064 ( .A(G16), .B(KEYINPUT56), .ZN(n999) );
  XOR2_X1 U1065 ( .A(G168), .B(G1966), .Z(n973) );
  XNOR2_X1 U1066 ( .A(KEYINPUT123), .B(n973), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(n976), .B(KEYINPUT57), .ZN(n997) );
  XNOR2_X1 U1069 ( .A(n977), .B(G1341), .ZN(n995) );
  XNOR2_X1 U1070 ( .A(G1348), .B(n978), .ZN(n990) );
  XNOR2_X1 U1071 ( .A(n979), .B(G1956), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G166), .B(G1971), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(KEYINPUT124), .B(n986), .ZN(n987) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n992) );
  XOR2_X1 U1079 ( .A(G171), .B(G1961), .Z(n991) );
  NOR2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(KEYINPUT125), .B(n993), .ZN(n994) );
  NOR2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1084 ( .A1(n999), .A2(n998), .ZN(n1025) );
  INV_X1 U1085 ( .A(G16), .ZN(n1023) );
  XNOR2_X1 U1086 ( .A(G1986), .B(G24), .ZN(n1004) );
  XNOR2_X1 U1087 ( .A(G1971), .B(G22), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(G1976), .B(G23), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(KEYINPUT127), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(KEYINPUT58), .B(n1005), .ZN(n1018) );
  XOR2_X1 U1093 ( .A(G1348), .B(KEYINPUT59), .Z(n1006) );
  XNOR2_X1 U1094 ( .A(G4), .B(n1006), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(G20), .B(G1956), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(G1341), .B(G19), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G1981), .B(G6), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(n1013), .B(KEYINPUT60), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(G1966), .B(KEYINPUT126), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(G21), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(G5), .B(G1961), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1112 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

