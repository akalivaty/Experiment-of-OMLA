

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784;

  BUF_X1 U372 ( .A(n720), .Z(n353) );
  XNOR2_X1 U373 ( .A(n591), .B(n410), .ZN(n582) );
  OR2_X1 U374 ( .A1(n654), .A2(G902), .ZN(n411) );
  XOR2_X1 U375 ( .A(G116), .B(KEYINPUT3), .Z(n527) );
  INV_X2 U376 ( .A(G125), .ZN(n399) );
  XNOR2_X1 U377 ( .A(n351), .B(n557), .ZN(n570) );
  NAND2_X1 U378 ( .A1(n556), .A2(n781), .ZN(n351) );
  XNOR2_X1 U379 ( .A(n352), .B(n472), .ZN(n761) );
  XNOR2_X1 U380 ( .A(n400), .B(n470), .ZN(n352) );
  INV_X2 U381 ( .A(G104), .ZN(n451) );
  NAND2_X1 U382 ( .A1(n441), .A2(n439), .ZN(n632) );
  INV_X1 U383 ( .A(G953), .ZN(n774) );
  XOR2_X1 U384 ( .A(n506), .B(G116), .Z(n354) );
  XNOR2_X2 U385 ( .A(n521), .B(n522), .ZN(n536) );
  INV_X1 U386 ( .A(n582), .ZN(n559) );
  INV_X1 U387 ( .A(n364), .ZN(n359) );
  INV_X4 U388 ( .A(G128), .ZN(n450) );
  AND2_X2 U389 ( .A1(n363), .A2(n371), .ZN(n420) );
  XNOR2_X1 U390 ( .A(n630), .B(n629), .ZN(n363) );
  NOR2_X1 U391 ( .A1(n386), .A2(n381), .ZN(n405) );
  AND2_X1 U392 ( .A1(n431), .A2(n430), .ZN(n402) );
  AND2_X1 U393 ( .A1(n433), .A2(n599), .ZN(n431) );
  NOR2_X1 U394 ( .A1(n597), .A2(n596), .ZN(n610) );
  OR2_X1 U395 ( .A1(n552), .A2(n416), .ZN(n415) );
  NOR2_X1 U396 ( .A1(n444), .A2(KEYINPUT1), .ZN(n442) );
  OR2_X2 U397 ( .A1(n661), .A2(n445), .ZN(n444) );
  XNOR2_X1 U398 ( .A(n506), .B(KEYINPUT4), .ZN(n521) );
  XNOR2_X1 U399 ( .A(n390), .B(G119), .ZN(n470) );
  NOR2_X1 U400 ( .A1(n404), .A2(G237), .ZN(n532) );
  XOR2_X1 U401 ( .A(G902), .B(KEYINPUT15), .Z(n641) );
  XNOR2_X1 U402 ( .A(KEYINPUT85), .B(KEYINPUT48), .ZN(n629) );
  INV_X1 U403 ( .A(KEYINPUT82), .ZN(n364) );
  NAND2_X1 U404 ( .A1(n355), .A2(n772), .ZN(n643) );
  NOR2_X1 U405 ( .A1(n360), .A2(n356), .ZN(n355) );
  NAND2_X1 U406 ( .A1(n358), .A2(n357), .ZN(n356) );
  NAND2_X1 U407 ( .A1(n574), .A2(n359), .ZN(n357) );
  NAND2_X1 U408 ( .A1(n645), .A2(n359), .ZN(n358) );
  NOR2_X1 U409 ( .A1(n645), .A2(n361), .ZN(n360) );
  NAND2_X1 U410 ( .A1(n362), .A2(n364), .ZN(n361) );
  INV_X1 U411 ( .A(n574), .ZN(n362) );
  XNOR2_X2 U412 ( .A(n420), .B(n640), .ZN(n772) );
  XNOR2_X2 U413 ( .A(n573), .B(n572), .ZN(n645) );
  BUF_X1 U414 ( .A(n490), .Z(n365) );
  XNOR2_X1 U415 ( .A(n451), .B(G113), .ZN(n490) );
  NOR2_X2 U416 ( .A1(n648), .A2(n693), .ZN(n366) );
  NOR2_X2 U417 ( .A1(n648), .A2(n693), .ZN(n367) );
  BUF_X1 U418 ( .A(n779), .Z(n368) );
  XNOR2_X1 U419 ( .A(n516), .B(G146), .ZN(n533) );
  NAND2_X1 U420 ( .A1(n440), .A2(n447), .ZN(n439) );
  NOR2_X1 U421 ( .A1(n443), .A2(n442), .ZN(n441) );
  AND2_X1 U422 ( .A1(n444), .A2(KEYINPUT1), .ZN(n440) );
  NOR2_X1 U423 ( .A1(n778), .A2(n377), .ZN(n384) );
  OR2_X1 U424 ( .A1(KEYINPUT69), .A2(n619), .ZN(n622) );
  NAND2_X1 U425 ( .A1(n618), .A2(n387), .ZN(n386) );
  AND2_X1 U426 ( .A1(n437), .A2(n448), .ZN(n447) );
  NAND2_X1 U427 ( .A1(n525), .A2(n446), .ZN(n445) );
  INV_X1 U428 ( .A(G902), .ZN(n446) );
  NAND2_X1 U429 ( .A1(n438), .A2(n373), .ZN(n443) );
  XNOR2_X1 U430 ( .A(G140), .B(KEYINPUT98), .ZN(n491) );
  XNOR2_X1 U431 ( .A(n501), .B(n408), .ZN(n561) );
  XNOR2_X1 U432 ( .A(n409), .B(G475), .ZN(n408) );
  INV_X1 U433 ( .A(KEYINPUT13), .ZN(n409) );
  NAND2_X1 U434 ( .A1(n447), .A2(n444), .ZN(n603) );
  INV_X1 U435 ( .A(KEYINPUT6), .ZN(n410) );
  XNOR2_X1 U436 ( .A(n535), .B(n534), .ZN(n537) );
  XNOR2_X1 U437 ( .A(n533), .B(n370), .ZN(n534) );
  XNOR2_X1 U438 ( .A(n426), .B(n467), .ZN(n425) );
  XNOR2_X1 U439 ( .A(n465), .B(G128), .ZN(n426) );
  XNOR2_X1 U440 ( .A(n391), .B(n388), .ZN(n466) );
  XNOR2_X1 U441 ( .A(n470), .B(n389), .ZN(n388) );
  INV_X1 U442 ( .A(KEYINPUT91), .ZN(n389) );
  INV_X1 U443 ( .A(n554), .ZN(n416) );
  XNOR2_X1 U444 ( .A(KEYINPUT30), .B(KEYINPUT105), .ZN(n592) );
  OR2_X1 U445 ( .A1(n461), .A2(n460), .ZN(n455) );
  NAND2_X1 U446 ( .A1(n385), .A2(n384), .ZN(n383) );
  NOR2_X1 U447 ( .A1(n715), .A2(n622), .ZN(n620) );
  NAND2_X1 U448 ( .A1(n449), .A2(G902), .ZN(n448) );
  XOR2_X1 U449 ( .A(KEYINPUT97), .B(G131), .Z(n494) );
  XOR2_X1 U450 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n492) );
  NAND2_X1 U451 ( .A1(n421), .A2(n545), .ZN(n694) );
  XNOR2_X1 U452 ( .A(G119), .B(G137), .ZN(n528) );
  INV_X1 U453 ( .A(G110), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n393), .B(n392), .ZN(n503) );
  INV_X1 U455 ( .A(KEYINPUT8), .ZN(n392) );
  NAND2_X1 U456 ( .A1(n774), .A2(G234), .ZN(n393) );
  XNOR2_X1 U457 ( .A(n412), .B(G107), .ZN(n502) );
  INV_X1 U458 ( .A(G122), .ZN(n412) );
  XNOR2_X1 U459 ( .A(n403), .B(KEYINPUT77), .ZN(n463) );
  NAND2_X1 U460 ( .A1(n464), .A2(G224), .ZN(n403) );
  XNOR2_X1 U461 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n462) );
  XNOR2_X1 U462 ( .A(n571), .B(KEYINPUT45), .ZN(n572) );
  NAND2_X1 U463 ( .A1(G237), .A2(G234), .ZN(n480) );
  NOR2_X1 U464 ( .A1(G237), .A2(G902), .ZN(n477) );
  INV_X1 U465 ( .A(KEYINPUT66), .ZN(n460) );
  XOR2_X1 U466 ( .A(G143), .B(G122), .Z(n497) );
  XOR2_X1 U467 ( .A(G107), .B(n533), .Z(n520) );
  NOR2_X1 U468 ( .A1(n603), .A2(n602), .ZN(n615) );
  XNOR2_X1 U469 ( .A(n394), .B(n376), .ZN(n602) );
  NOR2_X1 U470 ( .A1(n601), .A2(n701), .ZN(n394) );
  XNOR2_X1 U471 ( .A(n407), .B(n406), .ZN(n708) );
  INV_X1 U472 ( .A(KEYINPUT41), .ZN(n406) );
  NOR2_X1 U473 ( .A1(n714), .A2(n713), .ZN(n407) );
  INV_X1 U474 ( .A(n603), .ZN(n423) );
  XNOR2_X1 U475 ( .A(n469), .B(n468), .ZN(n650) );
  XNOR2_X1 U476 ( .A(n425), .B(n523), .ZN(n424) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n749) );
  XNOR2_X1 U478 ( .A(n505), .B(n419), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n354), .B(n504), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n507), .B(KEYINPUT7), .ZN(n419) );
  NOR2_X1 U481 ( .A1(G952), .A2(n774), .ZN(n754) );
  XNOR2_X1 U482 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U483 ( .A(n587), .B(KEYINPUT110), .ZN(n588) );
  INV_X1 U484 ( .A(KEYINPUT32), .ZN(n413) );
  NAND2_X1 U485 ( .A1(n456), .A2(n454), .ZN(n453) );
  AND2_X1 U486 ( .A1(n456), .A2(n452), .ZN(n369) );
  AND2_X1 U487 ( .A1(G210), .A2(n532), .ZN(n370) );
  AND2_X1 U488 ( .A1(n689), .A2(n688), .ZN(n371) );
  AND2_X1 U489 ( .A1(n626), .A2(KEYINPUT47), .ZN(n372) );
  BUF_X1 U490 ( .A(n549), .Z(n550) );
  OR2_X1 U491 ( .A1(n448), .A2(KEYINPUT1), .ZN(n373) );
  INV_X1 U492 ( .A(KEYINPUT1), .ZN(n526) );
  NAND2_X1 U493 ( .A1(n478), .A2(G210), .ZN(n374) );
  AND2_X1 U494 ( .A1(n449), .A2(n526), .ZN(n375) );
  INV_X1 U495 ( .A(n632), .ZN(n452) );
  XNOR2_X1 U496 ( .A(KEYINPUT107), .B(KEYINPUT28), .ZN(n376) );
  XNOR2_X1 U497 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n377) );
  XOR2_X1 U498 ( .A(n656), .B(n655), .Z(n378) );
  XOR2_X1 U499 ( .A(n663), .B(n662), .Z(n379) );
  XOR2_X1 U500 ( .A(n738), .B(n737), .Z(n380) );
  NAND2_X1 U501 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U502 ( .A1(n778), .A2(n377), .ZN(n382) );
  INV_X1 U503 ( .A(n784), .ZN(n385) );
  NAND2_X1 U504 ( .A1(n784), .A2(n377), .ZN(n387) );
  XNOR2_X1 U505 ( .A(n616), .B(n617), .ZN(n784) );
  XNOR2_X2 U506 ( .A(n614), .B(n613), .ZN(n778) );
  NAND2_X1 U507 ( .A1(n503), .A2(G221), .ZN(n391) );
  NAND2_X1 U508 ( .A1(n579), .A2(n697), .ZN(n601) );
  XNOR2_X2 U509 ( .A(n542), .B(n541), .ZN(n697) );
  INV_X1 U510 ( .A(n637), .ZN(n395) );
  BUF_X1 U511 ( .A(G104), .Z(n671) );
  XOR2_X1 U512 ( .A(KEYINPUT16), .B(KEYINPUT73), .Z(n471) );
  XNOR2_X1 U513 ( .A(n490), .B(n471), .ZN(n400) );
  NOR2_X1 U514 ( .A1(n455), .A2(n632), .ZN(n454) );
  OR2_X1 U515 ( .A1(n632), .A2(n461), .ZN(n459) );
  XNOR2_X1 U516 ( .A(n466), .B(n424), .ZN(n469) );
  XNOR2_X1 U517 ( .A(n537), .B(n536), .ZN(n654) );
  XNOR2_X2 U518 ( .A(n396), .B(n374), .ZN(n609) );
  NOR2_X2 U519 ( .A1(n735), .A2(n641), .ZN(n396) );
  BUF_X1 U520 ( .A(G953), .Z(n404) );
  XNOR2_X1 U521 ( .A(n414), .B(n413), .ZN(n780) );
  INV_X1 U522 ( .A(n435), .ZN(n397) );
  AND2_X1 U523 ( .A1(n398), .A2(n458), .ZN(n457) );
  NAND2_X1 U524 ( .A1(n553), .A2(n460), .ZN(n398) );
  NAND2_X1 U525 ( .A1(n459), .A2(n460), .ZN(n458) );
  NOR2_X2 U526 ( .A1(n564), .A2(n559), .ZN(n548) );
  NAND2_X1 U527 ( .A1(n546), .A2(n632), .ZN(n564) );
  XNOR2_X1 U528 ( .A(n436), .B(KEYINPUT35), .ZN(n779) );
  NOR2_X2 U529 ( .A1(n553), .A2(n415), .ZN(n414) );
  NAND2_X1 U530 ( .A1(n402), .A2(n432), .ZN(n436) );
  XNOR2_X2 U531 ( .A(n399), .B(G146), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n457), .A2(n453), .ZN(n543) );
  XNOR2_X1 U533 ( .A(n401), .B(n475), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(n401) );
  XNOR2_X1 U535 ( .A(n761), .B(n428), .ZN(n735) );
  XNOR2_X1 U536 ( .A(n463), .B(n462), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n476), .B(n521), .ZN(n428) );
  NAND2_X1 U538 ( .A1(n405), .A2(n628), .ZN(n630) );
  XNOR2_X1 U539 ( .A(n500), .B(n499), .ZN(n743) );
  XNOR2_X2 U540 ( .A(n411), .B(G472), .ZN(n591) );
  XNOR2_X2 U541 ( .A(n515), .B(KEYINPUT22), .ZN(n553) );
  NAND2_X1 U542 ( .A1(n420), .A2(KEYINPUT2), .ZN(n647) );
  INV_X1 U543 ( .A(n697), .ZN(n421) );
  NOR2_X2 U544 ( .A1(n697), .A2(n422), .ZN(n594) );
  NAND2_X1 U545 ( .A1(n423), .A2(n545), .ZN(n422) );
  INV_X1 U546 ( .A(n550), .ZN(n435) );
  AND2_X1 U547 ( .A1(n550), .A2(n551), .ZN(n429) );
  NAND2_X1 U548 ( .A1(n397), .A2(n705), .ZN(n565) );
  NAND2_X1 U549 ( .A1(n397), .A2(n594), .ZN(n566) );
  NAND2_X1 U550 ( .A1(n435), .A2(n434), .ZN(n433) );
  NAND2_X1 U551 ( .A1(n720), .A2(n429), .ZN(n430) );
  OR2_X1 U552 ( .A1(n720), .A2(n551), .ZN(n432) );
  INV_X1 U553 ( .A(n551), .ZN(n434) );
  NAND2_X1 U554 ( .A1(n661), .A2(n449), .ZN(n437) );
  NAND2_X1 U555 ( .A1(n661), .A2(n375), .ZN(n438) );
  INV_X1 U556 ( .A(n525), .ZN(n449) );
  XNOR2_X2 U557 ( .A(n536), .B(n523), .ZN(n767) );
  XNOR2_X2 U558 ( .A(n450), .B(G143), .ZN(n506) );
  INV_X1 U559 ( .A(n553), .ZN(n456) );
  INV_X1 U560 ( .A(n701), .ZN(n461) );
  NOR2_X1 U561 ( .A1(n746), .A2(n754), .ZN(n748) );
  XNOR2_X1 U562 ( .A(n745), .B(n744), .ZN(n746) );
  NAND2_X1 U563 ( .A1(n367), .A2(G475), .ZN(n745) );
  INV_X1 U564 ( .A(n516), .ZN(n474) );
  XNOR2_X1 U565 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U566 ( .A(KEYINPUT0), .B(KEYINPUT86), .ZN(n488) );
  XNOR2_X1 U567 ( .A(n498), .B(n497), .ZN(n499) );
  INV_X1 U568 ( .A(KEYINPUT36), .ZN(n587) );
  INV_X1 U569 ( .A(KEYINPUT83), .ZN(n640) );
  XNOR2_X1 U570 ( .A(n743), .B(n742), .ZN(n744) );
  XNOR2_X1 U571 ( .A(n540), .B(n539), .ZN(n541) );
  INV_X1 U572 ( .A(KEYINPUT123), .ZN(n652) );
  INV_X1 U573 ( .A(G953), .ZN(n464) );
  XOR2_X1 U574 ( .A(G137), .B(G140), .Z(n523) );
  INV_X1 U575 ( .A(KEYINPUT76), .ZN(n465) );
  INV_X1 U576 ( .A(KEYINPUT24), .ZN(n467) );
  XOR2_X1 U577 ( .A(KEYINPUT10), .B(n473), .Z(n768) );
  XNOR2_X1 U578 ( .A(n768), .B(KEYINPUT23), .ZN(n468) );
  XNOR2_X1 U579 ( .A(n502), .B(n527), .ZN(n472) );
  XNOR2_X2 U580 ( .A(KEYINPUT68), .B(G101), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n477), .B(KEYINPUT75), .ZN(n478) );
  NAND2_X1 U582 ( .A1(G214), .A2(n478), .ZN(n710) );
  NAND2_X1 U583 ( .A1(n609), .A2(n710), .ZN(n585) );
  INV_X1 U584 ( .A(KEYINPUT19), .ZN(n479) );
  XNOR2_X1 U585 ( .A(n585), .B(n479), .ZN(n604) );
  XOR2_X1 U586 ( .A(KEYINPUT89), .B(KEYINPUT14), .Z(n481) );
  XNOR2_X1 U587 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U588 ( .A(KEYINPUT74), .B(n482), .ZN(n483) );
  NAND2_X1 U589 ( .A1(G952), .A2(n483), .ZN(n726) );
  NOR2_X1 U590 ( .A1(n404), .A2(n726), .ZN(n577) );
  AND2_X1 U591 ( .A1(n483), .A2(n404), .ZN(n484) );
  NAND2_X1 U592 ( .A1(G902), .A2(n484), .ZN(n575) );
  NOR2_X1 U593 ( .A1(G898), .A2(n575), .ZN(n485) );
  NOR2_X1 U594 ( .A1(n577), .A2(n485), .ZN(n486) );
  XNOR2_X1 U595 ( .A(n486), .B(KEYINPUT90), .ZN(n487) );
  NOR2_X2 U596 ( .A1(n604), .A2(n487), .ZN(n489) );
  XNOR2_X1 U597 ( .A(n489), .B(n488), .ZN(n549) );
  XNOR2_X1 U598 ( .A(n365), .B(n768), .ZN(n500) );
  XNOR2_X1 U599 ( .A(n492), .B(n491), .ZN(n496) );
  NAND2_X1 U600 ( .A1(n532), .A2(G214), .ZN(n493) );
  XNOR2_X1 U601 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U602 ( .A(n496), .B(n495), .ZN(n498) );
  NOR2_X1 U603 ( .A1(G902), .A2(n743), .ZN(n501) );
  XOR2_X1 U604 ( .A(n502), .B(G134), .Z(n505) );
  NAND2_X1 U605 ( .A1(G217), .A2(n503), .ZN(n504) );
  XOR2_X1 U606 ( .A(KEYINPUT9), .B(KEYINPUT99), .Z(n507) );
  NOR2_X1 U607 ( .A1(n749), .A2(G902), .ZN(n508) );
  XNOR2_X1 U608 ( .A(n508), .B(G478), .ZN(n562) );
  NAND2_X1 U609 ( .A1(n561), .A2(n562), .ZN(n713) );
  XOR2_X1 U610 ( .A(KEYINPUT93), .B(KEYINPUT20), .Z(n510) );
  INV_X1 U611 ( .A(n641), .ZN(n574) );
  NAND2_X1 U612 ( .A1(G234), .A2(n574), .ZN(n509) );
  XNOR2_X1 U613 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U614 ( .A(KEYINPUT92), .B(n511), .ZN(n538) );
  NAND2_X1 U615 ( .A1(G221), .A2(n538), .ZN(n513) );
  XOR2_X1 U616 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n512) );
  XNOR2_X1 U617 ( .A(n513), .B(n512), .ZN(n698) );
  NOR2_X1 U618 ( .A1(n713), .A2(n698), .ZN(n514) );
  NAND2_X1 U619 ( .A1(n549), .A2(n514), .ZN(n515) );
  XNOR2_X1 U620 ( .A(G110), .B(n671), .ZN(n518) );
  NAND2_X1 U621 ( .A1(G227), .A2(n774), .ZN(n517) );
  XNOR2_X1 U622 ( .A(n520), .B(n519), .ZN(n524) );
  XNOR2_X1 U623 ( .A(G131), .B(G134), .ZN(n522) );
  XNOR2_X2 U624 ( .A(n767), .B(n524), .ZN(n661) );
  XNOR2_X1 U625 ( .A(KEYINPUT70), .B(G469), .ZN(n525) );
  XNOR2_X1 U626 ( .A(n527), .B(KEYINPUT96), .ZN(n531) );
  XOR2_X1 U627 ( .A(KEYINPUT5), .B(G113), .Z(n529) );
  XNOR2_X1 U628 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U629 ( .A(n531), .B(n530), .ZN(n535) );
  INV_X1 U630 ( .A(n591), .ZN(n701) );
  NOR2_X1 U631 ( .A1(n650), .A2(G902), .ZN(n542) );
  NAND2_X1 U632 ( .A1(G217), .A2(n538), .ZN(n540) );
  XOR2_X1 U633 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n539) );
  NAND2_X1 U634 ( .A1(n543), .A2(n697), .ZN(n544) );
  XNOR2_X1 U635 ( .A(n544), .B(KEYINPUT100), .ZN(n781) );
  INV_X1 U636 ( .A(n698), .ZN(n545) );
  INV_X1 U637 ( .A(n694), .ZN(n546) );
  XNOR2_X1 U638 ( .A(KEYINPUT101), .B(KEYINPUT33), .ZN(n547) );
  XNOR2_X2 U639 ( .A(n548), .B(n547), .ZN(n720) );
  XOR2_X1 U640 ( .A(KEYINPUT72), .B(KEYINPUT34), .Z(n551) );
  NOR2_X1 U641 ( .A1(n561), .A2(n562), .ZN(n599) );
  XNOR2_X1 U642 ( .A(KEYINPUT78), .B(n582), .ZN(n552) );
  AND2_X1 U643 ( .A1(n632), .A2(n697), .ZN(n554) );
  INV_X1 U644 ( .A(n780), .ZN(n555) );
  NOR2_X1 U645 ( .A1(n779), .A2(n555), .ZN(n556) );
  INV_X1 U646 ( .A(KEYINPUT44), .ZN(n557) );
  NAND2_X1 U647 ( .A1(n369), .A2(n559), .ZN(n560) );
  NOR2_X1 U648 ( .A1(n697), .A2(n560), .ZN(n668) );
  INV_X1 U649 ( .A(n561), .ZN(n563) );
  NAND2_X1 U650 ( .A1(n562), .A2(n563), .ZN(n580) );
  INV_X1 U651 ( .A(n580), .ZN(n680) );
  NOR2_X1 U652 ( .A1(n563), .A2(n562), .ZN(n682) );
  NOR2_X1 U653 ( .A1(n680), .A2(n682), .ZN(n715) );
  NOR2_X1 U654 ( .A1(n701), .A2(n564), .ZN(n705) );
  XNOR2_X1 U655 ( .A(n565), .B(KEYINPUT31), .ZN(n683) );
  NOR2_X1 U656 ( .A1(n591), .A2(n566), .ZN(n672) );
  NOR2_X1 U657 ( .A1(n683), .A2(n672), .ZN(n567) );
  NOR2_X1 U658 ( .A1(n715), .A2(n567), .ZN(n568) );
  NOR2_X1 U659 ( .A1(n668), .A2(n568), .ZN(n569) );
  NAND2_X1 U660 ( .A1(n570), .A2(n569), .ZN(n573) );
  INV_X1 U661 ( .A(KEYINPUT84), .ZN(n571) );
  INV_X1 U662 ( .A(KEYINPUT102), .ZN(n584) );
  NOR2_X1 U663 ( .A1(G900), .A2(n575), .ZN(n576) );
  NOR2_X1 U664 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U665 ( .A(KEYINPUT79), .B(n578), .Z(n597) );
  NOR2_X1 U666 ( .A1(n698), .A2(n597), .ZN(n579) );
  NOR2_X1 U667 ( .A1(n580), .A2(n601), .ZN(n581) );
  AND2_X1 U668 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U669 ( .A(n584), .B(n583), .ZN(n631) );
  BUF_X1 U670 ( .A(n585), .Z(n586) );
  NOR2_X1 U671 ( .A1(n631), .A2(n586), .ZN(n589) );
  NOR2_X1 U672 ( .A1(n452), .A2(n590), .ZN(n686) );
  NAND2_X1 U673 ( .A1(n591), .A2(n710), .ZN(n593) );
  XNOR2_X1 U674 ( .A(n593), .B(n592), .ZN(n595) );
  NAND2_X1 U675 ( .A1(n594), .A2(n595), .ZN(n596) );
  AND2_X1 U676 ( .A1(n395), .A2(n610), .ZN(n598) );
  NAND2_X1 U677 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U678 ( .A(KEYINPUT106), .B(n600), .ZN(n783) );
  BUF_X1 U679 ( .A(n604), .Z(n605) );
  INV_X1 U680 ( .A(n605), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n615), .A2(n606), .ZN(n619) );
  INV_X1 U682 ( .A(n619), .ZN(n678) );
  NAND2_X1 U683 ( .A1(n678), .A2(KEYINPUT81), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n783), .A2(n607), .ZN(n608) );
  NOR2_X1 U685 ( .A1(n686), .A2(n608), .ZN(n618) );
  INV_X1 U686 ( .A(n609), .ZN(n637) );
  XNOR2_X1 U687 ( .A(KEYINPUT38), .B(n637), .ZN(n711) );
  NAND2_X1 U688 ( .A1(n610), .A2(n711), .ZN(n612) );
  XOR2_X1 U689 ( .A(KEYINPUT71), .B(KEYINPUT39), .Z(n611) );
  XNOR2_X1 U690 ( .A(n612), .B(n611), .ZN(n639) );
  NAND2_X1 U691 ( .A1(n639), .A2(n680), .ZN(n614) );
  XOR2_X1 U692 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n613) );
  XNOR2_X1 U693 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n617) );
  NAND2_X1 U694 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U695 ( .A1(n615), .A2(n708), .ZN(n616) );
  NOR2_X1 U696 ( .A1(n620), .A2(KEYINPUT81), .ZN(n621) );
  NOR2_X1 U697 ( .A1(KEYINPUT47), .A2(n621), .ZN(n627) );
  INV_X1 U698 ( .A(KEYINPUT81), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n625) );
  INV_X1 U700 ( .A(n715), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U702 ( .A1(n627), .A2(n372), .ZN(n628) );
  NOR2_X1 U703 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n633), .A2(n710), .ZN(n636) );
  XOR2_X1 U705 ( .A(KEYINPUT43), .B(KEYINPUT103), .Z(n634) );
  XNOR2_X1 U706 ( .A(KEYINPUT104), .B(n634), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(n638) );
  NAND2_X1 U708 ( .A1(n638), .A2(n637), .ZN(n689) );
  NAND2_X1 U709 ( .A1(n682), .A2(n639), .ZN(n688) );
  NAND2_X1 U710 ( .A1(KEYINPUT2), .A2(n641), .ZN(n642) );
  NAND2_X1 U711 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U712 ( .A(n644), .B(KEYINPUT65), .ZN(n648) );
  BUF_X1 U713 ( .A(n645), .Z(n646) );
  NOR2_X1 U714 ( .A1(n646), .A2(n647), .ZN(n693) );
  NAND2_X1 U715 ( .A1(G217), .A2(n366), .ZN(n649) );
  XNOR2_X1 U716 ( .A(n650), .B(n649), .ZN(n651) );
  NOR2_X1 U717 ( .A1(n651), .A2(n754), .ZN(n653) );
  XNOR2_X1 U718 ( .A(n653), .B(n652), .ZN(G66) );
  INV_X1 U719 ( .A(KEYINPUT63), .ZN(n660) );
  NAND2_X1 U720 ( .A1(n366), .A2(G472), .ZN(n657) );
  XOR2_X1 U721 ( .A(KEYINPUT62), .B(KEYINPUT87), .Z(n656) );
  XNOR2_X1 U722 ( .A(n654), .B(KEYINPUT111), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n657), .B(n378), .ZN(n658) );
  NOR2_X1 U724 ( .A1(n658), .A2(n754), .ZN(n659) );
  XNOR2_X1 U725 ( .A(n659), .B(n660), .ZN(G57) );
  INV_X1 U726 ( .A(KEYINPUT121), .ZN(n667) );
  NAND2_X1 U727 ( .A1(n367), .A2(G469), .ZN(n664) );
  XNOR2_X1 U728 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n663) );
  XNOR2_X1 U729 ( .A(n661), .B(KEYINPUT57), .ZN(n662) );
  XNOR2_X1 U730 ( .A(n664), .B(n379), .ZN(n665) );
  NOR2_X1 U731 ( .A1(n665), .A2(n754), .ZN(n666) );
  XNOR2_X1 U732 ( .A(n666), .B(n667), .ZN(G54) );
  XOR2_X1 U733 ( .A(G101), .B(n668), .Z(G3) );
  NAND2_X1 U734 ( .A1(n672), .A2(n680), .ZN(n669) );
  XNOR2_X1 U735 ( .A(n669), .B(KEYINPUT112), .ZN(n670) );
  XNOR2_X1 U736 ( .A(n671), .B(n670), .ZN(G6) );
  XOR2_X1 U737 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n674) );
  NAND2_X1 U738 ( .A1(n672), .A2(n682), .ZN(n673) );
  XNOR2_X1 U739 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U740 ( .A(G107), .B(n675), .ZN(G9) );
  XOR2_X1 U741 ( .A(G128), .B(KEYINPUT29), .Z(n677) );
  NAND2_X1 U742 ( .A1(n678), .A2(n682), .ZN(n676) );
  XNOR2_X1 U743 ( .A(n677), .B(n676), .ZN(G30) );
  NAND2_X1 U744 ( .A1(n678), .A2(n680), .ZN(n679) );
  XNOR2_X1 U745 ( .A(n679), .B(G146), .ZN(G48) );
  NAND2_X1 U746 ( .A1(n683), .A2(n680), .ZN(n681) );
  XNOR2_X1 U747 ( .A(n681), .B(G113), .ZN(G15) );
  XOR2_X1 U748 ( .A(G116), .B(KEYINPUT113), .Z(n685) );
  NAND2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U750 ( .A(n685), .B(n684), .ZN(G18) );
  XNOR2_X1 U751 ( .A(G125), .B(n686), .ZN(n687) );
  XNOR2_X1 U752 ( .A(n687), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U753 ( .A(G134), .B(n688), .ZN(G36) );
  XNOR2_X1 U754 ( .A(G140), .B(n689), .ZN(G42) );
  INV_X1 U755 ( .A(n772), .ZN(n690) );
  NOR2_X1 U756 ( .A1(n690), .A2(n646), .ZN(n691) );
  NOR2_X1 U757 ( .A1(KEYINPUT2), .A2(n691), .ZN(n692) );
  NOR2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n731) );
  NAND2_X1 U759 ( .A1(n708), .A2(n353), .ZN(n729) );
  XOR2_X1 U760 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n696) );
  NAND2_X1 U761 ( .A1(n452), .A2(n694), .ZN(n695) );
  XNOR2_X1 U762 ( .A(n696), .B(n695), .ZN(n703) );
  NAND2_X1 U763 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U764 ( .A(KEYINPUT49), .B(n699), .Z(n700) );
  NAND2_X1 U765 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U767 ( .A1(n705), .A2(n704), .ZN(n707) );
  XOR2_X1 U768 ( .A(KEYINPUT51), .B(KEYINPUT115), .Z(n706) );
  XNOR2_X1 U769 ( .A(n707), .B(n706), .ZN(n709) );
  NAND2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n723) );
  NOR2_X1 U771 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U772 ( .A1(n713), .A2(n712), .ZN(n717) );
  NOR2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U774 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U775 ( .A(KEYINPUT116), .B(n718), .Z(n719) );
  NAND2_X1 U776 ( .A1(n353), .A2(n719), .ZN(n721) );
  XOR2_X1 U777 ( .A(KEYINPUT117), .B(n721), .Z(n722) );
  NAND2_X1 U778 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U779 ( .A(KEYINPUT52), .B(n724), .Z(n725) );
  NOR2_X1 U780 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U781 ( .A(KEYINPUT118), .B(n727), .Z(n728) );
  NAND2_X1 U782 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U783 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U784 ( .A1(n774), .A2(n732), .ZN(n733) );
  XNOR2_X1 U785 ( .A(n733), .B(KEYINPUT53), .ZN(n734) );
  XNOR2_X1 U786 ( .A(KEYINPUT119), .B(n734), .ZN(G75) );
  NAND2_X1 U787 ( .A1(n367), .A2(G210), .ZN(n739) );
  XNOR2_X1 U788 ( .A(KEYINPUT55), .B(KEYINPUT80), .ZN(n738) );
  BUF_X1 U789 ( .A(n735), .Z(n736) );
  XNOR2_X1 U790 ( .A(n736), .B(KEYINPUT54), .ZN(n737) );
  XNOR2_X1 U791 ( .A(n739), .B(n380), .ZN(n740) );
  NOR2_X1 U792 ( .A1(n740), .A2(n754), .ZN(n741) );
  XNOR2_X1 U793 ( .A(KEYINPUT56), .B(n741), .ZN(G51) );
  XOR2_X1 U794 ( .A(KEYINPUT59), .B(KEYINPUT88), .Z(n742) );
  XOR2_X1 U795 ( .A(KEYINPUT67), .B(KEYINPUT60), .Z(n747) );
  XNOR2_X1 U796 ( .A(n748), .B(n747), .ZN(G60) );
  XNOR2_X1 U797 ( .A(n749), .B(KEYINPUT122), .ZN(n752) );
  BUF_X1 U798 ( .A(n366), .Z(n750) );
  NAND2_X1 U799 ( .A1(G478), .A2(n750), .ZN(n751) );
  XNOR2_X1 U800 ( .A(n752), .B(n751), .ZN(n753) );
  NOR2_X1 U801 ( .A1(n754), .A2(n753), .ZN(G63) );
  NOR2_X1 U802 ( .A1(n404), .A2(n646), .ZN(n755) );
  XNOR2_X1 U803 ( .A(n755), .B(KEYINPUT125), .ZN(n760) );
  NAND2_X1 U804 ( .A1(n404), .A2(G224), .ZN(n756) );
  XNOR2_X1 U805 ( .A(KEYINPUT61), .B(n756), .ZN(n757) );
  NAND2_X1 U806 ( .A1(n757), .A2(G898), .ZN(n758) );
  XNOR2_X1 U807 ( .A(KEYINPUT124), .B(n758), .ZN(n759) );
  NAND2_X1 U808 ( .A1(n760), .A2(n759), .ZN(n766) );
  BUF_X1 U809 ( .A(n761), .Z(n762) );
  XNOR2_X1 U810 ( .A(n762), .B(G101), .ZN(n764) );
  NOR2_X1 U811 ( .A1(n774), .A2(G898), .ZN(n763) );
  NOR2_X1 U812 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U813 ( .A(n766), .B(n765), .ZN(G69) );
  XNOR2_X1 U814 ( .A(n768), .B(n767), .ZN(n773) );
  XOR2_X1 U815 ( .A(G227), .B(n773), .Z(n769) );
  NAND2_X1 U816 ( .A1(n769), .A2(G900), .ZN(n770) );
  NAND2_X1 U817 ( .A1(n770), .A2(n404), .ZN(n771) );
  XNOR2_X1 U818 ( .A(n771), .B(KEYINPUT126), .ZN(n777) );
  XNOR2_X1 U819 ( .A(n773), .B(n772), .ZN(n775) );
  NAND2_X1 U820 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U821 ( .A1(n777), .A2(n776), .ZN(G72) );
  XOR2_X1 U822 ( .A(G131), .B(n778), .Z(G33) );
  XOR2_X1 U823 ( .A(n368), .B(G122), .Z(G24) );
  XNOR2_X1 U824 ( .A(G119), .B(n780), .ZN(G21) );
  BUF_X1 U825 ( .A(n781), .Z(n782) );
  XNOR2_X1 U826 ( .A(G110), .B(n782), .ZN(G12) );
  XNOR2_X1 U827 ( .A(G143), .B(n783), .ZN(G45) );
  XOR2_X1 U828 ( .A(G137), .B(n784), .Z(G39) );
endmodule

