//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1284, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  NAND2_X1  g0001(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(KEYINPUT64), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G50), .ZN(new_n204));
  NOR2_X1   g0004(.A1(G58), .A2(G68), .ZN(new_n205));
  NAND3_X1  g0005(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0008(.A(G50), .B1(G58), .B2(G68), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT65), .Z(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n215), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n214), .B(new_n218), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n212), .A2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G159), .ZN(new_n246));
  OAI21_X1  g0046(.A(KEYINPUT77), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT77), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(new_n249), .A3(G159), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G68), .ZN(new_n252));
  AOI21_X1  g0052(.A(KEYINPUT76), .B1(new_n252), .B2(G20), .ZN(new_n253));
  AND2_X1   g0053(.A1(G58), .A2(G68), .ZN(new_n254));
  OAI211_X1 g0054(.A(KEYINPUT76), .B(G20), .C1(new_n254), .C2(new_n205), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n251), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT78), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(KEYINPUT7), .B1(new_n261), .B2(new_n212), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT7), .ZN(new_n263));
  NOR4_X1   g0063(.A1(new_n259), .A2(new_n260), .A3(new_n263), .A4(G20), .ZN(new_n264));
  OAI21_X1  g0064(.A(G68), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT78), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n266), .B(new_n251), .C1(new_n253), .C2(new_n256), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n258), .A2(KEYINPUT16), .A3(new_n265), .A4(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(G20), .B1(new_n254), .B2(new_n205), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT76), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n255), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n265), .A2(new_n272), .A3(new_n251), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT16), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT68), .B1(new_n215), .B2(new_n244), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT68), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n277), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(new_n211), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n268), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT8), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT8), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G58), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n281), .A2(G20), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT8), .B(G58), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n284), .A2(new_n291), .B1(new_n292), .B2(new_n283), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n280), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G87), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT79), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G1698), .ZN(new_n298));
  OAI211_X1 g0098(.A(G223), .B(new_n298), .C1(new_n259), .C2(new_n260), .ZN(new_n299));
  OAI211_X1 g0099(.A(G226), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT66), .B(G41), .ZN(new_n304));
  OAI211_X1 g0104(.A(KEYINPUT67), .B(new_n281), .C1(new_n304), .C2(G45), .ZN(new_n305));
  AND2_X1   g0105(.A1(KEYINPUT66), .A2(G41), .ZN(new_n306));
  NOR2_X1   g0106(.A1(KEYINPUT66), .A2(G41), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n281), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT67), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n281), .A2(G45), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G274), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n302), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n305), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G33), .A2(G41), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(G1), .A3(G13), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n281), .B1(G41), .B2(G45), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(G232), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT80), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT80), .A4(G232), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n303), .A2(new_n314), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G179), .ZN(new_n324));
  OR2_X1    g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(G169), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n294), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT18), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT18), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n294), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(G190), .B2(new_n323), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n280), .A2(new_n334), .A3(new_n293), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT17), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n280), .A2(new_n334), .A3(KEYINPUT17), .A4(new_n293), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n329), .A2(new_n331), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT81), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n244), .A2(G20), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G77), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n343), .A2(new_n344), .B1(new_n212), .B2(G68), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n245), .A2(new_n201), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n279), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT11), .ZN(new_n348));
  INV_X1    g0148(.A(G13), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(G1), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT69), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(G20), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n282), .A2(KEYINPUT69), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(new_n279), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(G68), .A3(new_n290), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT12), .ZN(new_n358));
  INV_X1    g0158(.A(G68), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n358), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  AND4_X1   g0160(.A1(new_n358), .A2(new_n350), .A3(G20), .A4(new_n359), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n348), .B(new_n357), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(G33), .A2(G97), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n229), .A2(G1698), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(G226), .B2(G1698), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n363), .B1(new_n365), .B2(new_n261), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n316), .A2(new_n317), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n366), .A2(new_n302), .B1(G238), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n369), .A3(new_n314), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n369), .B1(new_n368), .B2(new_n314), .ZN(new_n372));
  INV_X1    g0172(.A(G190), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n362), .A2(new_n374), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n305), .A2(new_n311), .A3(new_n313), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n316), .A2(G238), .A3(new_n317), .ZN(new_n377));
  INV_X1    g0177(.A(new_n363), .ZN(new_n378));
  NOR2_X1   g0178(.A1(G226), .A2(G1698), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n229), .B2(G1698), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT3), .B(G33), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n377), .B1(new_n382), .B2(new_n316), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT13), .B1(new_n376), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(KEYINPUT74), .A3(new_n370), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT74), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n368), .A2(new_n386), .A3(new_n369), .A4(new_n314), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(G200), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n375), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n356), .A2(G77), .A3(new_n290), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n289), .A2(new_n248), .B1(G20), .B2(G77), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT15), .B(G87), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n343), .B2(new_n392), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n393), .A2(new_n279), .B1(new_n344), .B2(new_n355), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G169), .ZN(new_n396));
  INV_X1    g0196(.A(G107), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n316), .B1(new_n261), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(G232), .A2(G1698), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n298), .A2(G238), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n381), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n398), .A2(new_n401), .B1(new_n367), .B2(G244), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n314), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n395), .B1(new_n396), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(G179), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT70), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G150), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n292), .A2(new_n343), .B1(new_n408), .B2(new_n245), .ZN(new_n409));
  XNOR2_X1  g0209(.A(KEYINPUT64), .B(G50), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n212), .B1(new_n410), .B2(new_n205), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n279), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n279), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n201), .B1(new_n281), .B2(G20), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n282), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n283), .A2(new_n201), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n412), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  OAI211_X1 g0218(.A(G222), .B(new_n298), .C1(new_n259), .C2(new_n260), .ZN(new_n419));
  OAI211_X1 g0219(.A(G223), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n419), .B(new_n420), .C1(new_n344), .C2(new_n381), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n302), .B1(G226), .B2(new_n367), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n314), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n418), .B1(new_n396), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(G179), .B2(new_n423), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n402), .A2(new_n314), .A3(G190), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n390), .A2(new_n394), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n403), .A2(G200), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n389), .A2(new_n407), .A3(new_n425), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT71), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT9), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(new_n417), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n417), .A2(new_n431), .A3(new_n432), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n332), .B1(new_n422), .B2(new_n314), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT73), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT10), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT72), .B1(new_n417), .B2(new_n432), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n289), .A2(new_n342), .B1(G150), .B2(new_n248), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n206), .A2(G20), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n443), .A2(new_n279), .B1(new_n201), .B2(new_n283), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT72), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT9), .A4(new_n415), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n422), .A2(G190), .A3(new_n314), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(new_n437), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n436), .A2(new_n439), .A3(new_n447), .A4(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n439), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n449), .ZN(new_n452));
  INV_X1    g0252(.A(new_n435), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n433), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n451), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n430), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n294), .A2(new_n327), .A3(new_n330), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n330), .B1(new_n294), .B2(new_n327), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n337), .A2(new_n338), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT81), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n371), .A2(new_n372), .A3(new_n324), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n385), .A2(G169), .A3(new_n387), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(KEYINPUT14), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT14), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n385), .A2(new_n465), .A3(G169), .A4(new_n387), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT75), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n466), .A2(new_n467), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n362), .ZN(new_n471));
  AND4_X1   g0271(.A1(new_n341), .A2(new_n456), .A3(new_n461), .A4(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G283), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT82), .B1(new_n244), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT82), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(G33), .A3(G283), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(G250), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n479));
  OAI211_X1 g0279(.A(G244), .B(new_n298), .C1(new_n259), .C2(new_n260), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT4), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n478), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n480), .A2(new_n481), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n302), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT5), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n281), .B(G45), .C1(new_n485), .C2(G41), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n485), .B1(new_n306), .B2(new_n307), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n302), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n486), .B1(new_n304), .B2(new_n485), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n489), .A2(G257), .B1(new_n490), .B2(new_n313), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n484), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G200), .ZN(new_n493));
  OAI21_X1  g0293(.A(G107), .B1(new_n262), .B2(new_n264), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT6), .ZN(new_n495));
  AND2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  NOR2_X1   g0296(.A1(G97), .A2(G107), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n397), .A2(KEYINPUT6), .A3(G97), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n500), .A2(G20), .B1(G77), .B2(new_n248), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G97), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n502), .A2(new_n279), .B1(new_n503), .B2(new_n283), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n284), .B(G97), .C1(G1), .C2(new_n244), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n484), .A2(new_n491), .A3(G190), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n493), .A2(new_n504), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n500), .A2(G20), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n248), .A2(G77), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n263), .B1(new_n381), .B2(G20), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n397), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n279), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n283), .A2(new_n503), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n505), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n492), .A2(new_n396), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n484), .A2(new_n491), .A3(new_n324), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n507), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(G238), .B(new_n298), .C1(new_n259), .C2(new_n260), .ZN(new_n521));
  OAI211_X1 g0321(.A(G244), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G116), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n302), .ZN(new_n525));
  INV_X1    g0325(.A(G250), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n302), .B1(new_n526), .B2(new_n310), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n281), .A2(new_n312), .A3(G45), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G200), .ZN(new_n531));
  AOI211_X1 g0331(.A(new_n283), .B(new_n279), .C1(new_n281), .C2(G33), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G87), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT19), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n342), .A2(new_n534), .A3(G97), .ZN(new_n535));
  INV_X1    g0335(.A(G87), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n497), .A2(new_n536), .B1(new_n363), .B2(new_n212), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n535), .B1(new_n537), .B2(new_n534), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n381), .A2(KEYINPUT84), .A3(new_n212), .A4(G68), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n212), .B(G68), .C1(new_n259), .C2(new_n260), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT84), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n543), .A2(new_n279), .B1(new_n355), .B2(new_n392), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n531), .A2(new_n533), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT85), .B1(new_n530), .B2(new_n373), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n524), .A2(new_n302), .B1(new_n527), .B2(new_n528), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT85), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n548), .A3(G190), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n547), .A2(KEYINPUT83), .A3(new_n324), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT83), .B1(new_n547), .B2(new_n324), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n392), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n284), .B(new_n554), .C1(G1), .C2(new_n244), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n544), .A2(new_n555), .B1(new_n396), .B2(new_n530), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n545), .A2(new_n550), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G257), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n558));
  OAI211_X1 g0358(.A(G250), .B(new_n298), .C1(new_n259), .C2(new_n260), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G294), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n302), .A2(new_n561), .B1(new_n489), .B2(G264), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n490), .A2(new_n313), .ZN(new_n563));
  AOI21_X1  g0363(.A(G169), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n302), .ZN(new_n565));
  OR2_X1    g0365(.A1(KEYINPUT66), .A2(G41), .ZN(new_n566));
  NAND2_X1  g0366(.A1(KEYINPUT66), .A2(G41), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT5), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G264), .B(new_n316), .C1(new_n568), .C2(new_n486), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n565), .A2(new_n563), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(G179), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n564), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n212), .B(G87), .C1(new_n259), .C2(new_n260), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT22), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT22), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n381), .A2(new_n575), .A3(new_n212), .A4(G87), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n212), .A2(KEYINPUT23), .A3(G107), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT23), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n578), .A2(KEYINPUT87), .B1(new_n579), .B2(new_n397), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n397), .A3(G20), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT87), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n583));
  OAI22_X1  g0383(.A1(new_n581), .A2(new_n582), .B1(new_n583), .B2(G20), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT24), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n577), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n586), .B1(new_n577), .B2(new_n585), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n279), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n283), .B(new_n397), .C1(KEYINPUT88), .C2(KEYINPUT25), .ZN(new_n590));
  NAND2_X1  g0390(.A1(KEYINPUT88), .A2(KEYINPUT25), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n532), .A2(G107), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n572), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n520), .A2(new_n557), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n562), .A2(new_n373), .A3(new_n563), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n570), .A2(new_n332), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n600), .A2(new_n589), .A3(new_n594), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT89), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT89), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n600), .A2(new_n603), .A3(new_n589), .A4(new_n594), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT21), .ZN(new_n606));
  INV_X1    g0406(.A(G116), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n355), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n607), .B1(new_n281), .B2(G33), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n413), .A2(new_n354), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(G20), .B1(new_n244), .B2(G97), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n478), .A2(new_n612), .B1(G20), .B2(new_n607), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT20), .B1(new_n613), .B2(new_n279), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(KEYINPUT20), .A3(new_n279), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n611), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(G264), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n618));
  OAI211_X1 g0418(.A(G257), .B(new_n298), .C1(new_n259), .C2(new_n260), .ZN(new_n619));
  XNOR2_X1  g0419(.A(KEYINPUT86), .B(G303), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n618), .B(new_n619), .C1(new_n381), .C2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n302), .ZN(new_n622));
  OAI211_X1 g0422(.A(G270), .B(new_n316), .C1(new_n568), .C2(new_n486), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(new_n563), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G169), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n606), .B1(new_n617), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n563), .A2(new_n623), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(G190), .A3(new_n622), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n624), .A2(G200), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n617), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n613), .A2(KEYINPUT20), .A3(new_n279), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n608), .B(new_n610), .C1(new_n632), .C2(new_n614), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n396), .B1(new_n628), .B2(new_n622), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT21), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n622), .A2(G179), .A3(new_n563), .A4(new_n623), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n626), .A2(new_n631), .A3(new_n635), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n605), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n473), .A2(new_n597), .A3(new_n640), .ZN(G372));
  INV_X1    g0441(.A(new_n425), .ZN(new_n642));
  INV_X1    g0442(.A(new_n389), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n471), .B1(new_n643), .B2(new_n407), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n460), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n459), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n455), .A2(KEYINPUT90), .A3(new_n450), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT90), .B1(new_n455), .B2(new_n450), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n642), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n507), .A2(new_n519), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n544), .A2(new_n555), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n530), .A2(new_n396), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n547), .A2(new_n324), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n547), .A2(new_n548), .A3(G190), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n548), .B1(new_n547), .B2(G190), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n531), .A2(new_n533), .A3(new_n544), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n651), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n596), .A2(new_n626), .A3(new_n638), .A4(new_n635), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n605), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n660), .B2(new_n519), .ZN(new_n665));
  INV_X1    g0465(.A(new_n519), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n545), .A2(new_n550), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n553), .A2(new_n556), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n666), .A2(new_n667), .A3(new_n668), .A4(KEYINPUT26), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n663), .A2(new_n670), .A3(new_n655), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n472), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n650), .A2(new_n672), .ZN(G369));
  NAND2_X1  g0473(.A1(new_n350), .A2(new_n212), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n633), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n639), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n626), .A2(new_n638), .A3(new_n635), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n681), .B1(new_n683), .B2(new_n680), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n595), .A2(new_n679), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n605), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n596), .ZN(new_n688));
  INV_X1    g0488(.A(new_n596), .ZN(new_n689));
  INV_X1    g0489(.A(new_n679), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n602), .A2(new_n604), .B1(new_n595), .B2(new_n679), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n694), .A2(new_n596), .A3(new_n682), .A4(new_n690), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n691), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n693), .A2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n304), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n216), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n281), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n497), .A2(new_n536), .A3(new_n607), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n701), .A2(new_n703), .B1(new_n210), .B2(new_n700), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  NAND2_X1  g0505(.A1(new_n671), .A2(new_n690), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(KEYINPUT29), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT26), .B1(new_n660), .B2(new_n519), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n557), .A2(new_n664), .A3(new_n666), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n663), .A2(new_n655), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n708), .B1(new_n711), .B2(new_n690), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n597), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(new_n605), .A3(new_n639), .A4(new_n690), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT91), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n565), .A2(new_n569), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n530), .B2(new_n717), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n484), .A2(new_n491), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n562), .A2(new_n547), .A3(KEYINPUT91), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n718), .A2(new_n637), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT30), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n492), .A2(new_n636), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(new_n720), .A4(new_n718), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT92), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n530), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n547), .A2(KEYINPUT92), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(new_n492), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n624), .A2(new_n324), .A3(new_n570), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n726), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT93), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n726), .B2(new_n733), .ZN(new_n737));
  AOI211_X1 g0537(.A(KEYINPUT93), .B(new_n732), .C1(new_n722), .C2(new_n725), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n737), .A2(new_n738), .A3(new_n690), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n715), .B(new_n735), .C1(new_n739), .C2(KEYINPUT31), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n713), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n705), .B1(new_n743), .B2(G1), .ZN(G364));
  NOR2_X1   g0544(.A1(new_n349), .A2(G20), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G45), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT95), .Z(new_n747));
  NAND2_X1  g0547(.A1(new_n701), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n381), .A2(new_n216), .ZN(new_n750));
  INV_X1    g0550(.A(G355), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n750), .A2(new_n751), .B1(G116), .B2(new_n216), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n239), .A2(G45), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n261), .A2(new_n216), .ZN(new_n754));
  INV_X1    g0554(.A(G45), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n754), .B1(new_n755), .B2(new_n210), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n752), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(G20), .B1(KEYINPUT96), .B2(G169), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(KEYINPUT96), .A2(G169), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n211), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n749), .B1(new_n757), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n212), .A2(G179), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(new_n373), .A3(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n474), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n212), .A2(new_n324), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(G190), .A3(new_n332), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G190), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n773), .A2(G322), .B1(new_n776), .B2(G329), .ZN(new_n777));
  INV_X1    g0577(.A(G311), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n771), .A2(new_n774), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n777), .B(new_n261), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n768), .A2(G190), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n770), .B(new_n780), .C1(G303), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n771), .A2(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n373), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G326), .ZN(new_n787));
  INV_X1    g0587(.A(G294), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n373), .A2(G179), .A3(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n212), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n786), .A2(new_n787), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n791), .A2(KEYINPUT98), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(KEYINPUT98), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n784), .A2(G190), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n794), .A2(KEYINPUT97), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(KEYINPUT97), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(G317), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n783), .A2(new_n792), .A3(new_n793), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n797), .A2(new_n359), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n775), .A2(new_n246), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT32), .ZN(new_n805));
  INV_X1    g0605(.A(new_n790), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n806), .A2(G97), .B1(new_n782), .B2(G87), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n381), .B1(new_n779), .B2(new_n344), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G58), .B2(new_n773), .ZN(new_n809));
  INV_X1    g0609(.A(new_n769), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n785), .A2(G50), .B1(new_n810), .B2(G107), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n805), .A2(new_n807), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n802), .B1(new_n803), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n767), .B1(new_n813), .B2(new_n761), .ZN(new_n814));
  INV_X1    g0614(.A(new_n764), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n684), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n684), .A2(G330), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT94), .Z(new_n818));
  NAND2_X1  g0618(.A1(new_n685), .A2(new_n748), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT100), .ZN(G396));
  AND3_X1   g0621(.A1(new_n404), .A2(new_n406), .A3(KEYINPUT101), .ZN(new_n822));
  AOI21_X1  g0622(.A(KEYINPUT101), .B1(new_n404), .B2(new_n406), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n429), .B1(new_n395), .B2(new_n690), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n671), .A2(new_n690), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n407), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n825), .B1(new_n828), .B2(new_n679), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n827), .B1(new_n706), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G330), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n640), .A2(new_n597), .A3(new_n679), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n734), .A2(KEYINPUT93), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n726), .A2(new_n736), .A3(new_n733), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n833), .A2(new_n679), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT31), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n832), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n831), .B1(new_n837), .B2(new_n735), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n830), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n830), .A2(new_n838), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n839), .A2(new_n748), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n761), .A2(new_n762), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(G77), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n798), .A2(G283), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n772), .A2(new_n788), .B1(new_n779), .B2(new_n607), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n381), .B(new_n846), .C1(G311), .C2(new_n776), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n806), .A2(G97), .B1(new_n782), .B2(G107), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n769), .A2(new_n536), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G303), .B2(new_n785), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n845), .A2(new_n847), .A3(new_n848), .A4(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n381), .B1(new_n775), .B2(new_n852), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n201), .A2(new_n781), .B1(new_n769), .B2(new_n359), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n853), .B(new_n854), .C1(G58), .C2(new_n806), .ZN(new_n855));
  INV_X1    g0655(.A(new_n779), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n773), .A2(G143), .B1(new_n856), .B2(G159), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n857), .B1(new_n858), .B2(new_n786), .C1(new_n797), .C2(new_n408), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n855), .B1(new_n860), .B2(KEYINPUT34), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT34), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n851), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n748), .B(new_n844), .C1(new_n864), .C2(new_n761), .ZN(new_n865));
  INV_X1    g0665(.A(new_n829), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n865), .B1(new_n866), .B2(new_n763), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n841), .A2(new_n867), .ZN(G384));
  NOR2_X1   g0668(.A1(new_n745), .A2(new_n281), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT105), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n471), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n470), .A2(KEYINPUT105), .A3(new_n362), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n362), .A2(new_n679), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n643), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n871), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n874), .B1(new_n470), .B2(new_n643), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n833), .A2(KEYINPUT31), .A3(new_n679), .A4(new_n834), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n879), .B(new_n715), .C1(new_n739), .C2(KEYINPUT31), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n878), .A2(new_n866), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT40), .ZN(new_n882));
  INV_X1    g0682(.A(new_n677), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n294), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n339), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n328), .A2(new_n884), .A3(new_n335), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n328), .A2(new_n884), .A3(new_n889), .A4(new_n335), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n267), .A2(new_n265), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n266), .B1(new_n272), .B2(new_n251), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n274), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(new_n279), .A3(new_n268), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n677), .B1(new_n898), .B2(new_n293), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n339), .A2(new_n899), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n280), .A2(new_n334), .A3(new_n293), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n898), .A2(new_n293), .B1(new_n326), .B2(new_n325), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n901), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n890), .B1(new_n903), .B2(new_n889), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n900), .A2(new_n904), .A3(KEYINPUT38), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n882), .B1(new_n894), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n829), .B1(new_n837), .B2(new_n879), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n901), .A2(new_n899), .ZN(new_n908));
  INV_X1    g0708(.A(new_n902), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n889), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n890), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n899), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n459), .B2(new_n460), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n893), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n905), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n907), .A2(new_n916), .A3(new_n878), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n881), .A2(new_n906), .B1(new_n917), .B2(new_n882), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT106), .Z(new_n919));
  NAND2_X1  g0719(.A1(new_n472), .A2(new_n880), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n831), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n919), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n690), .B1(new_n822), .B2(new_n823), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n876), .A2(new_n877), .B1(new_n826), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n459), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n925), .A2(new_n916), .B1(new_n926), .B2(new_n677), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT39), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n900), .A2(new_n904), .A3(KEYINPUT38), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n886), .B2(new_n891), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n915), .A2(KEYINPUT39), .A3(new_n905), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n470), .A2(KEYINPUT105), .A3(new_n362), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT105), .B1(new_n470), .B2(new_n362), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n690), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n931), .A2(new_n932), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n927), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n472), .B1(new_n712), .B2(new_n707), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n650), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n938), .B(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n869), .B1(new_n923), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n941), .B2(new_n923), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n209), .A2(new_n254), .A3(new_n344), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n944), .A2(KEYINPUT103), .B1(G68), .B2(new_n410), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(KEYINPUT103), .B2(new_n944), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(G1), .A3(new_n349), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT104), .Z(new_n948));
  INV_X1    g0748(.A(KEYINPUT102), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n950), .A2(G116), .A3(new_n213), .A4(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT36), .Z(new_n953));
  OAI21_X1  g0753(.A(new_n948), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n949), .B2(new_n953), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n943), .A2(new_n955), .ZN(G367));
  NAND2_X1  g0756(.A1(new_n516), .A2(new_n679), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n520), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n666), .A2(new_n679), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT107), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n693), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n962), .A2(new_n689), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n690), .B1(new_n964), .B2(new_n666), .ZN(new_n965));
  INV_X1    g0765(.A(new_n960), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n695), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT42), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n533), .A2(new_n544), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n679), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n667), .A2(new_n655), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n655), .B2(new_n971), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT43), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n965), .A2(new_n976), .A3(new_n968), .ZN(new_n977));
  XOR2_X1   g0777(.A(KEYINPUT108), .B(KEYINPUT109), .Z(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n975), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n979), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n963), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n977), .A2(new_n979), .ZN(new_n984));
  INV_X1    g0784(.A(new_n963), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n984), .A2(new_n985), .A3(new_n981), .A4(new_n975), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n747), .A2(G1), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT110), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n695), .A2(new_n691), .A3(new_n960), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT45), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT44), .B1(new_n696), .B2(new_n966), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT44), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n996), .B(new_n960), .C1(new_n695), .C2(new_n691), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n993), .A2(new_n994), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n693), .ZN(new_n999));
  INV_X1    g0799(.A(new_n693), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n995), .B2(new_n997), .C1(new_n994), .C2(new_n993), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n688), .A2(new_n691), .B1(new_n682), .B2(new_n690), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n695), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n685), .ZN(new_n1006));
  OAI211_X1 g0806(.A(G330), .B(new_n684), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1008), .A2(new_n713), .A3(new_n741), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n990), .B1(new_n1002), .B2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1011), .A2(new_n742), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1012), .A2(new_n999), .A3(KEYINPUT110), .A4(new_n1001), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n742), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n699), .B(KEYINPUT41), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n989), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n987), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n235), .A2(new_n754), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n765), .B1(new_n216), .B2(new_n392), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n749), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n781), .A2(new_n285), .B1(new_n775), .B2(new_n858), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n798), .A2(G159), .B1(KEYINPUT111), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(KEYINPUT111), .B2(new_n1021), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n381), .B1(new_n772), .B2(new_n408), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n410), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1024), .B1(new_n1025), .B2(new_n856), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n806), .A2(G68), .B1(new_n810), .B2(G77), .ZN(new_n1027));
  INV_X1    g0827(.A(G143), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1026), .B(new_n1027), .C1(new_n1028), .C2(new_n786), .ZN(new_n1029));
  INV_X1    g0829(.A(G317), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n779), .A2(new_n474), .B1(new_n775), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n261), .B1(new_n772), .B2(new_n620), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n781), .A2(new_n607), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1031), .B(new_n1032), .C1(KEYINPUT46), .C2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(KEYINPUT46), .B2(new_n1033), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n785), .A2(G311), .B1(new_n810), .B2(G97), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n397), .B2(new_n790), .C1(new_n797), .C2(new_n788), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1023), .A2(new_n1029), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT47), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1020), .B1(new_n1039), .B2(new_n761), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n973), .A2(new_n815), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1017), .A2(new_n1042), .ZN(G387));
  NAND2_X1  g0843(.A1(new_n1009), .A2(new_n700), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1044), .A2(KEYINPUT115), .B1(new_n742), .B2(new_n1011), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(KEYINPUT115), .B2(new_n1044), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n750), .A2(new_n703), .B1(G107), .B2(new_n216), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n232), .A2(G45), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT113), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n292), .A2(G50), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT50), .ZN(new_n1051));
  AOI211_X1 g0851(.A(G45), .B(new_n702), .C1(G68), .C2(G77), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n754), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1047), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n749), .B1(new_n1054), .B2(new_n766), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n761), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n785), .A2(G322), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n620), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n773), .A2(G317), .B1(new_n856), .B2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1057), .B(new_n1059), .C1(new_n797), .C2(new_n778), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n806), .A2(G283), .B1(new_n782), .B2(G294), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n261), .B1(new_n775), .B2(new_n787), .C1(new_n607), .C2(new_n769), .ZN(new_n1069));
  OR3_X1    g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n381), .B1(new_n775), .B2(new_n408), .C1(new_n359), .C2(new_n779), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n344), .A2(new_n781), .B1(new_n769), .B2(new_n503), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(G159), .C2(new_n785), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n790), .A2(new_n392), .B1(new_n772), .B2(new_n201), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT114), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1073), .B(new_n1075), .C1(new_n292), .C2(new_n797), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1056), .B1(new_n1070), .B2(new_n1076), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1055), .B(new_n1077), .C1(new_n692), .C2(new_n764), .ZN(new_n1078));
  OR3_X1    g0878(.A1(new_n1011), .A2(KEYINPUT112), .A3(new_n989), .ZN(new_n1079));
  OAI21_X1  g0879(.A(KEYINPUT112), .B1(new_n1011), .B2(new_n989), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1046), .A2(new_n1081), .ZN(G393));
  NAND2_X1  g0882(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT118), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1002), .A2(KEYINPUT118), .A3(new_n1009), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1087), .A2(new_n700), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT119), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n242), .A2(new_n754), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n765), .B1(new_n503), .B2(new_n216), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n749), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n781), .A2(new_n359), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n849), .B(new_n1095), .C1(G77), .C2(new_n806), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n381), .B1(new_n775), .B2(new_n1028), .C1(new_n292), .C2(new_n779), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1096), .B(new_n1098), .C1(new_n797), .C2(new_n410), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G150), .A2(new_n785), .B1(new_n773), .B2(G159), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT51), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n779), .A2(new_n788), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n381), .B(new_n1102), .C1(G322), .C2(new_n776), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n397), .A2(new_n769), .B1(new_n781), .B2(new_n474), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G116), .B2(new_n806), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(new_n797), .C2(new_n620), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G317), .A2(new_n785), .B1(new_n773), .B2(G311), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT52), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n1099), .A2(new_n1101), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1094), .B1(new_n1109), .B2(new_n761), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n962), .B2(new_n815), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT116), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n988), .B1(new_n1002), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(KEYINPUT116), .B1(new_n999), .B2(new_n1001), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1111), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT117), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g0917(.A(KEYINPUT117), .B(new_n1111), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1087), .A2(KEYINPUT119), .A3(new_n700), .A4(new_n1088), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1091), .A2(new_n1119), .A3(new_n1120), .ZN(G390));
  NAND2_X1  g0921(.A1(new_n826), .A2(new_n924), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n875), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n933), .A2(new_n934), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n877), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1122), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n935), .A2(new_n1126), .B1(new_n931), .B2(new_n932), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n740), .A2(G330), .A3(new_n866), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n933), .A2(new_n934), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1125), .B1(new_n1129), .B2(new_n875), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n711), .A2(new_n690), .A3(new_n825), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n876), .A2(new_n877), .B1(new_n1132), .B2(new_n924), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n935), .B1(new_n929), .B2(new_n930), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1127), .A2(new_n1131), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n907), .A2(G330), .A3(new_n878), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n915), .A2(KEYINPUT39), .A3(new_n905), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT39), .B1(new_n894), .B2(new_n905), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1138), .A2(new_n1139), .B1(new_n925), .B2(new_n936), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n894), .A2(new_n905), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1132), .A2(new_n924), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n935), .B(new_n1141), .C1(new_n1130), .C2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1137), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1136), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n472), .A2(G330), .A3(new_n880), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n650), .A2(new_n939), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n878), .B1(new_n838), .B2(new_n866), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n880), .A2(G330), .A3(new_n866), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1149), .A2(new_n1130), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1122), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n838), .A2(new_n866), .A3(new_n878), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1130), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(new_n1153), .A3(new_n1142), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1147), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n699), .B1(new_n1145), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1150), .B1(new_n1127), .B2(new_n1135), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1140), .A2(new_n1143), .A3(new_n1152), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1147), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1142), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n878), .B1(new_n907), .B2(G330), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1122), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1137), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1160), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT120), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1159), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1159), .B2(new_n1167), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1156), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n762), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n749), .B1(new_n289), .B2(new_n843), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n781), .A2(new_n408), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT53), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n261), .B1(new_n810), .B2(new_n1025), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1175), .B1(KEYINPUT121), .B2(new_n1176), .C1(new_n797), .C2(new_n858), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(KEYINPUT121), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G159), .A2(new_n806), .B1(new_n785), .B2(G128), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n773), .A2(G132), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT54), .B(G143), .Z(new_n1181));
  AOI22_X1  g0981(.A1(new_n856), .A2(new_n1181), .B1(new_n776), .B2(G125), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1182), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G77), .A2(new_n806), .B1(new_n785), .B2(G283), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n381), .B1(new_n776), .B2(G294), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n773), .A2(G116), .B1(new_n856), .B2(G97), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n782), .A2(G87), .B1(new_n810), .B2(G68), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n797), .A2(new_n397), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n1177), .A2(new_n1183), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1173), .B1(new_n1190), .B2(new_n761), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1145), .A2(new_n988), .B1(new_n1172), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1171), .A2(new_n1192), .ZN(G378));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1147), .B1(new_n1145), .B2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n418), .A2(new_n677), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n649), .B2(new_n425), .ZN(new_n1201));
  NOR4_X1   g1001(.A1(new_n647), .A2(new_n648), .A3(new_n642), .A4(new_n1199), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1198), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n649), .A2(new_n425), .A3(new_n1200), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n455), .A2(new_n450), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT90), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n455), .A2(KEYINPUT90), .A3(new_n450), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n425), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1199), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1204), .A2(new_n1210), .A3(new_n1197), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1203), .A2(KEYINPUT123), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n925), .A2(new_n916), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n926), .A2(new_n677), .ZN(new_n1214));
  AND4_X1   g1014(.A1(new_n937), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1212), .B1(new_n927), .B2(new_n937), .ZN(new_n1216));
  OAI211_X1 g1016(.A(G330), .B(new_n918), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1212), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n938), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n881), .A2(new_n906), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n917), .A2(new_n882), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1220), .A2(new_n1221), .A3(G330), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n927), .A2(new_n937), .A3(new_n1212), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1219), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1217), .A2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1194), .B1(new_n1196), .B2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1160), .B1(new_n1159), .B2(new_n1227), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1228), .A2(KEYINPUT57), .A3(new_n1217), .A4(new_n1224), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1226), .A2(new_n700), .A3(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1203), .A2(new_n762), .A3(new_n1211), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n749), .B1(new_n1025), .B2(new_n843), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n698), .B(new_n261), .C1(new_n781), .C2(new_n344), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n798), .A2(G97), .B1(KEYINPUT122), .B2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(KEYINPUT122), .B2(new_n1233), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n554), .A2(new_n856), .B1(new_n776), .B2(G283), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n397), .B2(new_n772), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G68), .A2(new_n806), .B1(new_n785), .B2(G116), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n285), .B2(new_n769), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1235), .A2(new_n1237), .A3(new_n1239), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1240), .B(KEYINPUT58), .Z(new_n1241));
  OAI221_X1 g1041(.A(new_n201), .B1(G33), .B2(G41), .C1(new_n381), .C2(new_n304), .ZN(new_n1242));
  INV_X1    g1042(.A(G128), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n772), .A2(new_n1243), .B1(new_n779), .B2(new_n858), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G150), .B2(new_n806), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n785), .A2(G125), .B1(new_n782), .B2(new_n1181), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(new_n797), .C2(new_n852), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(KEYINPUT59), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(KEYINPUT59), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n810), .A2(G159), .ZN(new_n1250));
  AOI211_X1 g1050(.A(G33), .B(G41), .C1(new_n776), .C2(G124), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1241), .B(new_n1242), .C1(new_n1248), .C2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1232), .B1(new_n1253), .B2(new_n761), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1231), .A2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1225), .B2(new_n989), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1230), .A2(new_n1257), .ZN(G375));
  NAND3_X1  g1058(.A1(new_n1151), .A2(new_n1147), .A3(new_n1154), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1015), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1167), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n381), .B1(new_n776), .B2(G303), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n1262), .B1(new_n397), .B2(new_n779), .C1(new_n474), .C2(new_n772), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n785), .A2(G294), .B1(new_n782), .B2(G97), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1264), .B1(new_n344), .B2(new_n769), .C1(new_n392), .C2(new_n790), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1263), .B(new_n1265), .C1(G116), .C2(new_n798), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(G150), .A2(new_n856), .B1(new_n776), .B2(G128), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1267), .B(new_n381), .C1(new_n858), .C2(new_n772), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n785), .A2(G132), .B1(new_n810), .B2(G58), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n1269), .B1(new_n201), .B2(new_n790), .C1(new_n246), .C2(new_n781), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1268), .B(new_n1270), .C1(new_n798), .C2(new_n1181), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n761), .B1(new_n1266), .B2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1272), .B(new_n749), .C1(G68), .C2(new_n843), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n1130), .B2(new_n762), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n1195), .B2(new_n988), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1261), .A2(new_n1275), .ZN(G381));
  AND2_X1   g1076(.A1(new_n1230), .A2(new_n1257), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n987), .A2(new_n1016), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1278));
  NOR4_X1   g1078(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(G390), .A2(G378), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .A4(new_n1280), .ZN(G407));
  INV_X1    g1081(.A(G378), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1277), .A2(G213), .A3(new_n678), .A4(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(G407), .A2(new_n1283), .A3(G213), .ZN(new_n1284));
  XOR2_X1   g1084(.A(new_n1284), .B(KEYINPUT124), .Z(G409));
  NAND3_X1  g1085(.A1(new_n1230), .A2(G378), .A3(new_n1257), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1196), .A2(new_n1225), .A3(new_n1015), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1171), .B(new_n1192), .C1(new_n1287), .C2(new_n1256), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n1286), .A2(new_n1288), .B1(G213), .B2(new_n678), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1151), .A2(KEYINPUT60), .A3(new_n1147), .A4(new_n1154), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1167), .A2(new_n1290), .A3(new_n700), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT60), .B1(new_n1227), .B2(new_n1147), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G384), .B(new_n1275), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT60), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1259), .A2(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1296), .A2(new_n700), .A3(new_n1167), .A4(new_n1290), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G384), .B1(new_n1297), .B2(new_n1275), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1294), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1289), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n678), .A2(G213), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1303), .B1(new_n1294), .B2(new_n1298), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n678), .A2(G213), .A3(G2897), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1275), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1306));
  INV_X1    g1106(.A(G384), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(KEYINPUT125), .A3(new_n1293), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1304), .A2(new_n1305), .A3(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1305), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1299), .A2(KEYINPUT125), .A3(new_n1311), .ZN(new_n1312));
  AOI22_X1  g1112(.A1(new_n1301), .A2(new_n1302), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT63), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1300), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  AND2_X1   g1115(.A1(G390), .A2(new_n1278), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(G390), .A2(new_n1278), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(G393), .A2(G396), .ZN(new_n1318));
  AND2_X1   g1118(.A1(G393), .A2(G396), .ZN(new_n1319));
  OAI22_X1  g1119(.A1(new_n1316), .A2(new_n1317), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT61), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(G387), .A2(new_n1322), .A3(new_n1091), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1319), .A2(new_n1318), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(G390), .A2(new_n1278), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1323), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1320), .A2(new_n1321), .A3(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT126), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1289), .A2(KEYINPUT63), .A3(new_n1299), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1320), .A2(KEYINPUT126), .A3(new_n1326), .A4(new_n1321), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1315), .A2(new_n1329), .A3(new_n1330), .A4(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1320), .A2(new_n1326), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT62), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1301), .A2(new_n1334), .A3(new_n1302), .A4(new_n1299), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1309), .A2(new_n1305), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1311), .B1(new_n1299), .B2(KEYINPUT125), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1336), .B1(new_n1337), .B2(new_n1304), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n1335), .B(new_n1321), .C1(new_n1289), .C2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1334), .B1(new_n1289), .B2(new_n1299), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1333), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1332), .A2(new_n1341), .ZN(G405));
  NAND2_X1  g1142(.A1(G375), .A2(new_n1282), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(new_n1286), .ZN(new_n1344));
  NOR3_X1   g1144(.A1(new_n1294), .A2(new_n1298), .A3(KEYINPUT127), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1345), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1343), .A2(new_n1286), .A3(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1346), .A2(new_n1348), .ZN(new_n1349));
  XNOR2_X1  g1149(.A(new_n1349), .B(new_n1333), .ZN(G402));
endmodule


