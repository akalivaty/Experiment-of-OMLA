//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n212), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n215), .B(new_n221), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT64), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n238), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT65), .ZN(new_n245));
  XOR2_X1   g0045(.A(G58), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n209), .A2(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G13), .ZN(new_n257));
  NOR3_X1   g0057(.A1(new_n257), .A2(new_n210), .A3(G1), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n219), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n256), .A2(new_n261), .B1(new_n258), .B2(new_n252), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G1), .A3(G13), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n267), .A3(G274), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n268), .B1(new_n270), .B2(new_n235), .ZN(new_n271));
  INV_X1    g0071(.A(G226), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G1698), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(G223), .B2(G1698), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  OAI22_X1  g0078(.A1(new_n274), .A2(new_n277), .B1(new_n278), .B2(new_n225), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n267), .B(KEYINPUT66), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n271), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G190), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(G200), .B2(new_n281), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT77), .ZN(new_n285));
  INV_X1    g0085(.A(new_n260), .ZN(new_n286));
  AOI21_X1  g0086(.A(KEYINPUT7), .B1(new_n277), .B2(new_n210), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT7), .ZN(new_n288));
  NOR4_X1   g0088(.A1(new_n275), .A2(new_n276), .A3(new_n288), .A4(G20), .ZN(new_n289));
  OAI21_X1  g0089(.A(G68), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G58), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(new_n223), .ZN(new_n292));
  OAI21_X1  g0092(.A(G20), .B1(new_n292), .B2(new_n201), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G159), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT16), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n286), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n290), .A2(KEYINPUT16), .A3(new_n297), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n285), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT3), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n278), .ZN(new_n304));
  NAND2_X1  g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n288), .B1(new_n306), .B2(G20), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n277), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n223), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n299), .B1(new_n309), .B2(new_n296), .ZN(new_n310));
  AND4_X1   g0110(.A1(new_n285), .A2(new_n310), .A3(new_n260), .A4(new_n301), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n262), .B(new_n284), .C1(new_n302), .C2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT17), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT18), .ZN(new_n314));
  INV_X1    g0114(.A(new_n262), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n310), .A2(new_n260), .A3(new_n301), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT77), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n310), .A2(new_n301), .A3(new_n285), .A4(new_n260), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT78), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n281), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  OR2_X1    g0122(.A1(new_n281), .A2(G169), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n320), .B1(new_n281), .B2(new_n321), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n314), .B1(new_n319), .B2(new_n325), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n319), .A2(new_n314), .A3(new_n325), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT79), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n262), .B1(new_n302), .B2(new_n311), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n323), .A2(new_n324), .ZN(new_n331));
  INV_X1    g0131(.A(new_n322), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(KEYINPUT18), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(KEYINPUT79), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n313), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n258), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(G68), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  OR3_X1    g0139(.A1(new_n339), .A2(KEYINPUT76), .A3(KEYINPUT12), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT76), .B1(new_n339), .B2(KEYINPUT12), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(KEYINPUT12), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n261), .A2(G68), .A3(new_n254), .ZN(new_n344));
  INV_X1    g0144(.A(new_n294), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n345), .A2(new_n202), .B1(new_n210), .B2(G68), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n210), .A2(G33), .ZN(new_n347));
  INV_X1    g0147(.A(G77), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n260), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT11), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n343), .A2(new_n344), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n268), .ZN(new_n353));
  INV_X1    g0153(.A(new_n270), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n353), .B1(G238), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(G232), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT72), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n306), .A2(KEYINPUT72), .A3(G232), .A4(G1698), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G97), .ZN(new_n360));
  INV_X1    g0160(.A(G1698), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n306), .A2(G226), .A3(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n358), .A2(new_n359), .A3(new_n360), .A4(new_n362), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n363), .A2(KEYINPUT73), .A3(new_n280), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT73), .B1(new_n363), .B2(new_n280), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n355), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT13), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT74), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(new_n355), .C1(new_n364), .C2(new_n365), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n367), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n366), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n352), .B1(new_n373), .B2(G200), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n367), .A2(G190), .A3(new_n370), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT75), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n375), .B(new_n376), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT70), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(KEYINPUT10), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n268), .B1(new_n270), .B2(new_n272), .ZN(new_n381));
  AOI21_X1  g0181(.A(G1698), .B1(new_n304), .B2(new_n305), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G222), .ZN(new_n383));
  INV_X1    g0183(.A(G223), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n306), .A2(G1698), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n383), .B1(new_n348), .B2(new_n306), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n381), .B1(new_n386), .B2(new_n280), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n387), .A2(G190), .ZN(new_n388));
  INV_X1    g0188(.A(G200), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n202), .B1(new_n209), .B2(G20), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n261), .A2(new_n393), .B1(new_n202), .B2(new_n258), .ZN(new_n394));
  INV_X1    g0194(.A(G150), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n252), .A2(new_n347), .B1(new_n395), .B2(new_n345), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(G20), .B2(new_n203), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n394), .B1(new_n397), .B2(new_n286), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT9), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT9), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n398), .A2(new_n401), .B1(new_n379), .B2(KEYINPUT10), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n380), .B1(new_n392), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n380), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n391), .A2(new_n405), .A3(new_n400), .A4(new_n402), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n387), .A2(new_n321), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(new_n398), .C1(G169), .C2(new_n387), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n353), .B1(G244), .B2(new_n354), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n385), .A2(new_n224), .B1(new_n206), .B2(new_n306), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n306), .A2(new_n361), .ZN(new_n412));
  OR3_X1    g0212(.A1(new_n412), .A2(KEYINPUT67), .A3(new_n235), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT67), .B1(new_n412), .B2(new_n235), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT66), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n267), .B(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n410), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G200), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT68), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n252), .B1(new_n420), .B2(new_n345), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n420), .B2(new_n345), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT15), .B(G87), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(new_n347), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(G20), .B2(G77), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n286), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n261), .A2(G77), .A3(new_n254), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n337), .A2(KEYINPUT69), .A3(G77), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT69), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n258), .B2(new_n348), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n427), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n419), .B(new_n432), .C1(new_n282), .C2(new_n418), .ZN(new_n433));
  INV_X1    g0233(.A(G169), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n432), .B1(new_n418), .B2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n321), .B(new_n410), .C1(new_n415), .C2(new_n417), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT71), .B1(new_n409), .B2(new_n438), .ZN(new_n439));
  OR3_X1    g0239(.A1(new_n409), .A2(KEYINPUT71), .A3(new_n438), .ZN(new_n440));
  AOI211_X1 g0240(.A(new_n336), .B(new_n378), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n371), .A2(G169), .A3(new_n372), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT14), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n371), .A2(KEYINPUT14), .A3(G169), .A4(new_n372), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n367), .A2(G179), .A3(new_n370), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n352), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n441), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT83), .ZN(new_n451));
  XNOR2_X1  g0251(.A(G97), .B(G107), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT6), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n453), .A2(new_n205), .A3(G107), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n457), .A2(G20), .B1(G77), .B2(new_n294), .ZN(new_n458));
  OAI21_X1  g0258(.A(G107), .B1(new_n287), .B2(new_n289), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n286), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n258), .A2(KEYINPUT80), .A3(new_n205), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(new_n337), .B2(G97), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n278), .A2(G1), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n258), .A2(new_n260), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n461), .B(new_n463), .C1(new_n466), .C2(new_n205), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n451), .B1(new_n460), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n467), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n455), .B1(new_n453), .B2(new_n452), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n470), .A2(new_n210), .B1(new_n348), .B2(new_n345), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n206), .B1(new_n307), .B2(new_n308), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n260), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(new_n473), .A3(KEYINPUT83), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  OAI211_X1 g0276(.A(G250), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n477));
  OAI211_X1 g0277(.A(G244), .B(new_n361), .C1(new_n275), .C2(new_n276), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT4), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n476), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT4), .B1(new_n382), .B2(G244), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n280), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n263), .A2(KEYINPUT5), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT82), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n483), .B(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n486));
  INV_X1    g0286(.A(G274), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n209), .B(G45), .C1(new_n263), .C2(KEYINPUT5), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n489), .A2(KEYINPUT81), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n489), .A2(KEYINPUT81), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n485), .B(new_n488), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n483), .ZN(new_n493));
  OAI211_X1 g0293(.A(G257), .B(new_n267), .C1(new_n493), .C2(new_n489), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n482), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G169), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n482), .A2(G179), .A3(new_n492), .A4(new_n494), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n475), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n460), .A2(new_n467), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n495), .A2(G200), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n500), .B(new_n501), .C1(new_n282), .C2(new_n495), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n306), .A2(G238), .A3(new_n361), .ZN(new_n503));
  OAI211_X1 g0303(.A(G244), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G116), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT84), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT84), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n503), .A2(new_n508), .A3(new_n504), .A4(new_n505), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n280), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n226), .B1(new_n264), .B2(G1), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n209), .A2(new_n487), .A3(G45), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n267), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n510), .A2(new_n321), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n306), .A2(new_n210), .A3(G68), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT19), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n210), .B1(new_n360), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(G87), .B2(new_n207), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n516), .B1(new_n347), .B2(new_n205), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n520), .A2(new_n260), .B1(new_n258), .B2(new_n423), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n423), .B2(new_n466), .ZN(new_n522));
  INV_X1    g0322(.A(new_n513), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n417), .B1(new_n506), .B2(KEYINPUT84), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n509), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n514), .B(new_n522), .C1(G169), .C2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n510), .A2(G190), .A3(new_n513), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n465), .A2(G87), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n527), .B(new_n529), .C1(new_n389), .C2(new_n525), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n499), .A2(new_n502), .A3(new_n526), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n465), .A2(G116), .ZN(new_n532));
  INV_X1    g0332(.A(G116), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n258), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(G20), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n260), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n476), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT20), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND4_X1   g0338(.A1(KEYINPUT20), .A2(new_n537), .A3(new_n260), .A4(new_n535), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n532), .B(new_n534), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(G264), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n541));
  OAI211_X1 g0341(.A(G257), .B(new_n361), .C1(new_n275), .C2(new_n276), .ZN(new_n542));
  INV_X1    g0342(.A(G303), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n541), .B(new_n542), .C1(new_n543), .C2(new_n306), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n280), .ZN(new_n545));
  OAI211_X1 g0345(.A(G270), .B(new_n267), .C1(new_n493), .C2(new_n489), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n492), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n540), .B1(new_n547), .B2(G200), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n282), .B2(new_n547), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n540), .A3(G169), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT21), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n547), .A2(new_n321), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n540), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n547), .A2(new_n540), .A3(KEYINPUT21), .A4(G169), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n549), .A2(new_n552), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(G264), .B(new_n267), .C1(new_n493), .C2(new_n489), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n492), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n382), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n306), .A2(G257), .A3(G1698), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n417), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n434), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G294), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n560), .B(new_n563), .C1(new_n412), .C2(new_n226), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n280), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n565), .A2(new_n321), .A3(new_n492), .A4(new_n557), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n306), .A2(new_n210), .A3(G87), .ZN(new_n568));
  XNOR2_X1  g0368(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n306), .A2(new_n569), .A3(new_n210), .A4(G87), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT24), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT23), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n210), .B2(G107), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n577));
  INV_X1    g0377(.A(new_n505), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n576), .A2(new_n577), .B1(new_n578), .B2(new_n210), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n573), .A2(new_n574), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n574), .B1(new_n573), .B2(new_n579), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n260), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT25), .B1(new_n258), .B2(new_n206), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n258), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n585), .A2(new_n586), .B1(new_n465), .B2(G107), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n567), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n558), .A2(new_n561), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G190), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n565), .A2(new_n492), .A3(new_n557), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G200), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n583), .A2(new_n591), .A3(new_n587), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  NOR4_X1   g0395(.A1(new_n450), .A2(new_n531), .A3(new_n556), .A4(new_n595), .ZN(G372));
  INV_X1    g0396(.A(new_n450), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n500), .B1(new_n496), .B2(new_n497), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT26), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n598), .A2(new_n526), .A3(new_n530), .A4(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n594), .B1(new_n588), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n600), .B1(new_n531), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n526), .A2(new_n530), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT26), .B1(new_n604), .B2(new_n499), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n526), .ZN(new_n606));
  OR2_X1    g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n597), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g0408(.A(new_n608), .B(KEYINPUT86), .Z(new_n609));
  INV_X1    g0409(.A(new_n352), .ZN(new_n610));
  INV_X1    g0410(.A(new_n447), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n444), .B2(new_n445), .ZN(new_n612));
  OAI22_X1  g0412(.A1(new_n378), .A2(new_n437), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n613), .A2(new_n313), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT18), .B1(new_n330), .B2(new_n333), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(new_n327), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n404), .B(new_n406), .C1(new_n614), .C2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n609), .A2(new_n408), .A3(new_n617), .ZN(G369));
  NAND3_X1  g0418(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n619), .A2(KEYINPUT27), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(KEYINPUT27), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(G213), .ZN(new_n622));
  INV_X1    g0422(.A(G343), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n540), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n601), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n556), .B2(new_n625), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(G330), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n624), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n583), .B2(new_n587), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n595), .A2(new_n632), .B1(new_n589), .B2(new_n631), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n601), .A2(new_n631), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n589), .A3(new_n594), .ZN(new_n638));
  XOR2_X1   g0438(.A(new_n624), .B(KEYINPUT87), .Z(new_n639));
  OAI21_X1  g0439(.A(new_n638), .B1(new_n589), .B2(new_n639), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n635), .A2(new_n640), .ZN(G399));
  INV_X1    g0441(.A(new_n213), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT88), .B1(new_n642), .B2(G41), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n642), .A2(KEYINPUT88), .A3(G41), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n225), .A2(new_n205), .A3(new_n206), .A4(new_n533), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n646), .A2(new_n209), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n218), .B2(new_n646), .ZN(new_n649));
  XOR2_X1   g0449(.A(new_n649), .B(KEYINPUT28), .Z(new_n650));
  INV_X1    g0450(.A(new_n639), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n607), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT29), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT90), .ZN(new_n655));
  OR3_X1    g0455(.A1(new_n531), .A2(new_n602), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n655), .B1(new_n531), .B2(new_n602), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n598), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT26), .B1(new_n604), .B2(new_n659), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n604), .A2(new_n499), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n526), .B(new_n660), .C1(new_n661), .C2(KEYINPUT26), .ZN(new_n662));
  OAI211_X1 g0462(.A(KEYINPUT29), .B(new_n631), .C1(new_n658), .C2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n654), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n595), .A2(new_n531), .A3(new_n556), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n651), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT31), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n547), .A2(new_n321), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(new_n495), .A3(new_n592), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n525), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n553), .A2(KEYINPUT89), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT89), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n547), .B2(new_n321), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n482), .A2(new_n494), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n525), .A2(new_n675), .A3(new_n590), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT30), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n676), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT30), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n678), .A2(new_n679), .A3(new_n673), .A4(new_n671), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n670), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n667), .B1(new_n681), .B2(new_n631), .ZN(new_n682));
  INV_X1    g0482(.A(new_n681), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n683), .A2(KEYINPUT31), .A3(new_n639), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n666), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n664), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT91), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n650), .B1(new_n688), .B2(G1), .ZN(G364));
  XOR2_X1   g0489(.A(new_n630), .B(KEYINPUT92), .Z(new_n690));
  INV_X1    g0490(.A(new_n646), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n257), .A2(G20), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n209), .B1(new_n692), .B2(G45), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n690), .B(new_n694), .C1(G330), .C2(new_n627), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n219), .B1(G20), .B2(new_n434), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n210), .A2(G179), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(G190), .A3(G200), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(new_n225), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n210), .A2(new_n321), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G200), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n282), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n699), .B1(G50), .B2(new_n702), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n282), .A2(G179), .A3(G200), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n210), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n697), .A2(new_n282), .A3(G200), .ZN(new_n706));
  OAI221_X1 g0506(.A(new_n703), .B1(new_n205), .B2(new_n705), .C1(new_n206), .C2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(G190), .A2(G200), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n697), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(G159), .ZN(new_n710));
  OAI21_X1  g0510(.A(KEYINPUT32), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OR3_X1    g0511(.A1(new_n709), .A2(KEYINPUT32), .A3(new_n710), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n701), .A2(G190), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n711), .B(new_n712), .C1(new_n714), .C2(new_n223), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n700), .A2(new_n708), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n700), .A2(G190), .A3(new_n389), .ZN(new_n717));
  OAI221_X1 g0517(.A(new_n306), .B1(new_n716), .B2(new_n348), .C1(new_n291), .C2(new_n717), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n707), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n698), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n702), .A2(G326), .B1(new_n720), .B2(G303), .ZN(new_n721));
  INV_X1    g0521(.A(G283), .ZN(new_n722));
  INV_X1    g0522(.A(G294), .ZN(new_n723));
  OAI221_X1 g0523(.A(new_n721), .B1(new_n722), .B2(new_n706), .C1(new_n723), .C2(new_n705), .ZN(new_n724));
  XNOR2_X1  g0524(.A(KEYINPUT33), .B(G317), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n713), .B1(new_n725), .B2(KEYINPUT94), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(KEYINPUT94), .B2(new_n725), .ZN(new_n727));
  INV_X1    g0527(.A(new_n717), .ZN(new_n728));
  INV_X1    g0528(.A(new_n709), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n728), .A2(G322), .B1(new_n729), .B2(G329), .ZN(new_n730));
  INV_X1    g0530(.A(G311), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n730), .B(new_n277), .C1(new_n731), .C2(new_n716), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n724), .A2(new_n727), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n696), .B1(new_n719), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n642), .A2(new_n277), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n735), .A2(G355), .B1(new_n533), .B2(new_n642), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n247), .A2(new_n264), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n642), .A2(new_n306), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(G45), .B2(new_n217), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n736), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n696), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT93), .Z(new_n745));
  AOI21_X1  g0545(.A(new_n694), .B1(new_n740), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n743), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n734), .B(new_n746), .C1(new_n627), .C2(new_n747), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n695), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(G396));
  INV_X1    g0550(.A(new_n716), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n728), .A2(G143), .B1(new_n751), .B2(G159), .ZN(new_n752));
  INV_X1    g0552(.A(new_n702), .ZN(new_n753));
  INV_X1    g0553(.A(G137), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n752), .B1(new_n753), .B2(new_n754), .C1(new_n395), .C2(new_n714), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT34), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  INV_X1    g0558(.A(G132), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n306), .B1(new_n709), .B2(new_n759), .C1(new_n705), .C2(new_n291), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n202), .A2(new_n698), .B1(new_n706), .B2(new_n223), .ZN(new_n761));
  NOR4_X1   g0561(.A1(new_n757), .A2(new_n758), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n713), .A2(G283), .B1(new_n751), .B2(G116), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT95), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n277), .B1(new_n709), .B2(new_n731), .C1(new_n717), .C2(new_n723), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n753), .A2(new_n543), .B1(new_n205), .B2(new_n705), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n225), .A2(new_n706), .B1(new_n698), .B2(new_n206), .ZN(new_n767));
  NOR4_X1   g0567(.A1(new_n764), .A2(new_n765), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n696), .B1(new_n762), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n694), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n696), .A2(new_n741), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n769), .B(new_n770), .C1(G77), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n418), .A2(new_n434), .ZN(new_n774));
  INV_X1    g0574(.A(new_n432), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n774), .A2(new_n436), .A3(new_n775), .A4(new_n624), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT96), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n435), .A2(KEYINPUT96), .A3(new_n436), .A4(new_n624), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n433), .B(new_n437), .C1(new_n432), .C2(new_n631), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n773), .B1(new_n783), .B2(new_n741), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n652), .A2(new_n783), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n782), .B(new_n651), .C1(new_n603), .C2(new_n606), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n770), .B1(new_n787), .B2(new_n686), .ZN(new_n788));
  INV_X1    g0588(.A(new_n686), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(new_n785), .A3(new_n786), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n784), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G384));
  NOR2_X1   g0592(.A1(new_n692), .A2(new_n209), .ZN(new_n793));
  INV_X1    g0593(.A(new_n622), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n330), .B1(new_n333), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT102), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n312), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n319), .A2(KEYINPUT102), .A3(new_n284), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n795), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(KEYINPUT37), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT103), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n799), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n803));
  AOI21_X1  g0603(.A(KEYINPUT37), .B1(new_n319), .B2(new_n284), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT104), .ZN(new_n805));
  AND3_X1   g0605(.A1(new_n795), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(new_n795), .B2(new_n804), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n802), .A2(new_n803), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT17), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n312), .B(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n330), .B(new_n794), .C1(new_n616), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT38), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT37), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n316), .A2(new_n262), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n794), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT100), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n319), .A2(new_n284), .B1(new_n333), .B2(new_n817), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n795), .A2(new_n804), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT38), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n819), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n336), .A2(KEYINPUT101), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(KEYINPUT101), .B1(new_n336), .B2(new_n825), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n815), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n683), .A2(KEYINPUT31), .A3(new_n624), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n666), .A2(new_n682), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n782), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT99), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n448), .A2(new_n833), .A3(new_n352), .ZN(new_n834));
  OAI21_X1  g0634(.A(KEYINPUT99), .B1(new_n612), .B2(new_n610), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n610), .A2(new_n631), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n374), .B2(new_n377), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n836), .B1(new_n378), .B2(new_n448), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n832), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n829), .A2(new_n840), .A3(KEYINPUT40), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT105), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT40), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n815), .B2(new_n828), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(KEYINPUT105), .A3(new_n840), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n821), .A2(new_n822), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT101), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n615), .B1(KEYINPUT79), .B2(new_n334), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n327), .A2(new_n328), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n811), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n849), .B1(new_n852), .B2(new_n819), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n336), .A2(KEYINPUT101), .A3(new_n825), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n848), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n828), .B1(new_n855), .B2(KEYINPUT38), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n840), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n844), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n847), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n597), .A2(new_n831), .ZN(new_n860));
  OAI21_X1  g0660(.A(G330), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n861), .A2(KEYINPUT106), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n861), .A2(KEYINPUT106), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n862), .B(new_n863), .C1(new_n859), .C2(new_n860), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n435), .A2(new_n436), .A3(new_n631), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n786), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT98), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT98), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n786), .A2(new_n869), .A3(new_n866), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n838), .A2(new_n839), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n856), .A2(new_n871), .B1(new_n616), .B2(new_n622), .ZN(new_n872));
  OAI211_X1 g0672(.A(KEYINPUT39), .B(new_n828), .C1(new_n855), .C2(KEYINPUT38), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n624), .B1(new_n834), .B2(new_n835), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT39), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n823), .B1(new_n853), .B2(new_n854), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT38), .B1(new_n809), .B2(new_n812), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n873), .A2(new_n874), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n872), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n441), .A2(new_n449), .A3(new_n654), .A4(new_n663), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n617), .A2(new_n408), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n880), .B(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n793), .B1(new_n865), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n883), .B2(new_n865), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n457), .A2(KEYINPUT35), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n457), .A2(KEYINPUT35), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n886), .A2(G116), .A3(new_n220), .A4(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT36), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n217), .A2(new_n348), .A3(new_n292), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n223), .A2(G50), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT97), .Z(new_n892));
  OAI211_X1 g0692(.A(G1), .B(new_n257), .C1(new_n890), .C2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n885), .A2(new_n889), .A3(new_n893), .ZN(G367));
  AND2_X1   g0694(.A1(new_n242), .A2(new_n738), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n744), .B1(new_n213), .B2(new_n423), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n770), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n717), .A2(new_n395), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n705), .A2(new_n223), .ZN(new_n899));
  AOI211_X1 g0699(.A(new_n898), .B(new_n899), .C1(G143), .C2(new_n702), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n901), .A2(KEYINPUT112), .ZN(new_n902));
  OAI221_X1 g0702(.A(new_n306), .B1(new_n709), .B2(new_n754), .C1(new_n202), .C2(new_n716), .ZN(new_n903));
  INV_X1    g0703(.A(new_n706), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(G77), .ZN(new_n905));
  OAI221_X1 g0705(.A(new_n905), .B1(new_n291), .B2(new_n698), .C1(new_n714), .C2(new_n710), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n902), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(KEYINPUT112), .B2(new_n901), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n698), .A2(new_n533), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n909), .A2(KEYINPUT46), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT110), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n277), .B1(new_n716), .B2(new_n722), .ZN(new_n912));
  XOR2_X1   g0712(.A(KEYINPUT111), .B(G317), .Z(new_n913));
  OAI22_X1  g0713(.A1(new_n717), .A2(new_n543), .B1(new_n913), .B2(new_n709), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n912), .B(new_n914), .C1(KEYINPUT46), .C2(new_n909), .ZN(new_n915));
  INV_X1    g0715(.A(new_n705), .ZN(new_n916));
  AOI22_X1  g0716(.A1(G107), .A2(new_n916), .B1(new_n702), .B2(G311), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n713), .A2(G294), .B1(new_n904), .B2(G97), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n911), .A2(new_n915), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n908), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT47), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n897), .B1(new_n921), .B2(new_n696), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n529), .A2(new_n631), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n526), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n526), .A2(new_n530), .A3(new_n923), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n922), .B1(new_n747), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n693), .B(KEYINPUT109), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n499), .B(new_n502), .C1(new_n651), .C2(new_n500), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT108), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n598), .B2(new_n639), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n640), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT44), .Z(new_n933));
  NOR2_X1   g0733(.A1(new_n931), .A2(new_n640), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT45), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n635), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n933), .A2(new_n634), .A3(new_n935), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n630), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n638), .B1(new_n633), .B2(new_n637), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n690), .B2(new_n941), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n688), .B1(new_n939), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n646), .B(KEYINPUT41), .Z(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n928), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n931), .A2(new_n638), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT42), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n499), .B1(new_n931), .B2(new_n589), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n651), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n926), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n954), .A2(KEYINPUT107), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(KEYINPUT107), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n955), .A2(new_n956), .A3(KEYINPUT43), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n957), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT43), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n960), .B2(new_n954), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n958), .B1(new_n953), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n931), .A2(new_n634), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n958), .B(new_n963), .C1(new_n953), .C2(new_n961), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n927), .B1(new_n948), .B2(new_n967), .ZN(G387));
  INV_X1    g0768(.A(new_n688), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n944), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n688), .A2(new_n943), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(new_n646), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n943), .A2(new_n928), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n735), .A2(new_n647), .B1(new_n206), .B2(new_n642), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n238), .A2(new_n264), .ZN(new_n975));
  AOI211_X1 g0775(.A(G45), .B(new_n647), .C1(G68), .C2(G77), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n253), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT50), .B1(new_n253), .B2(new_n202), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n738), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n974), .B1(new_n975), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n694), .B1(new_n981), .B2(new_n745), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n916), .A2(G283), .B1(new_n720), .B2(G294), .ZN(new_n983));
  INV_X1    g0783(.A(new_n913), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n728), .A2(new_n984), .B1(new_n751), .B2(G303), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n702), .A2(G322), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(new_n731), .C2(new_n714), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT48), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n983), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT114), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(new_n988), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(KEYINPUT49), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n306), .B1(new_n729), .B2(G326), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n533), .B2(new_n706), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n993), .B2(KEYINPUT49), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n705), .A2(new_n423), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n202), .B2(new_n717), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT113), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n714), .A2(new_n252), .B1(new_n706), .B2(new_n205), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n753), .A2(new_n710), .B1(new_n698), .B2(new_n348), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n306), .B1(new_n709), .B2(new_n395), .C1(new_n223), .C2(new_n716), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n994), .A2(new_n997), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n696), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n982), .B1(new_n633), .B2(new_n747), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n973), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n972), .A2(new_n1008), .ZN(G393));
  INV_X1    g0809(.A(new_n938), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n634), .B1(new_n933), .B2(new_n935), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n971), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n691), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n939), .A2(new_n971), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1012), .A2(new_n928), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n931), .A2(new_n743), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n738), .A2(new_n250), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n743), .B(new_n696), .C1(new_n642), .C2(G97), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n694), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n705), .A2(new_n533), .B1(new_n716), .B2(new_n723), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G317), .A2(new_n702), .B1(new_n728), .B2(G311), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT52), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1022), .B(new_n1024), .C1(G303), .C2(new_n713), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n306), .B1(new_n729), .B2(G322), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n206), .B2(new_n706), .C1(new_n722), .C2(new_n698), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT115), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n753), .A2(new_n395), .B1(new_n710), .B2(new_n717), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT51), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n714), .A2(new_n202), .B1(new_n706), .B2(new_n225), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n277), .B1(new_n729), .B2(G143), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n252), .B2(new_n716), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n705), .A2(new_n348), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n698), .A2(new_n223), .ZN(new_n1035));
  NOR4_X1   g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1025), .A2(new_n1028), .B1(new_n1030), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1018), .B(new_n1021), .C1(new_n1006), .C2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1016), .A2(new_n1017), .A3(new_n1038), .ZN(G390));
  NAND2_X1  g0839(.A1(new_n873), .A2(new_n878), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n741), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n713), .A2(G137), .B1(new_n904), .B2(G50), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n710), .B2(new_n705), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(KEYINPUT54), .B(G143), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n277), .B1(new_n751), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT53), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n698), .A2(new_n395), .ZN(new_n1048));
  INV_X1    g0848(.A(G125), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1046), .B1(new_n1047), .B2(new_n1048), .C1(new_n1049), .C2(new_n709), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1043), .B(new_n1050), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G128), .A2(new_n702), .B1(new_n728), .B2(G132), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT118), .Z(new_n1053));
  OAI22_X1  g0853(.A1(new_n706), .A2(new_n223), .B1(new_n709), .B2(new_n723), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT119), .Z(new_n1055));
  OAI22_X1  g0855(.A1(new_n206), .A2(new_n714), .B1(new_n753), .B2(new_n722), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n277), .B1(new_n716), .B2(new_n205), .C1(new_n533), .C2(new_n717), .ZN(new_n1057));
  NOR4_X1   g0857(.A1(new_n1056), .A2(new_n699), .A3(new_n1034), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1051), .A2(new_n1053), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n770), .B1(new_n253), .B2(new_n772), .C1(new_n1059), .C2(new_n1006), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT120), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1041), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n838), .A2(new_n839), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n868), .A2(new_n870), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n834), .A2(new_n835), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n631), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1040), .A2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n631), .B(new_n782), .C1(new_n658), .C2(new_n662), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n838), .A2(new_n839), .B1(new_n1070), .B2(new_n866), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n874), .B1(new_n815), .B2(new_n828), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n686), .A2(new_n783), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1072), .A2(new_n1073), .B1(new_n1063), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1069), .A2(KEYINPUT116), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT116), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n873), .A2(new_n878), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1074), .A2(new_n1063), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1067), .B1(new_n876), .B2(new_n877), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n1080), .B2(new_n1071), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1077), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1076), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n832), .A2(new_n629), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1084), .A2(new_n1063), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1080), .A2(new_n1071), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1085), .B1(new_n1078), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n928), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1062), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n441), .A2(G330), .A3(new_n449), .A4(new_n831), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n617), .A2(new_n408), .A3(new_n881), .A4(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1074), .A2(new_n1063), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1064), .B1(new_n1085), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1070), .A2(new_n866), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1079), .B(new_n1097), .C1(new_n1063), .C2(new_n1084), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1093), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT116), .B1(new_n1069), .B2(new_n1075), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n1078), .A2(new_n1081), .A3(new_n1077), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1099), .B(new_n1087), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT117), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n1103), .A3(new_n646), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1093), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1088), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1103), .B1(new_n1102), .B2(new_n646), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1091), .B1(new_n1109), .B2(new_n1110), .ZN(G378));
  XNOR2_X1  g0911(.A(new_n1093), .B(KEYINPUT123), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1102), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n629), .B1(new_n857), .B2(new_n844), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n847), .A2(new_n880), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n880), .B1(new_n847), .B2(new_n1114), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n399), .A2(new_n622), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n409), .B(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1118), .B(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1115), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n880), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n845), .A2(KEYINPUT105), .A3(new_n840), .ZN(new_n1124));
  AOI21_X1  g0924(.A(KEYINPUT105), .B1(new_n845), .B2(new_n840), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n858), .A2(G330), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1123), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n847), .A2(new_n880), .A3(new_n1114), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1120), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1113), .B(KEYINPUT57), .C1(new_n1122), .C2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1121), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1128), .A2(new_n1120), .A3(new_n1129), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1132), .A2(new_n1133), .B1(new_n1102), .B2(new_n1112), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1131), .B(new_n646), .C1(new_n1134), .C2(KEYINPUT57), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1121), .A2(new_n742), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n899), .B1(G116), .B2(new_n702), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT122), .Z(new_n1138));
  NOR2_X1   g0938(.A1(new_n706), .A2(new_n291), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT121), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n714), .A2(new_n205), .B1(new_n698), .B2(new_n348), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n277), .A2(new_n263), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n717), .A2(new_n206), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n716), .A2(new_n423), .B1(new_n709), .B2(new_n722), .ZN(new_n1144));
  NOR4_X1   g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1138), .A2(new_n1140), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(KEYINPUT58), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1142), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n1049), .A2(new_n753), .B1(new_n714), .B2(new_n759), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n728), .A2(G128), .B1(new_n751), .B2(G137), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n698), .B2(new_n1044), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(G150), .C2(new_n916), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n904), .A2(G159), .ZN(new_n1158));
  AOI211_X1 g0958(.A(G33), .B(G41), .C1(new_n729), .C2(G124), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1150), .B1(KEYINPUT58), .B2(new_n1147), .C1(new_n1156), .C2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n696), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1162), .B(new_n770), .C1(G50), .C2(new_n772), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1136), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n928), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1135), .A2(new_n1166), .ZN(G375));
  INV_X1    g0967(.A(new_n1105), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n1093), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1169), .A2(new_n947), .A3(new_n1107), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n838), .A2(new_n741), .A3(new_n839), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n770), .B1(G68), .B2(new_n772), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n533), .A2(new_n714), .B1(new_n753), .B2(new_n723), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G97), .B2(new_n720), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n717), .A2(new_n722), .B1(new_n716), .B2(new_n206), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n306), .B(new_n1175), .C1(G303), .C2(new_n729), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1174), .A2(new_n905), .A3(new_n998), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1140), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G132), .A2(new_n702), .B1(new_n713), .B2(new_n1045), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n277), .B1(new_n728), .B2(G137), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G150), .A2(new_n751), .B1(new_n729), .B2(G128), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n916), .A2(G50), .B1(new_n720), .B2(G159), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1177), .B1(new_n1178), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1172), .B1(new_n1184), .B2(new_n696), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1105), .A2(new_n928), .B1(new_n1171), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1170), .A2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT124), .ZN(G381));
  NAND3_X1  g0988(.A1(new_n972), .A2(new_n749), .A3(new_n1008), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(G384), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1190), .A2(KEYINPUT125), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(KEYINPUT125), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n969), .B1(new_n1012), .B2(new_n943), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1089), .B1(new_n1193), .B2(new_n946), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n965), .A2(new_n966), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1017), .A2(new_n1038), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1198), .A3(new_n927), .ZN(new_n1199));
  OR3_X1    g0999(.A1(new_n1191), .A2(new_n1192), .A3(new_n1199), .ZN(new_n1200));
  OR4_X1    g1000(.A1(G378), .A2(new_n1200), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1001(.A(G378), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n623), .A2(G213), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  OAI211_X1 g1005(.A(G407), .B(G213), .C1(G375), .C2(new_n1205), .ZN(G409));
  NAND2_X1  g1006(.A1(new_n1131), .A2(new_n646), .ZN(new_n1207));
  AOI21_X1  g1007(.A(KEYINPUT57), .B1(new_n1165), .B2(new_n1113), .ZN(new_n1208));
  OAI211_X1 g1008(.A(G378), .B(new_n1166), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1113), .B(new_n947), .C1(new_n1122), .C2(new_n1130), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n928), .B1(new_n1122), .B2(new_n1130), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1164), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1110), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1213), .A2(new_n1216), .A3(new_n1091), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1209), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1107), .A2(KEYINPUT60), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1169), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1168), .A2(KEYINPUT60), .A3(new_n1093), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1220), .A2(new_n646), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1186), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n791), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1220), .A2(new_n646), .A3(new_n1221), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1225), .A2(G384), .A3(new_n1186), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1218), .A2(new_n1203), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT62), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1218), .A2(new_n1203), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1204), .A2(G2897), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1227), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1224), .A2(new_n1226), .A3(new_n1232), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1231), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT61), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1204), .B1(new_n1209), .B2(new_n1217), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT62), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1240), .A3(new_n1228), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1230), .A2(new_n1237), .A3(new_n1238), .A4(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G387), .A2(G390), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G393), .A2(G396), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1189), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1199), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1199), .B2(new_n1243), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1242), .A2(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1250), .B(new_n1238), .C1(new_n1239), .C2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT126), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1204), .B(new_n1227), .C1(new_n1209), .C2(new_n1217), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1254), .B1(new_n1255), .B2(KEYINPUT63), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(KEYINPUT63), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT63), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1229), .A2(KEYINPUT126), .A3(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1253), .A2(new_n1256), .A3(new_n1257), .A4(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1249), .A2(new_n1260), .ZN(G405));
  INV_X1    g1061(.A(new_n1209), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G378), .B1(new_n1135), .B2(new_n1166), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1228), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G375), .A2(new_n1202), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(new_n1209), .A3(new_n1227), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1248), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1248), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT127), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1267), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  AOI211_X1 g1070(.A(KEYINPUT127), .B(new_n1248), .C1(new_n1264), .C2(new_n1266), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(G402));
endmodule


