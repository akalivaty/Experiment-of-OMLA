//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943;
  XOR2_X1   g000(.A(G43gat), .B(G50gat), .Z(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT89), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT15), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT15), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n202), .A2(KEYINPUT89), .A3(new_n205), .ZN(new_n206));
  OR3_X1    g005(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n207), .A2(new_n208), .B1(G29gat), .B2(G36gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n204), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT90), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  OR3_X1    g011(.A1(new_n209), .A2(new_n205), .A3(new_n202), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT17), .ZN(new_n215));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216));
  INV_X1    g015(.A(G85gat), .ZN(new_n217));
  INV_X1    g016(.A(G92gat), .ZN(new_n218));
  AOI22_X1  g017(.A1(KEYINPUT8), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(new_n217), .B2(new_n218), .ZN(new_n221));
  NAND4_X1  g020(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G99gat), .B(G106gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n219), .A2(new_n224), .A3(new_n221), .A4(new_n222), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XOR2_X1   g027(.A(new_n228), .B(KEYINPUT99), .Z(new_n229));
  NAND2_X1  g028(.A1(new_n215), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n229), .ZN(new_n231));
  AND2_X1   g030(.A1(G232gat), .A2(G233gat), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n214), .A2(new_n231), .B1(KEYINPUT41), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(G190gat), .B(G218gat), .Z(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n232), .A2(KEYINPUT41), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(G134gat), .B(G162gat), .Z(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n237), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n236), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n239), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G57gat), .ZN(new_n246));
  OR2_X1    g045(.A1(KEYINPUT95), .A2(G64gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(KEYINPUT95), .A2(G64gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT96), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT96), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(new_n246), .B2(G64gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n250), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(G71gat), .A2(G78gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT9), .ZN(new_n255));
  NAND2_X1  g054(.A1(G71gat), .A2(G78gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(G57gat), .B(G64gat), .Z(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT9), .ZN(new_n260));
  INV_X1    g059(.A(new_n256), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(new_n254), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(G231gat), .A2(G233gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G127gat), .B(G155gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n270), .B(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G8gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(G15gat), .B(G22gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT91), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G1gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT16), .ZN(new_n279));
  XOR2_X1   g078(.A(new_n279), .B(KEYINPUT92), .Z(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n274), .B1(new_n281), .B2(KEYINPUT93), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n281), .B1(G1gat), .B2(new_n277), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI221_X1 g083(.A(new_n281), .B1(KEYINPUT93), .B2(new_n274), .C1(G1gat), .C2(new_n277), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n253), .A2(new_n257), .B1(new_n260), .B2(new_n262), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n286), .B1(KEYINPUT21), .B2(new_n287), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n273), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n288), .ZN(new_n290));
  XOR2_X1   g089(.A(G183gat), .B(G211gat), .Z(new_n291));
  OR3_X1    g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n289), .B2(new_n290), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n245), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n228), .B1(new_n258), .B2(new_n263), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n227), .A2(KEYINPUT100), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n226), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n223), .A2(KEYINPUT100), .A3(new_n225), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n296), .B1(new_n287), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G230gat), .A2(G233gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n304), .B(KEYINPUT102), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT10), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n229), .A2(new_n306), .A3(new_n264), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT101), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n301), .B2(KEYINPUT10), .ZN(new_n309));
  INV_X1    g108(.A(new_n228), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n264), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n300), .A2(new_n287), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(KEYINPUT101), .A3(new_n306), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n307), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n302), .B(KEYINPUT103), .Z(new_n316));
  OAI21_X1  g115(.A(new_n305), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G120gat), .B(G148gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(G176gat), .B(G204gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n320), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n305), .B(new_n322), .C1(new_n303), .C2(new_n315), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n295), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n214), .A2(new_n286), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT94), .ZN(new_n327));
  INV_X1    g126(.A(new_n286), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n215), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G229gat), .A2(G233gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(KEYINPUT18), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n327), .A2(new_n329), .A3(new_n331), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT18), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n327), .B1(new_n214), .B2(new_n286), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n331), .B(KEYINPUT13), .Z(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n332), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G113gat), .B(G141gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT11), .ZN(new_n341));
  INV_X1    g140(.A(G169gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n343), .B(G197gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n344), .B(KEYINPUT12), .Z(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n345), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n332), .A2(new_n335), .A3(new_n338), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(KEYINPUT31), .B(G50gat), .Z(new_n351));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352));
  XNOR2_X1  g151(.A(G211gat), .B(G218gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n354));
  XNOR2_X1  g153(.A(G197gat), .B(G204gat), .ZN(new_n355));
  INV_X1    g154(.A(G211gat), .ZN(new_n356));
  INV_X1    g155(.A(G218gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT74), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G218gat), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n356), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n354), .B(new_n355), .C1(new_n361), .C2(KEYINPUT22), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT22), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT74), .B(G218gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n364), .B1(new_n365), .B2(new_n356), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n354), .B1(new_n366), .B2(new_n355), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n353), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n358), .A2(new_n360), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT22), .B1(new_n369), .B2(G211gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n355), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT75), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n353), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n362), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT29), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(KEYINPUT86), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT86), .ZN(new_n377));
  AOI211_X1 g176(.A(new_n377), .B(KEYINPUT29), .C1(new_n368), .C2(new_n374), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n352), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G155gat), .ZN(new_n380));
  INV_X1    g179(.A(G162gat), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT2), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G141gat), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n383), .A2(G148gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(G148gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n382), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G155gat), .B(G162gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(G155gat), .A2(G162gat), .ZN(new_n388));
  OR2_X1    g187(.A1(new_n388), .A2(KEYINPUT79), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n387), .B1(new_n386), .B2(new_n389), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n379), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(G228gat), .ZN(new_n395));
  INV_X1    g194(.A(G233gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n368), .A2(new_n374), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n352), .B1(new_n391), .B2(new_n392), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT29), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n398), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n394), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT85), .ZN(new_n406));
  XNOR2_X1  g205(.A(G141gat), .B(G148gat), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT2), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n408), .B1(G155gat), .B2(G162gat), .ZN(new_n409));
  OAI22_X1  g208(.A1(new_n407), .A2(new_n409), .B1(KEYINPUT79), .B2(new_n388), .ZN(new_n410));
  INV_X1    g209(.A(new_n387), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n390), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT29), .B1(new_n413), .B2(new_n352), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT84), .B1(new_n399), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n403), .A2(new_n416), .A3(new_n374), .A4(new_n368), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n393), .B1(new_n375), .B2(KEYINPUT3), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n406), .B1(new_n420), .B2(new_n398), .ZN(new_n421));
  AOI211_X1 g220(.A(KEYINPUT85), .B(new_n397), .C1(new_n418), .C2(new_n419), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n405), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(G22gat), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n372), .A2(new_n362), .A3(new_n373), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n373), .B1(new_n372), .B2(new_n362), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n402), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n352), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n393), .A2(new_n428), .B1(new_n415), .B2(new_n417), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT85), .B1(new_n429), .B2(new_n397), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n420), .A2(new_n406), .A3(new_n398), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(G22gat), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n405), .ZN(new_n434));
  XNOR2_X1  g233(.A(G78gat), .B(G106gat), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n424), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n424), .B2(new_n434), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n351), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  XOR2_X1   g237(.A(G127gat), .B(G134gat), .Z(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT69), .ZN(new_n440));
  XNOR2_X1  g239(.A(G127gat), .B(G134gat), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT69), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT68), .ZN(new_n444));
  INV_X1    g243(.A(G120gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(G113gat), .ZN(new_n446));
  INV_X1    g245(.A(G113gat), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT68), .B1(new_n447), .B2(G120gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(G120gat), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT1), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n440), .A2(new_n443), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G113gat), .B(G120gat), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n439), .B1(new_n453), .B2(KEYINPUT1), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n393), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n413), .A2(new_n454), .A3(new_n452), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G225gat), .A2(G233gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT80), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT5), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n393), .A2(new_n455), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n460), .B1(new_n463), .B2(KEYINPUT4), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT82), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n412), .A2(KEYINPUT3), .A3(new_n390), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n401), .A2(new_n455), .A3(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n468));
  NAND2_X1  g267(.A1(new_n457), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n464), .A2(new_n465), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n467), .ZN(new_n471));
  INV_X1    g270(.A(new_n460), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT4), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n472), .B1(new_n457), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT82), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n462), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n467), .B1(new_n457), .B2(new_n468), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n463), .A2(KEYINPUT4), .ZN(new_n478));
  NOR4_X1   g277(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT5), .A4(new_n460), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  XOR2_X1   g279(.A(G1gat), .B(G29gat), .Z(new_n481));
  XNOR2_X1  g280(.A(G57gat), .B(G85gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n484));
  XOR2_X1   g283(.A(new_n483), .B(new_n484), .Z(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n485), .B1(new_n476), .B2(new_n479), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n489), .A2(new_n488), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G226gat), .A2(G233gat), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n493), .B(KEYINPUT76), .Z(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT23), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(G169gat), .B2(G176gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT65), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(KEYINPUT67), .B(G190gat), .Z(new_n501));
  INV_X1    g300(.A(G183gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G183gat), .A2(G190gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT24), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n500), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G169gat), .A2(G176gat), .ZN(new_n507));
  INV_X1    g306(.A(G176gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n342), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n507), .B1(new_n509), .B2(new_n497), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT66), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n496), .B1(new_n506), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(G169gat), .A2(G176gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT26), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n507), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G183gat), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n501), .A2(KEYINPUT28), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT28), .B1(new_n501), .B2(new_n517), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n504), .B(new_n516), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n505), .B1(G183gat), .B2(G190gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n498), .B(KEYINPUT65), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT64), .B(G169gat), .Z(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(KEYINPUT23), .A3(new_n508), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT25), .B1(G169gat), .B2(G176gat), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n521), .A2(new_n522), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n513), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n495), .B1(new_n528), .B2(KEYINPUT29), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT77), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n528), .B2(new_n495), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n503), .A2(new_n505), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n512), .A2(new_n522), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT25), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(new_n520), .A3(new_n526), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(KEYINPUT77), .A3(new_n494), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n529), .A2(new_n531), .A3(new_n536), .A4(new_n399), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n494), .B1(new_n535), .B2(new_n402), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n528), .A2(new_n495), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n400), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G8gat), .B(G36gat), .Z(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT78), .ZN(new_n542));
  XOR2_X1   g341(.A(G64gat), .B(G92gat), .Z(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n537), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n546), .A2(KEYINPUT30), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n537), .B2(new_n540), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(KEYINPUT30), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n492), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT70), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n553), .B(new_n455), .C1(new_n513), .C2(new_n527), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n535), .B2(new_n455), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n455), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G227gat), .A2(G233gat), .ZN(new_n559));
  AOI211_X1 g358(.A(KEYINPUT72), .B(KEYINPUT34), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT34), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n513), .A2(new_n527), .A3(new_n455), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n557), .B1(KEYINPUT70), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n559), .A3(new_n554), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT72), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G15gat), .B(G43gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT71), .ZN(new_n569));
  XOR2_X1   g368(.A(G71gat), .B(G99gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n559), .B1(new_n563), .B2(new_n554), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(KEYINPUT33), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT32), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT32), .B1(new_n558), .B2(new_n559), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT33), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n578), .B1(new_n558), .B2(new_n559), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n577), .B1(new_n579), .B2(new_n571), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n567), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n573), .A2(new_n575), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n577), .A3(new_n571), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n582), .B(new_n583), .C1(new_n566), .C2(new_n560), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n435), .ZN(new_n586));
  INV_X1    g385(.A(new_n404), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n379), .B2(new_n393), .ZN(new_n588));
  AOI211_X1 g387(.A(G22gat), .B(new_n588), .C1(new_n430), .C2(new_n431), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n433), .B1(new_n432), .B2(new_n405), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n424), .A2(new_n434), .A3(new_n435), .ZN(new_n592));
  INV_X1    g391(.A(new_n351), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n438), .A2(new_n552), .A3(new_n585), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT35), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT35), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n550), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT6), .B1(new_n480), .B2(new_n486), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT88), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n470), .A2(new_n475), .ZN(new_n601));
  INV_X1    g400(.A(new_n462), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n479), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT87), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT87), .B1(new_n476), .B2(new_n479), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n600), .B1(new_n608), .B2(new_n485), .ZN(new_n609));
  AOI211_X1 g408(.A(KEYINPUT88), .B(new_n486), .C1(new_n606), .C2(new_n607), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n599), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n598), .B1(new_n611), .B2(new_n491), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n612), .A2(new_n585), .A3(new_n594), .A4(new_n438), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n581), .A2(new_n584), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT36), .B1(new_n615), .B2(KEYINPUT73), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT73), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n618));
  AOI211_X1 g417(.A(new_n617), .B(new_n618), .C1(new_n581), .C2(new_n584), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT38), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT37), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n537), .A2(new_n540), .A3(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n623), .A2(new_n544), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n537), .A2(new_n540), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT37), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n621), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n529), .A2(new_n531), .A3(new_n536), .A4(new_n400), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n399), .B1(new_n538), .B2(new_n539), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n629), .A3(KEYINPUT37), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n630), .A2(new_n623), .A3(new_n621), .A4(new_n544), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n546), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n611), .A2(new_n491), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n550), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n460), .B1(new_n477), .B2(new_n478), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n636), .B(KEYINPUT39), .C1(new_n460), .C2(new_n458), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n637), .B(new_n486), .C1(KEYINPUT39), .C2(new_n636), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT40), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n635), .B(new_n639), .C1(new_n609), .C2(new_n610), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n634), .A2(new_n640), .A3(new_n594), .A4(new_n438), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n438), .A2(new_n594), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n551), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n620), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n350), .B1(new_n614), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n325), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n492), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(new_n278), .ZN(G1324gat));
  NAND2_X1  g447(.A1(new_n274), .A2(KEYINPUT42), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n646), .A2(new_n550), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n650), .A2(KEYINPUT104), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(KEYINPUT104), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT16), .B(G8gat), .Z(new_n654));
  NAND3_X1  g453(.A1(new_n650), .A2(KEYINPUT42), .A3(new_n654), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n653), .B(new_n655), .C1(KEYINPUT42), .C2(new_n654), .ZN(G1325gat));
  INV_X1    g455(.A(new_n646), .ZN(new_n657));
  AOI21_X1  g456(.A(G15gat), .B1(new_n657), .B2(new_n585), .ZN(new_n658));
  INV_X1    g457(.A(new_n620), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(G15gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT105), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n658), .B1(new_n657), .B2(new_n661), .ZN(G1326gat));
  INV_X1    g461(.A(new_n642), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n646), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT43), .B(G22gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  NAND2_X1  g465(.A1(new_n241), .A2(new_n244), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n596), .A2(new_n668), .A3(new_n613), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n644), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n596), .B2(new_n613), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n667), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n614), .A2(new_n644), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(KEYINPUT44), .A3(new_n667), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n294), .A2(new_n350), .A3(new_n324), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n492), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(G29gat), .ZN(new_n682));
  INV_X1    g481(.A(new_n294), .ZN(new_n683));
  INV_X1    g482(.A(new_n324), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n667), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT106), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n645), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n687), .A2(G29gat), .A3(new_n492), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n682), .A2(new_n690), .ZN(G1328gat));
  INV_X1    g490(.A(G36gat), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n692), .B1(new_n679), .B2(new_n635), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n686), .A2(new_n645), .A3(new_n692), .A4(new_n635), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT46), .ZN(new_n695));
  OR3_X1    g494(.A1(new_n693), .A2(KEYINPUT109), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT109), .B1(new_n693), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(G1329gat));
  INV_X1    g497(.A(G43gat), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n677), .A2(new_n659), .A3(new_n678), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n700), .A2(KEYINPUT110), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(KEYINPUT110), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n687), .A2(G43gat), .A3(new_n615), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT47), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n700), .B2(G43gat), .ZN(new_n707));
  OAI22_X1  g506(.A1(new_n703), .A2(new_n706), .B1(KEYINPUT47), .B2(new_n707), .ZN(G1330gat));
  NAND3_X1  g507(.A1(new_n679), .A2(G50gat), .A3(new_n642), .ZN(new_n709));
  INV_X1    g508(.A(G50gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(new_n687), .B2(new_n663), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g512(.A1(new_n614), .A2(KEYINPUT108), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(new_n644), .A3(new_n669), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n295), .A2(new_n349), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n324), .A3(new_n716), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n717), .A2(new_n492), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g518(.A(new_n717), .B(KEYINPUT111), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n720), .A2(new_n635), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n721), .A2(KEYINPUT49), .A3(G64gat), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT49), .B(G64gat), .Z(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n721), .B2(new_n723), .ZN(G1333gat));
  NAND3_X1  g523(.A1(new_n720), .A2(G71gat), .A3(new_n659), .ZN(new_n725));
  INV_X1    g524(.A(G71gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n717), .B2(new_n615), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g528(.A1(new_n720), .A2(new_n642), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g530(.A1(new_n294), .A2(new_n349), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n324), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT112), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n677), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735), .B2(new_n492), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n715), .A2(new_n667), .A3(new_n732), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n715), .A2(KEYINPUT51), .A3(new_n667), .A4(new_n732), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n741), .A2(new_n217), .A3(new_n680), .A4(new_n324), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n736), .A2(new_n742), .ZN(G1336gat));
  NOR3_X1   g542(.A1(new_n684), .A2(G92gat), .A3(new_n550), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n674), .A2(new_n635), .A3(new_n676), .A4(new_n734), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G92gat), .ZN(new_n747));
  XOR2_X1   g546(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n748));
  NAND3_X1  g547(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n739), .A2(KEYINPUT114), .A3(new_n740), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n737), .A2(new_n751), .A3(new_n738), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n744), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n746), .A2(KEYINPUT113), .A3(G92gat), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT113), .B1(new_n746), .B2(G92gat), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n756), .A2(KEYINPUT115), .A3(KEYINPUT52), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT115), .B1(new_n756), .B2(KEYINPUT52), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n749), .B1(new_n757), .B2(new_n758), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n735), .B2(new_n620), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n615), .A2(G99gat), .A3(new_n684), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n741), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(G1338gat));
  OAI21_X1  g562(.A(G106gat), .B1(new_n735), .B2(new_n663), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n663), .A2(G106gat), .A3(new_n684), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n752), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT53), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT53), .B1(new_n741), .B2(new_n765), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n764), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(G1339gat));
  OAI22_X1  g570(.A1(new_n330), .A2(new_n331), .B1(new_n336), .B2(new_n337), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n344), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n348), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n241), .B2(new_n244), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT118), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n231), .A2(KEYINPUT10), .A3(new_n287), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT101), .B1(new_n313), .B2(new_n306), .ZN(new_n778));
  AOI211_X1 g577(.A(new_n308), .B(KEYINPUT10), .C1(new_n311), .C2(new_n312), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n777), .B(new_n316), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n780), .B(KEYINPUT54), .C1(new_n315), .C2(new_n303), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  INV_X1    g582(.A(new_n316), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n781), .A2(new_n320), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(KEYINPUT117), .A3(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n781), .A2(KEYINPUT55), .A3(new_n320), .A4(new_n785), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n323), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT117), .B1(new_n786), .B2(new_n787), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n776), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n791), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n789), .A2(new_n323), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n793), .A2(new_n794), .A3(KEYINPUT118), .A4(new_n788), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n775), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n792), .A2(new_n349), .A3(new_n795), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n348), .A2(new_n773), .A3(new_n324), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(KEYINPUT119), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n245), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT119), .B1(new_n797), .B2(new_n798), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n796), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n683), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n716), .A2(new_n684), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n642), .A2(new_n615), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n680), .A3(new_n806), .ZN(new_n807));
  OR3_X1    g606(.A1(new_n807), .A2(KEYINPUT120), .A3(new_n635), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT120), .B1(new_n807), .B2(new_n635), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n350), .A2(new_n447), .ZN(new_n811));
  INV_X1    g610(.A(new_n807), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n550), .A3(new_n349), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n810), .A2(new_n811), .B1(new_n447), .B2(new_n813), .ZN(G1340gat));
  NOR2_X1   g613(.A1(new_n684), .A2(new_n445), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(new_n550), .A3(new_n324), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n810), .A2(new_n815), .B1(new_n445), .B2(new_n816), .ZN(G1341gat));
  AOI21_X1  g616(.A(new_n683), .B1(new_n808), .B2(new_n809), .ZN(new_n818));
  INV_X1    g617(.A(G127gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n812), .A2(new_n550), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n294), .A2(new_n819), .ZN(new_n821));
  OAI22_X1  g620(.A1(new_n818), .A2(new_n819), .B1(new_n820), .B2(new_n821), .ZN(G1342gat));
  NOR2_X1   g621(.A1(new_n245), .A2(new_n635), .ZN(new_n823));
  INV_X1    g622(.A(G134gat), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT56), .B1(new_n807), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT121), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n807), .A2(new_n825), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n245), .B1(new_n808), .B2(new_n809), .ZN(new_n829));
  OAI221_X1 g628(.A(new_n827), .B1(KEYINPUT56), .B2(new_n828), .C1(new_n824), .C2(new_n829), .ZN(G1343gat));
  NAND2_X1  g629(.A1(new_n786), .A2(new_n787), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n349), .A2(new_n831), .A3(new_n794), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n798), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n245), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n294), .B1(new_n796), .B2(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n295), .A2(new_n349), .A3(new_n324), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n642), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT57), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n659), .A2(new_n492), .A3(new_n635), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n797), .A2(new_n798), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n245), .A3(new_n799), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n294), .B1(new_n843), .B2(new_n796), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n642), .B1(new_n844), .B2(new_n836), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n838), .B(new_n839), .C1(KEYINPUT57), .C2(new_n845), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n846), .A2(new_n383), .A3(new_n350), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n659), .A2(new_n663), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(KEYINPUT122), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n805), .A2(new_n680), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n635), .ZN(new_n851));
  AOI21_X1  g650(.A(G141gat), .B1(new_n851), .B2(new_n349), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853));
  OR3_X1    g652(.A1(new_n847), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n847), .B2(new_n852), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1344gat));
  INV_X1    g655(.A(KEYINPUT59), .ZN(new_n857));
  AOI211_X1 g656(.A(new_n857), .B(G148gat), .C1(new_n851), .C2(new_n324), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n846), .B2(new_n684), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n642), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n790), .A2(new_n791), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n775), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n834), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n683), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n861), .B1(new_n804), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n845), .B2(KEYINPUT57), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n867), .A2(KEYINPUT59), .A3(new_n324), .A4(new_n839), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n859), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n858), .B1(new_n869), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g669(.A(G155gat), .B1(new_n846), .B2(new_n683), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n851), .A2(new_n380), .A3(new_n294), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1346gat));
  OAI21_X1  g672(.A(G162gat), .B1(new_n846), .B2(new_n245), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n823), .A2(new_n381), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n850), .B2(new_n875), .ZN(G1347gat));
  NOR2_X1   g675(.A1(new_n680), .A2(new_n550), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n878), .B1(new_n803), .B2(new_n804), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n806), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n350), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n523), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n882), .B1(new_n342), .B2(new_n881), .ZN(G1348gat));
  NOR2_X1   g682(.A1(new_n880), .A2(new_n684), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(new_n508), .ZN(G1349gat));
  NOR2_X1   g684(.A1(new_n880), .A2(new_n683), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n517), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n502), .B2(new_n886), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g688(.A1(new_n879), .A2(new_n806), .A3(new_n667), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n891), .A3(G190gat), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n891), .B1(new_n890), .B2(G190gat), .ZN(new_n894));
  INV_X1    g693(.A(new_n501), .ZN(new_n895));
  OAI22_X1  g694(.A1(new_n893), .A2(new_n894), .B1(new_n895), .B2(new_n890), .ZN(G1351gat));
  AOI21_X1  g695(.A(new_n294), .B1(new_n863), .B2(new_n834), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n860), .B(new_n642), .C1(new_n836), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n659), .A2(new_n878), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n663), .B1(new_n803), .B2(new_n804), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n898), .B(new_n899), .C1(new_n900), .C2(new_n860), .ZN(new_n901));
  INV_X1    g700(.A(G197gat), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n901), .A2(new_n902), .A3(new_n350), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n848), .B(new_n877), .C1(new_n844), .C2(new_n836), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(G197gat), .B1(new_n905), .B2(new_n349), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n903), .A2(new_n906), .ZN(G1352gat));
  NAND3_X1  g706(.A1(new_n867), .A2(new_n324), .A3(new_n899), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(G204gat), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n684), .A2(G204gat), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n910), .B1(new_n904), .B2(new_n912), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n879), .A2(KEYINPUT123), .A3(new_n848), .A4(new_n911), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT62), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT62), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n909), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT124), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n909), .B(new_n919), .C1(new_n915), .C2(new_n916), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1353gat));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n922));
  OAI21_X1  g721(.A(G211gat), .B1(new_n901), .B2(new_n683), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT63), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n867), .A2(new_n294), .A3(new_n899), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n926), .A2(KEYINPUT125), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n923), .A2(new_n924), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n905), .A2(new_n356), .A3(new_n294), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1354gat));
  AOI21_X1  g730(.A(G218gat), .B1(new_n905), .B2(new_n667), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n901), .A2(KEYINPUT126), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n867), .A2(new_n935), .A3(new_n899), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n245), .A2(new_n365), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  OAI211_X1 g738(.A(KEYINPUT127), .B(new_n933), .C1(new_n937), .C2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n934), .B2(new_n936), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n932), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n940), .A2(new_n943), .ZN(G1355gat));
endmodule


