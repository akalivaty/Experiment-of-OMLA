//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n450, new_n451, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n633, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g024(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n450));
  AND2_X1   g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(G223));
  NAND2_X1  g027(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g028(.A1(new_n451), .A2(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n456), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT66), .Z(new_n462));
  AND2_X1   g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XOR2_X1   g038(.A(new_n463), .B(KEYINPUT67), .Z(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n469), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n472), .A2(new_n465), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n468), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n470), .A2(new_n475), .ZN(new_n480));
  INV_X1    g055(.A(G125), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n478), .B1(new_n485), .B2(new_n486), .ZN(G160));
  OAI21_X1  g062(.A(KEYINPUT70), .B1(G100), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NOR3_X1   g064(.A1(KEYINPUT70), .A2(G100), .A3(G2105), .ZN(new_n490));
  OAI221_X1 g065(.A(G2104), .B1(G112), .B2(new_n465), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G124), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n472), .A2(G2105), .A3(new_n473), .A4(new_n475), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n476), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(G136), .B2(new_n495), .ZN(G162));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n465), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  OAI22_X1  g074(.A1(new_n493), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n470), .A2(new_n475), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(new_n465), .A3(G138), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT71), .B1(new_n480), .B2(new_n504), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G138), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT4), .B1(new_n476), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n500), .B1(new_n508), .B2(new_n510), .ZN(G164));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g089(.A(G543), .B1(KEYINPUT74), .B2(KEYINPUT5), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(KEYINPUT74), .B2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT72), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(KEYINPUT73), .B1(new_n522), .B2(KEYINPUT5), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT5), .ZN(new_n525));
  AOI211_X1 g100(.A(new_n524), .B(new_n525), .C1(new_n519), .C2(new_n521), .ZN(new_n526));
  OAI211_X1 g101(.A(G62), .B(new_n517), .C1(new_n523), .C2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n514), .B1(new_n527), .B2(KEYINPUT75), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT72), .B(G543), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n524), .B1(new_n529), .B2(new_n525), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n520), .A2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n518), .A2(KEYINPUT72), .ZN(new_n532));
  OAI211_X1 g107(.A(KEYINPUT73), .B(KEYINPUT5), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n516), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n534), .A2(new_n535), .A3(G62), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n512), .B1(new_n528), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT6), .B(G651), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n538), .A2(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G50), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n534), .A2(new_n538), .ZN(new_n541));
  INV_X1    g116(.A(G88), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n537), .A2(new_n543), .ZN(G166));
  AND2_X1   g119(.A1(new_n534), .A2(new_n538), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G89), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n534), .A2(G63), .A3(G651), .ZN(new_n547));
  NAND3_X1  g122(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(KEYINPUT7), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n548), .A2(KEYINPUT7), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n539), .A2(G51), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n546), .A2(new_n547), .A3(new_n551), .ZN(G286));
  INV_X1    g127(.A(G286), .ZN(G168));
  AOI22_X1  g128(.A1(new_n534), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n512), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n539), .A2(G52), .ZN(new_n556));
  INV_X1    g131(.A(G90), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n541), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(G171));
  AOI22_X1  g134(.A1(new_n534), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n512), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n539), .A2(G43), .ZN(new_n562));
  INV_X1    g137(.A(G81), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n541), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  AOI22_X1  g145(.A1(new_n534), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(new_n512), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n538), .A2(G53), .A3(G543), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(G91), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n541), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  INV_X1    g154(.A(G166), .ZN(G303));
  OAI21_X1  g155(.A(G651), .B1(new_n534), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n538), .A2(G49), .A3(G543), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT76), .Z(new_n583));
  NAND3_X1  g158(.A1(new_n534), .A2(G87), .A3(new_n538), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(G288));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  AOI211_X1 g161(.A(new_n586), .B(new_n516), .C1(new_n530), .C2(new_n533), .ZN(new_n587));
  INV_X1    g162(.A(G73), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n518), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n538), .A2(G48), .A3(G543), .ZN(new_n591));
  XOR2_X1   g166(.A(new_n591), .B(KEYINPUT78), .Z(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n530), .A2(new_n533), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n594), .A2(G86), .A3(new_n517), .A4(new_n538), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT77), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n534), .A2(new_n597), .A3(G86), .A4(new_n538), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n590), .A2(new_n593), .A3(new_n596), .A4(new_n598), .ZN(G305));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n601));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n534), .B2(G60), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n601), .B1(new_n604), .B2(new_n512), .ZN(new_n605));
  INV_X1    g180(.A(G60), .ZN(new_n606));
  AOI211_X1 g181(.A(new_n606), .B(new_n516), .C1(new_n530), .C2(new_n533), .ZN(new_n607));
  OAI211_X1 g182(.A(KEYINPUT79), .B(G651), .C1(new_n607), .C2(new_n603), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n534), .A2(G85), .A3(new_n538), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n539), .A2(G47), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n600), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  AOI211_X1 g189(.A(KEYINPUT80), .B(new_n612), .C1(new_n605), .C2(new_n608), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(G290));
  NAND2_X1  g192(.A1(G301), .A2(G868), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n534), .A2(G92), .A3(new_n538), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT10), .Z(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n594), .A2(new_n517), .ZN(new_n622));
  INV_X1    g197(.A(G66), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n624), .A2(G651), .B1(G54), .B2(new_n539), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n618), .B1(new_n627), .B2(G868), .ZN(G284));
  OAI21_X1  g203(.A(new_n618), .B1(new_n627), .B2(G868), .ZN(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n577), .B2(G868), .ZN(G297));
  OAI21_X1  g206(.A(new_n630), .B1(new_n577), .B2(G868), .ZN(G280));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n627), .B1(new_n633), .B2(G860), .ZN(G148));
  NAND3_X1  g209(.A1(new_n620), .A2(new_n625), .A3(new_n633), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G868), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n495), .A2(G135), .ZN(new_n639));
  INV_X1    g214(.A(G123), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n465), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  OAI221_X1 g217(.A(new_n639), .B1(new_n640), .B2(new_n493), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n643), .A2(KEYINPUT81), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(KEYINPUT81), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  NOR2_X1   g222(.A1(new_n480), .A2(new_n466), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT13), .B(G2100), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n651), .ZN(G156));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n658), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(G401));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT82), .ZN(new_n670));
  NOR2_X1   g245(.A1(G2072), .A2(G2078), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n444), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n668), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(KEYINPUT17), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n673), .B1(new_n670), .B2(new_n674), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n668), .B(new_n669), .C1(new_n444), .C2(new_n671), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT18), .Z(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n670), .A3(new_n668), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2096), .B(G2100), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1971), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(new_n686), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  AOI211_X1 g266(.A(new_n688), .B(new_n691), .C1(new_n683), .C2(new_n687), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT84), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT85), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(G229));
  INV_X1    g275(.A(KEYINPUT24), .ZN(new_n701));
  INV_X1    g276(.A(G34), .ZN(new_n702));
  AOI21_X1  g277(.A(G29), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n701), .B2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(G160), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(G2084), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT94), .Z(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G5), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G171), .B2(new_n709), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n708), .B1(G1961), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(G162), .A2(G29), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G29), .B2(G35), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G2090), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n712), .B(new_n718), .C1(G1961), .C2(new_n711), .ZN(new_n719));
  NAND2_X1  g294(.A1(G168), .A2(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G16), .B2(G21), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT93), .B(G1966), .Z(new_n722));
  NOR2_X1   g297(.A1(G27), .A2(G29), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G164), .B2(G29), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n721), .A2(new_n722), .B1(G2078), .B2(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(G2078), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n725), .B(new_n726), .C1(new_n722), .C2(new_n721), .ZN(new_n727));
  INV_X1    g302(.A(new_n646), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n728), .A2(G29), .B1(G2084), .B2(new_n706), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n705), .A2(G32), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT26), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n733), .A2(new_n734), .B1(G105), .B2(new_n467), .ZN(new_n735));
  INV_X1    g310(.A(G129), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n493), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G141), .B2(new_n495), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n730), .B1(new_n738), .B2(new_n705), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT27), .B(G1996), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT92), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n739), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n705), .A2(G26), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT28), .ZN(new_n744));
  OR2_X1    g319(.A1(G104), .A2(G2105), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n745), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n746));
  INV_X1    g321(.A(G128), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n493), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G140), .B2(new_n495), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n744), .B1(new_n749), .B2(new_n705), .ZN(new_n750));
  INV_X1    g325(.A(G2067), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n705), .A2(G33), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n495), .A2(G139), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n755));
  NAND3_X1  g330(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n501), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n754), .B(new_n757), .C1(new_n465), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n753), .B1(new_n759), .B2(G29), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(new_n442), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n442), .ZN(new_n762));
  INV_X1    g337(.A(G28), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(KEYINPUT30), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n763), .B2(KEYINPUT30), .ZN(new_n765));
  OR2_X1    g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  NAND2_X1  g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n764), .A2(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AND3_X1   g343(.A1(new_n761), .A2(new_n762), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n729), .A2(new_n742), .A3(new_n752), .A4(new_n769), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n719), .A2(new_n727), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n627), .A2(new_n709), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G4), .B2(new_n709), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT89), .B(G1348), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G16), .A2(G19), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n565), .B2(G16), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT90), .B(G1341), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n773), .A2(new_n774), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n771), .A2(new_n775), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n709), .A2(G20), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT23), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n577), .B2(new_n709), .ZN(new_n784));
  INV_X1    g359(.A(G1956), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n717), .B2(new_n716), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT96), .Z(new_n788));
  NOR2_X1   g363(.A1(new_n781), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n709), .A2(G22), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G166), .B2(new_n709), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1971), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(KEYINPUT87), .ZN(new_n794));
  INV_X1    g369(.A(G1971), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n792), .B(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT87), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n709), .A2(G23), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G288), .B2(G16), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT33), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1976), .ZN(new_n806));
  MUX2_X1   g381(.A(G6), .B(G305), .S(G16), .Z(new_n807));
  XOR2_X1   g382(.A(KEYINPUT32), .B(G1981), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n794), .A2(new_n798), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT88), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT34), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n810), .A2(new_n811), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n810), .A2(new_n811), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n815), .A2(KEYINPUT34), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n616), .A2(G16), .ZN(new_n818));
  NOR2_X1   g393(.A1(G16), .A2(G24), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n818), .A2(G1986), .A3(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(G25), .A2(G29), .ZN(new_n823));
  INV_X1    g398(.A(G119), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n465), .A2(G107), .ZN(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n826));
  OAI22_X1  g401(.A1(new_n493), .A2(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G131), .B2(new_n495), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n823), .B1(new_n828), .B2(G29), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT86), .Z(new_n830));
  XOR2_X1   g405(.A(KEYINPUT35), .B(G1991), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(G1986), .B1(new_n818), .B2(new_n820), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n822), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n814), .A2(new_n817), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT36), .ZN(new_n836));
  INV_X1    g411(.A(new_n834), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n812), .B2(new_n813), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT36), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n838), .A2(new_n839), .A3(new_n817), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n790), .B1(new_n836), .B2(new_n840), .ZN(G311));
  AND3_X1   g416(.A1(new_n838), .A2(new_n839), .A3(new_n817), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n839), .B1(new_n838), .B2(new_n817), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n789), .B1(new_n842), .B2(new_n843), .ZN(G150));
  NOR2_X1   g419(.A1(new_n626), .A2(new_n633), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n539), .A2(G55), .ZN(new_n848));
  INV_X1    g423(.A(G93), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n541), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n534), .A2(G67), .ZN(new_n851));
  NAND2_X1  g426(.A1(G80), .A2(G543), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n512), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n565), .A2(new_n854), .ZN(new_n855));
  OAI22_X1  g430(.A1(new_n561), .A2(new_n564), .B1(new_n850), .B2(new_n853), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n847), .B(new_n857), .Z(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n859));
  INV_X1    g434(.A(G860), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n854), .A2(new_n860), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(new_n646), .B(KEYINPUT98), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G162), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G160), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n510), .A2(new_n507), .A3(new_n506), .ZN(new_n869));
  INV_X1    g444(.A(new_n500), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n749), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n759), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n738), .ZN(new_n874));
  INV_X1    g449(.A(G130), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n465), .A2(G118), .ZN(new_n876));
  OAI21_X1  g451(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n877));
  OAI22_X1  g452(.A1(new_n493), .A2(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(G142), .B2(new_n495), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(new_n649), .Z(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n828), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n874), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n868), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n874), .A2(new_n881), .ZN(new_n884));
  AOI21_X1  g459(.A(G37), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT99), .B1(new_n874), .B2(new_n881), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n882), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n868), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n885), .A2(KEYINPUT40), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT40), .B1(new_n885), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(G395));
  NAND2_X1  g466(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n892));
  OR2_X1    g467(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n893));
  INV_X1    g468(.A(G288), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n614), .B2(new_n615), .ZN(new_n895));
  OAI22_X1  g470(.A1(new_n622), .A2(new_n586), .B1(new_n588), .B2(new_n518), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n592), .B1(new_n896), .B2(G651), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n596), .A2(new_n598), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n897), .B(new_n898), .C1(new_n537), .C2(new_n543), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n527), .A2(KEYINPUT75), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n536), .A3(new_n513), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(G651), .ZN(new_n902));
  INV_X1    g477(.A(new_n543), .ZN(new_n903));
  NAND3_X1  g478(.A1(G305), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g480(.A(G60), .B(new_n517), .C1(new_n523), .C2(new_n526), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n602), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT79), .B1(new_n907), .B2(G651), .ZN(new_n908));
  AOI211_X1 g483(.A(new_n601), .B(new_n512), .C1(new_n906), .C2(new_n602), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n613), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT80), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n609), .A2(new_n600), .A3(new_n613), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(G288), .A3(new_n912), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n895), .A2(new_n905), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n905), .B1(new_n895), .B2(new_n913), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n892), .B(new_n893), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n905), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n614), .A2(new_n615), .A3(new_n894), .ZN(new_n918));
  AOI21_X1  g493(.A(G288), .B1(new_n911), .B2(new_n912), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n895), .A2(new_n913), .A3(new_n905), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n920), .A2(KEYINPUT100), .A3(KEYINPUT42), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n916), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n627), .A2(new_n577), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n577), .B1(new_n620), .B2(new_n625), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(KEYINPUT41), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n626), .A2(G299), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n928), .B1(new_n929), .B2(new_n925), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n635), .B1(new_n856), .B2(new_n855), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n857), .B1(new_n633), .B2(new_n627), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n927), .B(new_n930), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n931), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n929), .A2(new_n925), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n923), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT102), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n937), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT101), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n941), .A2(new_n916), .A3(new_n942), .A4(new_n922), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT101), .B1(new_n923), .B2(new_n937), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n923), .A2(KEYINPUT102), .A3(new_n937), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n940), .A2(new_n943), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(G868), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n854), .A2(G868), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(G295));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n947), .B2(new_n949), .ZN(new_n952));
  AOI211_X1 g527(.A(KEYINPUT103), .B(new_n948), .C1(new_n946), .C2(G868), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(G331));
  NAND3_X1  g529(.A1(new_n855), .A2(G301), .A3(new_n856), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(G301), .B1(new_n855), .B2(new_n856), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n956), .A2(G286), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n857), .A2(G171), .ZN(new_n959));
  AOI21_X1  g534(.A(G168), .B1(new_n959), .B2(new_n955), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n935), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(G286), .B1(new_n956), .B2(new_n957), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(G168), .A3(new_n955), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n962), .A2(new_n927), .A3(new_n963), .A4(new_n930), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n920), .A2(new_n921), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n961), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(G37), .B1(new_n966), .B2(KEYINPUT104), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n961), .A2(new_n964), .ZN(new_n968));
  INV_X1    g543(.A(new_n965), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n961), .A2(new_n964), .A3(new_n965), .A4(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n967), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n961), .A2(new_n964), .A3(KEYINPUT105), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n975), .B(new_n969), .C1(KEYINPUT105), .C2(new_n961), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n976), .A2(new_n967), .A3(new_n977), .A4(new_n972), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n973), .A2(new_n977), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n976), .A2(new_n967), .A3(KEYINPUT43), .A4(new_n972), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  MUX2_X1   g557(.A(new_n979), .B(new_n982), .S(KEYINPUT44), .Z(G397));
  INV_X1    g558(.A(G1986), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n616), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n616), .A2(new_n984), .ZN(new_n987));
  OR3_X1    g562(.A1(new_n986), .A2(KEYINPUT106), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(G160), .A2(G40), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(G164), .B2(G1384), .ZN(new_n991));
  AOI211_X1 g566(.A(new_n989), .B(new_n991), .C1(new_n987), .C2(KEYINPUT106), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n989), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n738), .B(G1996), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n749), .B(G2067), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n828), .A2(new_n831), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n828), .A2(new_n831), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n988), .A2(new_n992), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT107), .Z(new_n1000));
  INV_X1    g575(.A(KEYINPUT125), .ZN(new_n1001));
  XOR2_X1   g576(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1002), .B1(G166), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n1005));
  OAI221_X1 g580(.A(G8), .B1(new_n1005), .B2(KEYINPUT55), .C1(new_n537), .C2(new_n543), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1384), .B1(new_n869), .B2(new_n870), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1012));
  INV_X1    g587(.A(G40), .ZN(new_n1013));
  AOI211_X1 g588(.A(new_n1013), .B(new_n478), .C1(new_n485), .C2(new_n486), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT110), .B(G2090), .Z(new_n1015));
  NAND4_X1  g590(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n990), .A2(G1384), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT109), .B1(new_n871), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1018), .ZN(new_n1021));
  NOR3_X1   g596(.A1(G164), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n1009), .B2(KEYINPUT45), .ZN(new_n1025));
  OAI211_X1 g600(.A(KEYINPUT108), .B(new_n990), .C1(G164), .C2(G1384), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1023), .A2(new_n1014), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1017), .B1(new_n1027), .B2(new_n795), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT113), .B(G8), .Z(new_n1029));
  OAI21_X1  g604(.A(new_n1008), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n871), .A2(KEYINPUT109), .A3(new_n1018), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1020), .B1(G164), .B2(new_n1021), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n1033), .A3(new_n1014), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n795), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1384), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n871), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n989), .B1(new_n1037), .B2(KEYINPUT50), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n1011), .A4(new_n1015), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1016), .A2(KEYINPUT111), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1035), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(G8), .A3(new_n1007), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n894), .A2(G1976), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1029), .B1(new_n1014), .B2(new_n1009), .ZN(new_n1045));
  INV_X1    g620(.A(G1976), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(G288), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1048), .B(KEYINPUT114), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1045), .ZN(new_n1050));
  INV_X1    g625(.A(G1981), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n897), .A2(new_n898), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n590), .A2(new_n593), .ZN(new_n1053));
  INV_X1    g628(.A(new_n595), .ZN(new_n1054));
  OAI21_X1  g629(.A(G1981), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT49), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1050), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1052), .A2(new_n1055), .A3(KEYINPUT49), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1058), .A2(new_n1059), .B1(KEYINPUT52), .B2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1030), .A2(new_n1043), .A3(new_n1049), .A4(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1032), .A2(new_n1033), .A3(new_n1014), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1065), .A2(new_n443), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1067));
  INV_X1    g642(.A(G1961), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1038), .A2(new_n1011), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1066), .A2(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n871), .A2(new_n1071), .A3(new_n1018), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(G164), .B2(new_n1021), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n991), .A2(new_n1014), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1076));
  OR3_X1    g651(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(G301), .B1(new_n1070), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1069), .A2(new_n1068), .ZN(new_n1079));
  INV_X1    g654(.A(new_n483), .ZN(new_n1080));
  NOR4_X1   g655(.A1(new_n1080), .A2(new_n478), .A3(new_n1013), .A4(new_n1076), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1023), .A2(new_n991), .A3(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1031), .A2(new_n1034), .A3(G2078), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1067), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1079), .B(new_n1082), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(G171), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1064), .B1(new_n1078), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(G171), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1077), .B(new_n1079), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1088), .B(KEYINPUT54), .C1(G171), .C2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1063), .A2(new_n1087), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n722), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n1093));
  INV_X1    g668(.A(G2084), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1011), .A2(new_n1012), .A3(new_n1094), .A4(new_n1014), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1092), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1093), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1096), .A2(new_n1097), .A3(new_n1003), .ZN(new_n1098));
  NOR2_X1   g673(.A1(G168), .A2(new_n1029), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT51), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1029), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1099), .A2(KEYINPUT51), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1029), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1099), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT123), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1101), .A2(KEYINPUT121), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1092), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1099), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT122), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n1099), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1100), .A2(new_n1112), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1001), .B1(new_n1091), .B2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1065), .A2(new_n1025), .A3(new_n1026), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1069), .A2(new_n785), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n577), .B(KEYINPUT57), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(KEYINPUT118), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1011), .A2(new_n1014), .A3(new_n1012), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1014), .A2(new_n1009), .ZN(new_n1129));
  OAI22_X1  g704(.A1(new_n1128), .A2(G1348), .B1(G2067), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n627), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1125), .B(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1127), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(KEYINPUT61), .B(new_n1126), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1130), .A2(KEYINPUT60), .A3(new_n626), .ZN(new_n1138));
  INV_X1    g713(.A(G1348), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1129), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1069), .A2(new_n1139), .B1(new_n751), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n626), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1131), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1138), .B1(new_n1143), .B2(KEYINPUT60), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1027), .A2(G1996), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(G1341), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1140), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n565), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1149), .A2(KEYINPUT59), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(KEYINPUT59), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1137), .B(new_n1144), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n1134), .A2(new_n1125), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT61), .B1(new_n1127), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1136), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1089), .A2(G171), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1156), .A2(new_n1064), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1062), .B1(new_n1088), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1113), .A2(G8), .A3(new_n1114), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1109), .B1(new_n1159), .B2(new_n1108), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1118), .B1(new_n1117), .B2(new_n1099), .ZN(new_n1162));
  NOR4_X1   g737(.A1(new_n1096), .A2(new_n1097), .A3(KEYINPUT122), .A4(new_n1108), .ZN(new_n1163));
  OAI22_X1  g738(.A1(new_n1160), .A2(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1158), .A2(new_n1164), .A3(KEYINPUT125), .A4(new_n1087), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1121), .A2(new_n1155), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(KEYINPUT62), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1119), .A2(new_n1116), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1168), .B(new_n1169), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1063), .A2(new_n1078), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1167), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1107), .A2(G168), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1173), .B1(new_n1062), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(KEYINPUT117), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT117), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1177), .B(new_n1173), .C1(new_n1062), .C2(new_n1174), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1042), .A2(G8), .A3(new_n1007), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1179), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1042), .A2(G8), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1008), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1060), .A2(KEYINPUT52), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1183), .A2(new_n1049), .A3(new_n1184), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1185), .A2(KEYINPUT115), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1185), .A2(KEYINPUT115), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1180), .B(new_n1182), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1176), .A2(new_n1178), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1183), .A2(new_n1046), .A3(new_n894), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1050), .B1(new_n1190), .B2(new_n1052), .ZN(new_n1191));
  OR2_X1    g766(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1191), .B1(new_n1192), .B2(new_n1179), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1172), .A2(new_n1189), .A3(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1000), .B1(new_n1166), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n749), .A2(new_n751), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n994), .A2(new_n995), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1196), .B1(new_n1197), .B2(new_n996), .ZN(new_n1198));
  AND2_X1   g773(.A1(new_n1198), .A2(new_n993), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n995), .A2(new_n738), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n993), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n1201), .B(KEYINPUT126), .Z(new_n1202));
  NOR3_X1   g777(.A1(new_n991), .A2(new_n989), .A3(G1996), .ZN(new_n1203));
  XOR2_X1   g778(.A(new_n1203), .B(KEYINPUT46), .Z(new_n1204));
  NAND2_X1  g779(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g780(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n1205), .B(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n998), .A2(new_n993), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n986), .A2(new_n993), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT48), .ZN(new_n1210));
  AOI211_X1 g785(.A(new_n1199), .B(new_n1207), .C1(new_n1208), .C2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1195), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g787(.A1(new_n885), .A2(new_n888), .ZN(new_n1214));
  INV_X1    g788(.A(new_n463), .ZN(new_n1215));
  NOR4_X1   g789(.A1(G229), .A2(new_n1215), .A3(G401), .A4(G227), .ZN(new_n1216));
  NAND3_X1  g790(.A1(new_n1214), .A2(new_n1216), .A3(new_n979), .ZN(G225));
  INV_X1    g791(.A(G225), .ZN(G308));
endmodule


