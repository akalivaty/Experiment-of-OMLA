//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n526, new_n527,
    new_n528, new_n529, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n540, new_n541, new_n542, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n552, new_n553, new_n554,
    new_n555, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n590, new_n591, new_n594, new_n596, new_n597, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT65), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n466), .A2(new_n472), .A3(G125), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n466), .A2(new_n472), .A3(KEYINPUT66), .A4(G125), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n461), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  INV_X1    g054(.A(G101), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n461), .A2(G2104), .ZN(new_n481));
  OAI22_X1  g056(.A1(new_n478), .A2(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n477), .A2(new_n482), .ZN(G160));
  AOI21_X1  g058(.A(new_n461), .B1(new_n469), .B2(new_n471), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n485), .B(new_n487), .C1(new_n488), .C2(new_n478), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n491), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n466), .A2(new_n472), .A3(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n461), .C1(new_n464), .C2(new_n465), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n498));
  OAI211_X1 g073(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n505));
  XNOR2_X1  g080(.A(new_n505), .B(KEYINPUT67), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n506), .A2(G543), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n506), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G88), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n513), .A2(new_n504), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n509), .A2(new_n512), .A3(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT68), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n518), .A2(KEYINPUT7), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(KEYINPUT7), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n508), .A2(G51), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(G63), .A2(G651), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n511), .A2(G89), .B1(new_n510), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(G168));
  NAND2_X1  g100(.A1(new_n511), .A2(G90), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n508), .A2(G52), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n504), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(G301));
  INV_X1    g105(.A(G301), .ZN(G171));
  AOI22_X1  g106(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n504), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT69), .ZN(new_n534));
  AOI22_X1  g109(.A1(G43), .A2(new_n508), .B1(new_n511), .B2(G81), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  NAND4_X1  g113(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT70), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT8), .ZN(new_n542));
  NAND4_X1  g117(.A1(G319), .A2(G483), .A3(G661), .A4(new_n542), .ZN(G188));
  NAND2_X1  g118(.A1(new_n508), .A2(G53), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT9), .ZN(new_n545));
  NAND2_X1  g120(.A1(G78), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(new_n510), .ZN(new_n547));
  XNOR2_X1  g122(.A(KEYINPUT71), .B(G65), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n511), .A2(G91), .B1(G651), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n545), .A2(new_n550), .ZN(G299));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n524), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n521), .A2(new_n523), .A3(KEYINPUT72), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(G286));
  NAND2_X1  g131(.A1(new_n511), .A2(G87), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n511), .A2(KEYINPUT73), .A3(G87), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n510), .A2(G74), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n508), .A2(G49), .B1(G651), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(G288));
  NAND2_X1  g139(.A1(new_n508), .A2(G48), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n511), .A2(G86), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n504), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(G305));
  NAND2_X1  g144(.A1(new_n511), .A2(G85), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n508), .A2(G47), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(new_n504), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(G301), .A2(G868), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n511), .A2(G92), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT10), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n511), .A2(KEYINPUT10), .A3(G92), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(G79), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G66), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n547), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n508), .A2(G54), .B1(G651), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n576), .B1(new_n587), .B2(G868), .ZN(G284));
  OAI21_X1  g163(.A(new_n576), .B1(new_n587), .B2(G868), .ZN(G321));
  NAND2_X1  g164(.A1(new_n555), .A2(G868), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(G868), .B2(G299), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT74), .ZN(G297));
  XOR2_X1   g167(.A(new_n591), .B(KEYINPUT75), .Z(G280));
  INV_X1    g168(.A(G559), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n587), .B1(new_n594), .B2(G860), .ZN(G148));
  NAND2_X1  g170(.A1(new_n587), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G868), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(G868), .B2(new_n537), .ZN(G323));
  XNOR2_X1  g173(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g174(.A1(new_n466), .A2(new_n472), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n481), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT12), .Z(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT13), .ZN(new_n603));
  INV_X1    g178(.A(G2100), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n484), .A2(G123), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n461), .A2(G111), .ZN(new_n608));
  OAI21_X1  g183(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n609));
  INV_X1    g184(.A(G135), .ZN(new_n610));
  OAI221_X1 g185(.A(new_n607), .B1(new_n608), .B2(new_n609), .C1(new_n610), .C2(new_n478), .ZN(new_n611));
  INV_X1    g186(.A(G2096), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n605), .A2(new_n606), .A3(new_n613), .ZN(G156));
  XNOR2_X1  g189(.A(G2427), .B(G2430), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT78), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT77), .B(G2438), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2435), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT14), .ZN(new_n622));
  XOR2_X1   g197(.A(G1341), .B(G1348), .Z(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n622), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2451), .B(G2454), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(G14), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(new_n629), .B2(new_n626), .ZN(G401));
  INV_X1    g206(.A(KEYINPUT18), .ZN(new_n632));
  XOR2_X1   g207(.A(G2084), .B(G2090), .Z(new_n633));
  XNOR2_X1  g208(.A(G2067), .B(G2678), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(KEYINPUT17), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n633), .A2(new_n634), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n632), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(new_n604), .ZN(new_n639));
  XOR2_X1   g214(.A(G2072), .B(G2078), .Z(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n635), .B2(KEYINPUT18), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(new_n612), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n639), .B(new_n642), .ZN(G227));
  XOR2_X1   g218(.A(G1971), .B(G1976), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT19), .ZN(new_n645));
  XOR2_X1   g220(.A(G1956), .B(G2474), .Z(new_n646));
  XOR2_X1   g221(.A(G1961), .B(G1966), .Z(new_n647));
  AND2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT20), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n646), .A2(new_n647), .ZN(new_n651));
  NOR3_X1   g226(.A1(new_n645), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n645), .B2(new_n651), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n654), .B(new_n655), .Z(new_n656));
  XNOR2_X1  g231(.A(G1991), .B(G1996), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1981), .B(G1986), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G229));
  INV_X1    g236(.A(KEYINPUT36), .ZN(new_n662));
  INV_X1    g237(.A(G16), .ZN(new_n663));
  OR2_X1    g238(.A1(G305), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT32), .ZN(new_n665));
  OR2_X1    g240(.A1(G6), .A2(G16), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n665), .B1(new_n664), .B2(new_n666), .ZN(new_n668));
  OAI21_X1  g243(.A(G1981), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n664), .A2(new_n666), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT32), .ZN(new_n671));
  INV_X1    g246(.A(G1981), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n663), .A2(G23), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(G288), .B2(G16), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT33), .B(G1976), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(G166), .A2(G16), .ZN(new_n681));
  OR2_X1    g256(.A1(G16), .A2(G22), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT81), .B(G1971), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT82), .ZN(new_n684));
  AND3_X1   g259(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n681), .B2(new_n682), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n677), .A2(new_n679), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n680), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g264(.A(KEYINPUT83), .B1(new_n675), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n687), .A2(new_n688), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n669), .A2(new_n674), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT83), .ZN(new_n693));
  NAND4_X1  g268(.A1(new_n691), .A2(new_n692), .A3(new_n693), .A4(new_n680), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT34), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n690), .A2(new_n694), .A3(KEYINPUT34), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G25), .ZN(new_n700));
  INV_X1    g275(.A(new_n478), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G131), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT79), .ZN(new_n703));
  OAI21_X1  g278(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n704));
  INV_X1    g279(.A(G107), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(G2105), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n484), .A2(G119), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n703), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n700), .B1(new_n709), .B2(new_n699), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  XOR2_X1   g286(.A(new_n710), .B(new_n711), .Z(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(KEYINPUT80), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(KEYINPUT80), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n663), .A2(G24), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(new_n574), .B2(new_n663), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1986), .ZN(new_n717));
  NOR3_X1   g292(.A1(new_n713), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n697), .A2(new_n698), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n662), .B1(new_n719), .B2(KEYINPUT84), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n697), .A2(new_n721), .A3(new_n718), .A4(new_n698), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n720), .A2(KEYINPUT85), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n697), .A2(new_n662), .A3(new_n718), .A4(new_n698), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT85), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n720), .B2(new_n722), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n663), .A2(G21), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G168), .B2(new_n663), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1966), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n701), .A2(G141), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G129), .B2(new_n484), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT88), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT26), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(new_n699), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n699), .B2(G32), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT27), .B(G1996), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT31), .B(G11), .Z(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT30), .B(G28), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n745), .B1(new_n699), .B2(new_n746), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n744), .B(new_n747), .C1(new_n699), .C2(new_n611), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n663), .A2(G4), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n587), .B2(new_n663), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G1348), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n484), .A2(G128), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n461), .A2(G116), .ZN(new_n753));
  OAI21_X1  g328(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n754));
  INV_X1    g329(.A(G140), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n752), .B1(new_n753), .B2(new_n754), .C1(new_n755), .C2(new_n478), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G29), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n699), .A2(G26), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT28), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G2067), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n742), .B2(new_n743), .ZN(new_n763));
  OR4_X1    g338(.A1(new_n731), .A2(new_n748), .A3(new_n751), .A4(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G171), .A2(new_n663), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G5), .B2(new_n663), .ZN(new_n766));
  INV_X1    g341(.A(G1961), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT89), .Z(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G34), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(G29), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G160), .B2(G29), .ZN(new_n773));
  INV_X1    g348(.A(G2084), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n663), .A2(G20), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT23), .Z(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G299), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1956), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n769), .A2(new_n775), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n663), .A2(G19), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n537), .B2(new_n663), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(G1341), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n699), .A2(G35), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G162), .B2(new_n699), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT91), .B(G2090), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n783), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n766), .A2(new_n767), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n699), .A2(G27), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G164), .B2(new_n699), .ZN(new_n793));
  INV_X1    g368(.A(G2078), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT86), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT25), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n701), .A2(G139), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n466), .A2(new_n472), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n800), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n798), .B(new_n799), .C1(new_n801), .C2(new_n461), .ZN(new_n802));
  MUX2_X1   g377(.A(G33), .B(new_n802), .S(G29), .Z(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(G2072), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(G2072), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n791), .A2(new_n795), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n764), .A2(new_n780), .A3(new_n790), .A4(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n724), .A2(new_n728), .A3(new_n808), .ZN(G311));
  AND2_X1   g384(.A1(new_n720), .A2(new_n722), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n723), .B(new_n807), .C1(new_n810), .C2(new_n727), .ZN(G150));
  XOR2_X1   g386(.A(KEYINPUT92), .B(G93), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n511), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n508), .A2(G55), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(new_n504), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G860), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  NOR2_X1   g394(.A1(new_n586), .A2(new_n594), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n536), .A2(new_n817), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n814), .A2(new_n816), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n823), .A2(new_n535), .A3(new_n534), .A4(new_n813), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n821), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT39), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT93), .ZN(new_n830));
  INV_X1    g405(.A(G860), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n827), .B2(new_n828), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n819), .B1(new_n830), .B2(new_n832), .ZN(G145));
  XOR2_X1   g408(.A(new_n756), .B(new_n502), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n802), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n739), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n709), .B(new_n602), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n484), .A2(G130), .ZN(new_n838));
  OR2_X1    g413(.A1(G106), .A2(G2105), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n839), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n840));
  INV_X1    g415(.A(G142), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n838), .B(new_n840), .C1(new_n841), .C2(new_n478), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n837), .B(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n836), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n836), .A2(new_n843), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n844), .A2(KEYINPUT94), .A3(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(G160), .B(new_n611), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G162), .ZN(new_n848));
  OR3_X1    g423(.A1(new_n836), .A2(KEYINPUT94), .A3(new_n843), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(G37), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n844), .A2(new_n845), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n850), .B(new_n851), .C1(new_n848), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g429(.A(new_n826), .B(new_n596), .ZN(new_n855));
  NAND2_X1  g430(.A1(G299), .A2(new_n586), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n545), .A2(new_n581), .A3(new_n550), .A4(new_n585), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n856), .A2(KEYINPUT41), .A3(new_n857), .ZN(new_n861));
  AOI21_X1  g436(.A(KEYINPUT41), .B1(new_n856), .B2(new_n857), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n860), .B1(new_n855), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT95), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n561), .A2(new_n574), .A3(new_n563), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n574), .B1(new_n561), .B2(new_n563), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(G288), .A2(G290), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(KEYINPUT95), .A3(new_n867), .ZN(new_n872));
  XNOR2_X1  g447(.A(G303), .B(G305), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n873), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n875), .B(new_n866), .C1(new_n869), .C2(new_n868), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT42), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n865), .B(new_n878), .ZN(new_n879));
  MUX2_X1   g454(.A(new_n817), .B(new_n879), .S(G868), .Z(G295));
  MUX2_X1   g455(.A(new_n817), .B(new_n879), .S(G868), .Z(G331));
  INV_X1    g456(.A(new_n554), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT72), .B1(new_n521), .B2(new_n523), .ZN(new_n883));
  OAI21_X1  g458(.A(G171), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n524), .A2(G301), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n884), .A2(new_n822), .A3(new_n824), .A4(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(G301), .B1(new_n553), .B2(new_n554), .ZN(new_n887));
  INV_X1    g462(.A(new_n885), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n825), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n886), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n826), .A2(KEYINPUT97), .A3(new_n884), .A4(new_n885), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n858), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n874), .A2(new_n876), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n886), .A2(new_n889), .A3(KEYINPUT96), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT96), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n825), .B(new_n897), .C1(new_n887), .C2(new_n888), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n863), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n851), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n863), .A2(new_n896), .A3(new_n898), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT98), .B1(new_n903), .B2(new_n893), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT98), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n894), .A2(new_n905), .A3(new_n899), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT99), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n874), .A2(new_n907), .A3(new_n876), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n907), .B1(new_n874), .B2(new_n876), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n904), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n902), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT43), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n863), .A2(new_n891), .A3(new_n892), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n896), .A2(new_n898), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n915), .B1(new_n916), .B2(new_n858), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n910), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n918), .B1(new_n917), .B2(new_n910), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n902), .B(new_n914), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n913), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n917), .A2(new_n910), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT100), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n901), .B1(new_n927), .B2(new_n919), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n925), .B1(new_n928), .B2(new_n914), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n902), .B1(new_n920), .B2(new_n921), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n930), .A2(KEYINPUT101), .A3(KEYINPUT43), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n902), .A2(new_n911), .A3(new_n914), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n924), .B1(new_n933), .B2(KEYINPUT44), .ZN(G397));
  NOR2_X1   g509(.A1(G290), .A2(G1986), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT103), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(G1986), .B2(G290), .ZN(new_n937));
  INV_X1    g512(.A(G1996), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n739), .B(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n756), .B(new_n761), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n709), .B(new_n711), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT104), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n937), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n473), .A2(new_n474), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(new_n476), .A3(new_n462), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(G2105), .ZN(new_n947));
  INV_X1    g522(.A(G40), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n482), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(KEYINPUT102), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT102), .ZN(new_n951));
  INV_X1    g526(.A(new_n949), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n477), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G1384), .B1(new_n496), .B2(new_n501), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n954), .A2(KEYINPUT45), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n944), .A2(new_n956), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n950), .A2(new_n953), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n959));
  INV_X1    g534(.A(G1384), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n502), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT105), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n502), .A2(new_n960), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT50), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n955), .A2(new_n965), .A3(new_n959), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n962), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n958), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n962), .A2(new_n964), .A3(new_n966), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT115), .B1(new_n954), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n767), .A3(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n955), .B(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(new_n953), .A3(new_n950), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n973), .B1(new_n976), .B2(G2078), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n972), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n794), .A2(KEYINPUT53), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n978), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(G171), .ZN(new_n981));
  INV_X1    g556(.A(G8), .ZN(new_n982));
  NOR2_X1   g557(.A1(G168), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(G1966), .B1(new_n958), .B2(new_n975), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n954), .A2(new_n970), .A3(G2084), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT119), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n954), .A2(new_n970), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n774), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT119), .ZN(new_n990));
  INV_X1    g565(.A(G1966), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n976), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n984), .B1(new_n987), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n987), .A2(new_n993), .A3(G168), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n996), .A2(KEYINPUT120), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(KEYINPUT120), .ZN(new_n998));
  OAI21_X1  g573(.A(G8), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n995), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n989), .A2(new_n992), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G8), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n983), .A2(KEYINPUT51), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n994), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT62), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n981), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT124), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1010));
  INV_X1    g585(.A(G2090), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n988), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1971), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n976), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n982), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT106), .B(KEYINPUT55), .Z(new_n1016));
  AND3_X1   g591(.A1(G303), .A2(G8), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT106), .ZN(new_n1018));
  AOI22_X1  g593(.A1(G303), .A2(G8), .B1(new_n1018), .B2(KEYINPUT55), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1015), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n950), .A2(new_n953), .A3(new_n961), .A4(new_n964), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1014), .B1(G2090), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(new_n1023), .B2(G8), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1976), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G288), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1026), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n950), .A2(new_n953), .A3(new_n955), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT107), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1030), .A2(new_n1031), .A3(G8), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n1030), .B2(G8), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1028), .B(new_n1029), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G305), .A2(G1981), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n565), .A2(new_n566), .A3(new_n672), .A4(new_n568), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1036), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1039));
  OAI22_X1  g614(.A1(new_n1032), .A2(new_n1033), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1034), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1030), .A2(G8), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT107), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1030), .A2(new_n1031), .A3(G8), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n1028), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT52), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1041), .A2(new_n1047), .A3(KEYINPUT109), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1027), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1034), .B(new_n1040), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT109), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1025), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n995), .A2(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT124), .B(KEYINPUT62), .C1(new_n1055), .C2(new_n994), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1008), .A2(new_n1010), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT108), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT108), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1051), .A2(new_n1059), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1040), .A2(new_n1026), .A3(new_n561), .A4(new_n563), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1037), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1061), .A2(new_n1021), .B1(new_n1045), .B2(new_n1063), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT56), .B(G2072), .Z(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n975), .A2(new_n953), .A3(new_n950), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1067), .A2(KEYINPUT113), .ZN(new_n1071));
  INV_X1    g646(.A(G1956), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1022), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n545), .A2(new_n1075), .A3(new_n550), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1075), .B1(new_n545), .B2(new_n550), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1074), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1348), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n969), .A2(new_n971), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n958), .A2(new_n761), .A3(new_n955), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1080), .B1(new_n1084), .B2(new_n586), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1070), .A2(new_n1078), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1068), .A2(new_n1069), .B1(new_n1072), .B2(new_n1022), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1089), .A2(KEYINPUT114), .A3(new_n1078), .A4(new_n1071), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1085), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT60), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1093), .B1(new_n587), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1082), .A2(new_n1083), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT60), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n586), .A2(KEYINPUT117), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1096), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1084), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1100), .A2(new_n1101), .A3(KEYINPUT118), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT118), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT61), .B1(new_n1091), .B2(new_n1080), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1080), .A2(KEYINPUT61), .A3(new_n1086), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT58), .B(G1341), .Z(new_n1108));
  NAND2_X1  g683(.A1(new_n1030), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n975), .A2(new_n938), .A3(new_n953), .A4(new_n950), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n536), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1107), .B1(new_n1111), .B2(KEYINPUT116), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(KEYINPUT116), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1111), .A2(KEYINPUT116), .A3(new_n1107), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1106), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1105), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1092), .B1(new_n1104), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1006), .ZN(new_n1119));
  XOR2_X1   g694(.A(G301), .B(KEYINPUT54), .Z(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n477), .A2(new_n952), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1122), .A2(KEYINPUT122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(KEYINPUT122), .ZN(new_n1124));
  INV_X1    g699(.A(new_n979), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1123), .A2(new_n975), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1120), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n1127), .B2(new_n1126), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n980), .A2(new_n1121), .B1(new_n978), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1054), .A2(new_n1119), .A3(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1057), .B(new_n1064), .C1(new_n1118), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT111), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1017), .A2(new_n1019), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1015), .A2(new_n1135), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n982), .B(new_n1134), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1002), .A2(KEYINPUT63), .A3(G8), .A4(new_n555), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT112), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT112), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1142), .B(new_n1139), .C1(new_n1058), .C2(new_n1060), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1003), .A2(G286), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1148), .A2(KEYINPUT110), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT63), .B1(new_n1148), .B2(KEYINPUT110), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1144), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n957), .B1(new_n1132), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n956), .ZN(new_n1153));
  OR3_X1    g728(.A1(new_n1153), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT46), .B1(new_n1153), .B2(G1996), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n740), .A2(new_n940), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1154), .A2(new_n1155), .B1(new_n956), .B2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g732(.A(new_n1157), .B(KEYINPUT47), .Z(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT48), .B1(new_n936), .B2(new_n956), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n943), .A2(new_n941), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n1160), .B2(new_n956), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n936), .A2(KEYINPUT48), .A3(new_n956), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n709), .A2(new_n711), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(KEYINPUT125), .Z(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n941), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(G2067), .B2(new_n756), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1161), .A2(new_n1162), .B1(new_n956), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1158), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT126), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1152), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g745(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1172));
  NAND2_X1  g746(.A1(new_n660), .A2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g747(.A(new_n1173), .B(KEYINPUT127), .Z(new_n1174));
  NAND2_X1  g748(.A1(new_n913), .A2(new_n922), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n1174), .A2(new_n853), .A3(new_n1175), .ZN(G225));
  INV_X1    g750(.A(G225), .ZN(G308));
endmodule


