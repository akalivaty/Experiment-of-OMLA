//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968;
  XOR2_X1   g000(.A(G155gat), .B(G162gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G141gat), .B(G148gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT79), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT80), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G155gat), .B(G162gat), .ZN(new_n209));
  INV_X1    g008(.A(G155gat), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT2), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G141gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT80), .A3(G148gat), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n208), .A2(new_n209), .A3(new_n212), .A4(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n202), .B(new_n216), .C1(new_n203), .C2(new_n204), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n206), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G197gat), .B(G204gat), .ZN(new_n219));
  INV_X1    g018(.A(G211gat), .ZN(new_n220));
  INV_X1    g019(.A(G218gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n219), .B1(KEYINPUT22), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G211gat), .B(G218gat), .Z(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT29), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n218), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G228gat), .ZN(new_n230));
  INV_X1    g029(.A(G233gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n206), .A2(new_n228), .A3(new_n215), .A4(new_n217), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n225), .B1(new_n233), .B2(new_n226), .ZN(new_n234));
  OR3_X1    g033(.A1(new_n229), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  OAI211_X1 g034(.A(G228gat), .B(G233gat), .C1(new_n229), .C2(new_n234), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT31), .B(G50gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n238), .B1(new_n235), .B2(new_n236), .ZN(new_n241));
  XOR2_X1   g040(.A(G78gat), .B(G106gat), .Z(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT85), .B(G22gat), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n242), .B(new_n243), .Z(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n240), .A2(new_n241), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n235), .A2(new_n236), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n237), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n244), .B1(new_n248), .B2(new_n239), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G1gat), .B(G29gat), .ZN(new_n251));
  INV_X1    g050(.A(G85gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT0), .B(G57gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n253), .B(new_n254), .Z(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT83), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n258));
  INV_X1    g057(.A(G120gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G113gat), .ZN(new_n260));
  INV_X1    g059(.A(G113gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G120gat), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT1), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G127gat), .B(G134gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n261), .A2(KEYINPUT73), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n261), .A2(KEYINPUT73), .ZN(new_n267));
  OAI21_X1  g066(.A(G120gat), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT1), .B1(new_n268), .B2(new_n260), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n265), .B1(new_n269), .B2(new_n264), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n258), .B1(new_n218), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n206), .A2(new_n215), .A3(new_n217), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT73), .B(G113gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n260), .B1(new_n273), .B2(new_n259), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n275), .A3(new_n264), .ZN(new_n276));
  INV_X1    g075(.A(new_n265), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n272), .A2(new_n278), .A3(KEYINPUT4), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n257), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n218), .A2(new_n258), .A3(new_n270), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT4), .B1(new_n272), .B2(new_n278), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(KEYINPUT83), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G225gat), .A2(G233gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT81), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(new_n218), .B2(new_n228), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n272), .A2(KEYINPUT81), .A3(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n233), .A2(new_n278), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n286), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n284), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n272), .A2(KEYINPUT81), .A3(KEYINPUT3), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT81), .B1(new_n272), .B2(KEYINPUT3), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n291), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n298), .A3(new_n285), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n270), .A2(new_n215), .A3(new_n206), .A4(new_n217), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n272), .A2(new_n278), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n285), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT82), .B1(new_n302), .B2(new_n293), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n272), .A2(new_n278), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n272), .A2(new_n278), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n286), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT82), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT5), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n299), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n256), .B1(new_n294), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT6), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT84), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n294), .A2(new_n309), .A3(new_n256), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(new_n310), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT6), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NOR4_X1   g115(.A1(new_n313), .A2(new_n310), .A3(KEYINPUT84), .A4(KEYINPUT6), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n311), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT28), .ZN(new_n319));
  INV_X1    g118(.A(G190gat), .ZN(new_n320));
  AND2_X1   g119(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n325), .B1(new_n323), .B2(new_n324), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n319), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G169gat), .ZN(new_n329));
  INV_X1    g128(.A(G176gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT26), .ZN(new_n331));
  NAND2_X1  g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT26), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n333), .B1(G169gat), .B2(G176gat), .ZN(new_n334));
  AND2_X1   g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n331), .B(new_n332), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT72), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n329), .A2(new_n330), .ZN(new_n338));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n333), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n340), .A2(new_n341), .A3(new_n332), .A4(new_n331), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  OR2_X1    g142(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n345));
  AOI21_X1  g144(.A(G190gat), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT71), .B1(new_n346), .B2(KEYINPUT70), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(KEYINPUT28), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n328), .A2(new_n343), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G183gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n320), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT69), .B1(G183gat), .B2(G190gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT24), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n354), .ZN(new_n355));
  OAI221_X1 g154(.A(new_n352), .B1(new_n353), .B2(new_n354), .C1(new_n355), .C2(KEYINPUT69), .ZN(new_n356));
  INV_X1    g155(.A(new_n338), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n335), .B1(new_n357), .B2(KEYINPUT23), .ZN(new_n358));
  AND2_X1   g157(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n359));
  NOR2_X1   g158(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n338), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT68), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT68), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n338), .B(new_n363), .C1(new_n359), .C2(new_n360), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n356), .A2(new_n358), .A3(new_n362), .A4(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT25), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT66), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n332), .A2(new_n354), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n369), .B1(new_n351), .B2(new_n320), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT25), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n371), .A2(new_n358), .A3(new_n362), .A4(new_n364), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n350), .A2(new_n366), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n226), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n350), .A2(new_n372), .A3(new_n374), .A4(new_n366), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n225), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT75), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n376), .A2(new_n225), .A3(new_n377), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n378), .A2(KEYINPUT75), .A3(new_n379), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G8gat), .B(G36gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(G64gat), .B(G92gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT77), .B(KEYINPUT30), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(new_n385), .B2(new_n389), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n382), .A2(new_n381), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n225), .B1(new_n376), .B2(new_n377), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n384), .ZN(new_n396));
  OAI211_X1 g195(.A(KEYINPUT30), .B(new_n389), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT76), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n388), .B1(new_n383), .B2(new_n384), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(KEYINPUT76), .A3(KEYINPUT30), .ZN(new_n401));
  AOI211_X1 g200(.A(new_n390), .B(new_n392), .C1(new_n399), .C2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n250), .B1(new_n318), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n373), .A2(new_n270), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n350), .A2(new_n372), .A3(new_n278), .A4(new_n366), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(G227gat), .A2(G233gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n407), .B(KEYINPUT64), .Z(new_n408));
  XOR2_X1   g207(.A(new_n408), .B(KEYINPUT65), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT32), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n412), .B1(new_n406), .B2(new_n410), .ZN(new_n413));
  XNOR2_X1  g212(.A(G15gat), .B(G43gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G71gat), .B(G99gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  NAND3_X1  g215(.A1(new_n411), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n416), .ZN(new_n418));
  OAI221_X1 g217(.A(KEYINPUT32), .B1(new_n412), .B2(new_n418), .C1(new_n406), .C2(new_n410), .ZN(new_n419));
  INV_X1    g218(.A(new_n408), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n406), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n409), .A2(KEYINPUT34), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n421), .A2(KEYINPUT34), .B1(new_n406), .B2(new_n422), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n417), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n423), .B1(new_n417), .B2(new_n419), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n426), .A2(KEYINPUT36), .ZN(new_n427));
  AOI211_X1 g226(.A(KEYINPUT74), .B(new_n423), .C1(new_n419), .C2(new_n417), .ZN(new_n428));
  INV_X1    g227(.A(new_n423), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n417), .A2(new_n419), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT74), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n427), .B1(new_n433), .B2(KEYINPUT36), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n403), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n285), .B1(new_n284), .B2(new_n297), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT39), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n255), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n304), .A2(new_n305), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n437), .B1(new_n439), .B2(new_n285), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n440), .B(KEYINPUT86), .Z(new_n441));
  OAI21_X1  g240(.A(new_n438), .B1(new_n441), .B2(new_n436), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT40), .ZN(new_n443));
  INV_X1    g242(.A(new_n392), .ZN(new_n444));
  INV_X1    g243(.A(new_n390), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n397), .A2(new_n398), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT76), .B1(new_n400), .B2(KEYINPUT30), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n444), .B(new_n445), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n294), .A2(new_n309), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n255), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n443), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n294), .A2(new_n309), .A3(new_n256), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n315), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n311), .ZN(new_n454));
  INV_X1    g253(.A(new_n400), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT37), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n389), .B1(new_n385), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n383), .A2(KEYINPUT37), .A3(new_n384), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n457), .A2(KEYINPUT38), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n380), .A2(KEYINPUT87), .A3(new_n382), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n460), .B(KEYINPUT37), .C1(KEYINPUT87), .C2(new_n380), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT38), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n455), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n451), .B(new_n250), .C1(new_n454), .C2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n246), .A2(new_n249), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n428), .A2(new_n432), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n318), .A2(new_n402), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT35), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT35), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n454), .A2(new_n426), .A3(new_n469), .A4(new_n250), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(new_n448), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n435), .A2(new_n464), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT17), .ZN(new_n474));
  OR3_X1    g273(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G29gat), .A2(G36gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G50gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G43gat), .ZN(new_n482));
  INV_X1    g281(.A(G43gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G50gat), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n482), .A2(new_n484), .A3(KEYINPUT88), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT88), .B1(new_n482), .B2(new_n484), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G43gat), .B(G50gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n489), .A2(KEYINPUT15), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n480), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(KEYINPUT88), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n483), .A2(G50gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n481), .A2(G43gat), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n492), .A2(new_n496), .A3(KEYINPUT15), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n479), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n474), .B1(new_n499), .B2(KEYINPUT89), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n488), .A2(new_n480), .ZN(new_n501));
  INV_X1    g300(.A(new_n490), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n479), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT89), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT17), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G15gat), .B(G22gat), .ZN(new_n508));
  INV_X1    g307(.A(G1gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(KEYINPUT16), .A3(new_n509), .ZN(new_n510));
  OAI221_X1 g309(.A(new_n510), .B1(KEYINPUT90), .B2(G8gat), .C1(new_n509), .C2(new_n508), .ZN(new_n511));
  NAND2_X1  g310(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n511), .B(new_n512), .Z(new_n513));
  NAND2_X1  g312(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n513), .A2(new_n499), .ZN(new_n515));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(KEYINPUT91), .A2(KEYINPUT18), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n513), .B(new_n499), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(new_n516), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n517), .A2(new_n518), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n519), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  INV_X1    g325(.A(G197gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT11), .B(G169gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT12), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n531), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n519), .A2(new_n523), .A3(new_n524), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT8), .ZN(new_n540));
  NAND2_X1  g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT7), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G92gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n252), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n540), .A2(new_n543), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G99gat), .B(G106gat), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT97), .ZN(new_n550));
  AOI22_X1  g349(.A1(KEYINPUT8), .A2(new_n539), .B1(new_n252), .B2(new_n544), .ZN(new_n551));
  XNOR2_X1  g350(.A(G99gat), .B(G106gat), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n551), .A2(new_n552), .A3(new_n543), .A4(new_n546), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  OR3_X1    g353(.A1(new_n547), .A2(new_n550), .A3(new_n548), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n538), .B1(new_n507), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n499), .A2(new_n556), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n320), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n554), .A2(new_n555), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n500), .B2(new_n506), .ZN(new_n562));
  NOR4_X1   g361(.A1(new_n562), .A2(G190gat), .A3(new_n538), .A4(new_n558), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n221), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT17), .B1(new_n504), .B2(new_n505), .ZN(new_n566));
  NOR4_X1   g365(.A1(new_n501), .A2(new_n503), .A3(KEYINPUT89), .A4(new_n474), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n556), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n537), .A3(new_n559), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(G190gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n557), .A2(new_n320), .A3(new_n559), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n571), .A3(G218gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n564), .A2(new_n565), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n574), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n564), .A2(new_n572), .A3(new_n565), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n575), .A2(new_n577), .A3(new_n579), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G127gat), .B(G155gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT93), .ZN(new_n589));
  NOR2_X1   g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n588), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n592), .A2(KEYINPUT9), .ZN(new_n593));
  XNOR2_X1  g392(.A(G57gat), .B(G64gat), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n589), .B(new_n591), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G57gat), .B(G64gat), .Z(new_n596));
  INV_X1    g395(.A(KEYINPUT94), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(KEYINPUT94), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n592), .A2(KEYINPUT9), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n591), .A2(new_n602), .A3(new_n588), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT95), .B1(new_n592), .B2(new_n590), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n595), .B1(new_n600), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n513), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G183gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(new_n220), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n612), .A2(new_n614), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n587), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(new_n586), .A3(new_n615), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n605), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n594), .B(new_n597), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g423(.A1(new_n624), .A2(new_n595), .B1(new_n554), .B2(new_n555), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n549), .A2(new_n553), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n606), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT98), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n625), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n561), .A2(new_n606), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n624), .A2(new_n626), .A3(new_n595), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT10), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT10), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n556), .A2(new_n638), .A3(new_n606), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n631), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n632), .A2(new_n633), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n634), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT100), .ZN(new_n644));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  NOR2_X1   g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n642), .A2(new_n646), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n583), .A2(new_n621), .A3(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n473), .A2(new_n536), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n318), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n448), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n653), .A2(KEYINPUT101), .A3(new_n448), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT16), .B(G8gat), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n659), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(new_n662), .B2(G8gat), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n665), .B1(new_n657), .B2(new_n666), .ZN(G1325gat));
  AOI21_X1  g466(.A(G15gat), .B1(new_n653), .B2(new_n426), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n434), .A2(G15gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT102), .Z(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n653), .B2(new_n670), .ZN(G1326gat));
  NAND2_X1  g470(.A1(new_n653), .A2(new_n465), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT103), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT43), .B(G22gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n673), .B(new_n674), .Z(G1327gat));
  NOR2_X1   g474(.A1(new_n473), .A2(new_n536), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677));
  INV_X1    g476(.A(new_n621), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n651), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n679), .B2(new_n583), .ZN(new_n680));
  INV_X1    g479(.A(new_n679), .ZN(new_n681));
  INV_X1    g480(.A(new_n583), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(KEYINPUT104), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n676), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n684), .A2(G29gat), .A3(new_n318), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT45), .Z(new_n686));
  NAND2_X1  g485(.A1(new_n435), .A2(new_n464), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n688));
  AOI211_X1 g487(.A(new_n688), .B(new_n471), .C1(KEYINPUT35), .C2(new_n467), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT105), .B1(new_n468), .B2(new_n472), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n687), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n682), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT44), .B1(new_n473), .B2(new_n583), .ZN(new_n694));
  AOI211_X1 g493(.A(new_n536), .B(new_n679), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n654), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G29gat), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n686), .A2(new_n697), .ZN(G1328gat));
  NAND2_X1  g497(.A1(new_n695), .A2(new_n448), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n695), .A2(KEYINPUT108), .A3(new_n448), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(G36gat), .A3(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n684), .A2(G36gat), .A3(new_n402), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n704), .B1(KEYINPUT107), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n703), .A2(new_n706), .A3(new_n708), .ZN(G1329gat));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n483), .B1(new_n695), .B2(new_n434), .ZN(new_n711));
  INV_X1    g510(.A(new_n426), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n684), .A2(G43gat), .A3(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n710), .B(KEYINPUT47), .C1(new_n711), .C2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n693), .A2(new_n694), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n716), .A2(new_n434), .A3(new_n535), .A4(new_n681), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n713), .B1(new_n717), .B2(G43gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n715), .B1(new_n718), .B2(KEYINPUT109), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n714), .A2(new_n719), .ZN(G1330gat));
  NAND3_X1  g519(.A1(new_n695), .A2(G50gat), .A3(new_n465), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n481), .B1(new_n684), .B2(new_n250), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n723), .B1(new_n721), .B2(new_n722), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(G1331gat));
  AND2_X1   g525(.A1(new_n691), .A2(new_n536), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n583), .A2(new_n621), .A3(new_n650), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n654), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g532(.A1(new_n730), .A2(new_n402), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  AND2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n734), .B2(new_n735), .ZN(G1333gat));
  INV_X1    g537(.A(G71gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n730), .B2(new_n712), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n727), .A2(G71gat), .A3(new_n729), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n742), .B2(new_n434), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n727), .A2(G71gat), .A3(new_n729), .ZN(new_n744));
  INV_X1    g543(.A(new_n434), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n744), .A2(KEYINPUT111), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n740), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT50), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n749), .B(new_n740), .C1(new_n743), .C2(new_n746), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(G1334gat));
  NAND2_X1  g550(.A1(new_n731), .A2(new_n465), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g552(.A1(new_n621), .A2(new_n535), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n716), .A2(new_n650), .A3(new_n754), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n755), .A2(new_n252), .A3(new_n318), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n691), .A2(new_n682), .A3(new_n754), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(KEYINPUT112), .A3(new_n760), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n760), .A2(KEYINPUT112), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n761), .A2(new_n762), .A3(new_n654), .A4(new_n650), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n756), .B1(new_n763), .B2(new_n252), .ZN(G1336gat));
  NOR2_X1   g563(.A1(new_n402), .A2(G92gat), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n761), .A2(new_n762), .A3(new_n650), .A4(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n716), .A2(new_n448), .A3(new_n650), .A4(new_n754), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(new_n767), .B2(G92gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n651), .B1(new_n759), .B2(new_n760), .ZN(new_n771));
  AOI22_X1  g570(.A1(new_n771), .A2(new_n765), .B1(new_n767), .B2(G92gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n770), .B2(new_n772), .ZN(G1337gat));
  OR3_X1    g572(.A1(new_n755), .A2(KEYINPUT113), .A3(new_n745), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT114), .B(G99gat), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT113), .B1(new_n755), .B2(new_n745), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n712), .A2(new_n775), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n761), .A2(new_n762), .A3(new_n650), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1338gat));
  NOR2_X1   g579(.A1(new_n250), .A2(G106gat), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n761), .A2(new_n762), .A3(new_n650), .A4(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n716), .A2(new_n465), .A3(new_n650), .A4(new_n754), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT53), .B1(new_n783), .B2(G106gat), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n771), .A2(new_n781), .B1(new_n783), .B2(G106gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(G1339gat));
  OAI21_X1  g587(.A(new_n638), .B1(new_n625), .B2(new_n628), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n607), .A2(new_n561), .A3(KEYINPUT10), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n630), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n640), .A2(new_n791), .A3(KEYINPUT54), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT115), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n640), .A2(new_n791), .A3(new_n794), .A4(KEYINPUT54), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n646), .B1(new_n640), .B2(KEYINPUT54), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(KEYINPUT55), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n648), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n797), .B1(new_n793), .B2(new_n795), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(KEYINPUT55), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT116), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n801), .A2(KEYINPUT55), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n647), .B1(new_n801), .B2(KEYINPUT55), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n803), .A2(new_n535), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n520), .A2(new_n522), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n516), .B1(new_n514), .B2(new_n515), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n530), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n534), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n650), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n808), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n583), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n803), .A2(new_n807), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n817), .A2(new_n582), .A3(new_n581), .A4(new_n813), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n621), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n583), .A2(new_n621), .A3(new_n536), .A4(new_n651), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT117), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823));
  INV_X1    g622(.A(new_n582), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n579), .B1(new_n575), .B2(new_n577), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n824), .A2(new_n825), .A3(new_n812), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n826), .A2(new_n817), .B1(new_n815), .B2(new_n583), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n823), .B(new_n820), .C1(new_n827), .C2(new_n621), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n822), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n466), .ZN(new_n830));
  NOR4_X1   g629(.A1(new_n829), .A2(new_n318), .A3(new_n448), .A4(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n831), .B(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n833), .B(new_n535), .C1(new_n266), .C2(new_n267), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n822), .A2(new_n828), .A3(new_n250), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n318), .A2(new_n448), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n822), .A2(new_n828), .A3(KEYINPUT118), .A4(new_n250), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n837), .A2(new_n426), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G113gat), .B1(new_n840), .B2(new_n536), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n834), .A2(new_n841), .ZN(G1340gat));
  NAND3_X1  g641(.A1(new_n833), .A2(new_n259), .A3(new_n650), .ZN(new_n843));
  OAI21_X1  g642(.A(G120gat), .B1(new_n840), .B2(new_n651), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1341gat));
  INV_X1    g644(.A(G127gat), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n840), .A2(new_n846), .A3(new_n678), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n621), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n848), .B(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n847), .B1(new_n850), .B2(new_n846), .ZN(G1342gat));
  INV_X1    g650(.A(G134gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n831), .A2(new_n852), .A3(new_n682), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n853), .A2(KEYINPUT56), .ZN(new_n854));
  OAI21_X1  g653(.A(G134gat), .B1(new_n840), .B2(new_n583), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(KEYINPUT56), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(G1343gat));
  NAND2_X1  g656(.A1(new_n745), .A2(new_n838), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n822), .A2(new_n828), .A3(new_n465), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n800), .B1(KEYINPUT121), .B2(new_n802), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n802), .A2(KEYINPUT121), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n535), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n814), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT122), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n864), .A2(new_n867), .A3(new_n814), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n583), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n621), .B1(new_n869), .B2(new_n818), .ZN(new_n870));
  OAI211_X1 g669(.A(KEYINPUT57), .B(new_n465), .C1(new_n870), .C2(new_n821), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n858), .B1(new_n861), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n213), .B1(new_n872), .B2(new_n535), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n858), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(G141gat), .A3(new_n536), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n874), .A2(new_n875), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT58), .B1(new_n873), .B2(new_n878), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1344gat));
  AOI21_X1  g681(.A(G148gat), .B1(new_n876), .B2(new_n650), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT59), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n859), .A2(KEYINPUT57), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n826), .A2(new_n805), .A3(new_n804), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n621), .B1(new_n869), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n860), .B(new_n465), .C1(new_n888), .C2(new_n821), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n858), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n890), .A2(KEYINPUT59), .A3(new_n650), .A4(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n872), .A2(new_n650), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(KEYINPUT59), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n885), .B1(new_n894), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g694(.A(new_n210), .B1(new_n877), .B2(new_n678), .ZN(new_n896));
  INV_X1    g695(.A(new_n872), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n621), .A2(G155gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n896), .B(KEYINPUT123), .C1(new_n897), .C2(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1346gat));
  AOI21_X1  g702(.A(G162gat), .B1(new_n876), .B2(new_n682), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n583), .A2(new_n211), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n872), .B2(new_n905), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n654), .A2(new_n402), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n837), .A2(new_n426), .A3(new_n839), .A4(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(G169gat), .B1(new_n908), .B2(new_n536), .ZN(new_n909));
  INV_X1    g708(.A(new_n907), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n829), .A2(new_n830), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n329), .A3(new_n535), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n912), .ZN(G1348gat));
  OAI21_X1  g712(.A(G176gat), .B1(new_n908), .B2(new_n651), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n330), .A3(new_n650), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT124), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n914), .A2(new_n918), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1349gat));
  AND3_X1   g719(.A1(new_n822), .A2(new_n828), .A3(new_n466), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n344), .A2(new_n345), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n921), .A2(new_n922), .A3(new_n621), .A4(new_n907), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n911), .A2(new_n925), .A3(new_n922), .A4(new_n621), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G183gat), .B1(new_n908), .B2(new_n678), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT60), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT60), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1350gat));
  OAI21_X1  g732(.A(G190gat), .B1(new_n908), .B2(new_n583), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT61), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n936), .B(G190gat), .C1(new_n908), .C2(new_n583), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n911), .A2(new_n320), .A3(new_n682), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1351gat));
  NOR2_X1   g739(.A1(new_n910), .A2(new_n434), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n886), .A2(new_n889), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n536), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n859), .A2(new_n434), .A3(new_n910), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n527), .A3(new_n535), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1352gat));
  INV_X1    g745(.A(new_n944), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n947), .A2(G204gat), .A3(new_n651), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n890), .A2(new_n650), .A3(new_n941), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G204gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(G1353gat));
  NAND4_X1  g753(.A1(new_n886), .A2(new_n621), .A3(new_n889), .A4(new_n941), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G211gat), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n955), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n958), .A2(KEYINPUT126), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n220), .A3(new_n621), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n956), .A2(new_n962), .A3(new_n957), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(G1354gat));
  NAND3_X1  g763(.A1(new_n944), .A2(new_n221), .A3(new_n682), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n942), .A2(KEYINPUT127), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n942), .A2(KEYINPUT127), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n966), .A2(new_n967), .A3(new_n583), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n965), .B1(new_n968), .B2(new_n221), .ZN(G1355gat));
endmodule


