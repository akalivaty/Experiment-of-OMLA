//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n543, new_n544,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n557, new_n558, new_n559, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT66), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT67), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT68), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT69), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G221), .A3(G218), .A4(G220), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT70), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT71), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n463), .A2(G137), .A3(new_n462), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n462), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n476), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n462), .A2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n478), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT72), .ZN(G162));
  NAND4_X1  g059(.A1(new_n473), .A2(new_n475), .A3(G126), .A4(G2105), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(new_n488), .A3(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n473), .A2(new_n475), .A3(G138), .A4(new_n462), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n463), .A2(new_n493), .A3(G138), .A4(new_n462), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(G164));
  XNOR2_X1  g070(.A(KEYINPUT5), .B(G543), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n496), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n497));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT73), .A2(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT6), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT73), .A3(G651), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n501), .A2(new_n503), .A3(G50), .A4(G543), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n501), .A2(new_n503), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n499), .A2(new_n511), .ZN(G166));
  NAND3_X1  g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT7), .ZN(new_n514));
  INV_X1    g089(.A(G89), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n501), .A2(new_n503), .A3(G51), .A4(G543), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n506), .A2(new_n508), .A3(G63), .A4(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n517), .A2(KEYINPUT74), .A3(new_n518), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n516), .B1(new_n521), .B2(new_n522), .ZN(G168));
  NAND4_X1  g098(.A1(new_n496), .A2(G90), .A3(new_n501), .A4(new_n503), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n501), .A2(new_n503), .A3(G52), .A4(G543), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT75), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n506), .A2(new_n508), .A3(G64), .ZN(new_n528));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n528), .A2(new_n527), .A3(new_n529), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G651), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n526), .B1(new_n530), .B2(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  NAND4_X1  g109(.A1(new_n496), .A2(G81), .A3(new_n501), .A4(new_n503), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n501), .A2(new_n503), .A3(G43), .A4(G543), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n496), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n535), .B(new_n536), .C1(new_n537), .C2(new_n498), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G860), .ZN(G153));
  AND3_X1   g115(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G36), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n544), .ZN(G188));
  INV_X1    g120(.A(new_n509), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G91), .ZN(new_n547));
  NAND2_X1  g122(.A1(G78), .A2(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n506), .A2(new_n508), .ZN(new_n549));
  INV_X1    g124(.A(G65), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G651), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n501), .A2(new_n503), .A3(G53), .A4(G543), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n547), .B(new_n552), .C1(new_n554), .C2(new_n555), .ZN(G299));
  NAND2_X1  g131(.A1(new_n546), .A2(G89), .ZN(new_n557));
  INV_X1    g132(.A(new_n522), .ZN(new_n558));
  AOI21_X1  g133(.A(KEYINPUT74), .B1(new_n517), .B2(new_n518), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n557), .B(new_n514), .C1(new_n558), .C2(new_n559), .ZN(G286));
  OAI221_X1 g135(.A(new_n504), .B1(new_n509), .B2(new_n510), .C1(new_n497), .C2(new_n498), .ZN(G303));
  OAI21_X1  g136(.A(G651), .B1(new_n496), .B2(G74), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n496), .A2(G87), .A3(new_n501), .A4(new_n503), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n501), .A2(new_n503), .A3(G49), .A4(G543), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(G288));
  NAND3_X1  g140(.A1(new_n546), .A2(KEYINPUT76), .A3(G86), .ZN(new_n566));
  NAND2_X1  g141(.A1(G73), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G61), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n549), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n501), .A2(new_n503), .A3(G543), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G48), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n509), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n566), .A2(new_n570), .A3(new_n573), .A4(new_n576), .ZN(G305));
  NAND4_X1  g152(.A1(new_n496), .A2(G85), .A3(new_n501), .A4(new_n503), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n501), .A2(new_n503), .A3(G47), .A4(G543), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n496), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n498), .ZN(G290));
  NAND2_X1  g156(.A1(G301), .A2(G868), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n506), .A2(new_n508), .A3(G66), .ZN(new_n583));
  NAND2_X1  g158(.A1(G79), .A2(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT78), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n583), .A2(new_n587), .A3(new_n584), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(G651), .A3(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n509), .B2(new_n591), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n501), .A2(new_n503), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n593), .A2(KEYINPUT10), .A3(G92), .A4(new_n496), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(KEYINPUT77), .A3(G543), .ZN(new_n596));
  INV_X1    g171(.A(G54), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n597), .B1(new_n571), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n589), .A2(new_n595), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n582), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n582), .B1(new_n602), .B2(G868), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT9), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n553), .B(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n496), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G91), .ZN(new_n609));
  OAI22_X1  g184(.A1(new_n608), .A2(new_n498), .B1(new_n609), .B2(new_n509), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n605), .B1(G868), .B2(new_n611), .ZN(G297));
  OAI21_X1  g187(.A(new_n605), .B1(G868), .B2(new_n611), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n602), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n602), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n539), .ZN(G323));
  XOR2_X1   g193(.A(KEYINPUT79), .B(KEYINPUT11), .Z(new_n619));
  XNOR2_X1  g194(.A(G323), .B(new_n619), .ZN(G282));
  NAND2_X1  g195(.A1(new_n463), .A2(new_n469), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT13), .Z(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n477), .A2(G123), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n479), .A2(G135), .ZN(new_n626));
  OR2_X1    g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n623), .A2(G2100), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n624), .A2(new_n630), .A3(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2435), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2443), .B(G2446), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT80), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT17), .ZN(new_n651));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n652), .B2(new_n650), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n653), .B1(KEYINPUT81), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(KEYINPUT81), .B2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n651), .A2(new_n654), .A3(new_n652), .ZN(new_n658));
  INV_X1    g233(.A(new_n654), .ZN(new_n659));
  NOR3_X1   g234(.A1(new_n659), .A2(new_n652), .A3(new_n650), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT18), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n657), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n666), .A2(new_n670), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n674));
  OAI221_X1 g249(.A(new_n671), .B1(new_n666), .B2(new_n669), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n674), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT83), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT82), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n680), .B(new_n683), .ZN(G229));
  MUX2_X1   g259(.A(G6), .B(G305), .S(G16), .Z(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT32), .B(G1981), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT85), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G22), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n689), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(G1971), .Z(new_n692));
  NOR2_X1   g267(.A1(G16), .A2(G23), .ZN(new_n693));
  INV_X1    g268(.A(G288), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n693), .B1(new_n694), .B2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT33), .B(G1976), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n688), .A2(new_n692), .A3(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT34), .Z(new_n699));
  AND2_X1   g274(.A1(new_n689), .A2(G24), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G290), .B2(G16), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G1986), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G25), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n479), .A2(G131), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n477), .A2(G119), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT84), .ZN(new_n708));
  OR3_X1    g283(.A1(new_n708), .A2(G95), .A3(G2105), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(G95), .B2(G2105), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n462), .A2(G107), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n709), .A2(new_n710), .A3(G2104), .A4(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n706), .A2(new_n707), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n705), .B1(new_n714), .B2(new_n704), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT35), .B(G1991), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n702), .A2(G1986), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n699), .A2(new_n703), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT36), .Z(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT26), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n477), .A2(G129), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n479), .A2(G141), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI211_X1 g300(.A(new_n722), .B(new_n725), .C1(G105), .C2(new_n469), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G29), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G29), .B2(G32), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT27), .B(G1996), .Z(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n629), .A2(new_n704), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT31), .B(G11), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT90), .ZN(new_n734));
  OR2_X1    g309(.A1(KEYINPUT30), .A2(G28), .ZN(new_n735));
  NAND2_X1  g310(.A1(KEYINPUT30), .A2(G28), .ZN(new_n736));
  AOI21_X1  g311(.A(G29), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR4_X1   g312(.A1(new_n731), .A2(new_n732), .A3(new_n734), .A4(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G16), .A2(G21), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G168), .B2(G16), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G1966), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n539), .A2(new_n689), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n689), .B2(G19), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT86), .B(G1341), .Z(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n738), .A2(new_n741), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n704), .A2(G27), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G164), .B2(new_n704), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2078), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT24), .ZN(new_n751));
  INV_X1    g326(.A(G34), .ZN(new_n752));
  AOI21_X1  g327(.A(G29), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n751), .B2(new_n752), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G160), .B2(new_n704), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n728), .A2(new_n730), .B1(G2084), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G2084), .B2(new_n755), .ZN(new_n757));
  NOR2_X1   g332(.A1(G5), .A2(G16), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G171), .B2(G16), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1961), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n747), .A2(new_n750), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G29), .A2(G35), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G162), .B2(G29), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2090), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n689), .A2(G4), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n602), .B2(new_n689), .ZN(new_n769));
  INV_X1    g344(.A(G1348), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n766), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n740), .A2(G1966), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT91), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n704), .A2(G26), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n477), .A2(G128), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n479), .A2(G140), .ZN(new_n778));
  OR2_X1    g353(.A1(G104), .A2(G2105), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n779), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n776), .B1(new_n782), .B2(new_n704), .ZN(new_n783));
  MUX2_X1   g358(.A(new_n776), .B(new_n783), .S(KEYINPUT28), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2067), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n704), .A2(G33), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n469), .A2(G103), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT88), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n479), .A2(G139), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(KEYINPUT89), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(KEYINPUT89), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n462), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n788), .A2(new_n789), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n792), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n786), .B1(new_n797), .B2(new_n704), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2072), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n689), .A2(G20), .ZN(new_n800));
  OAI211_X1 g375(.A(KEYINPUT23), .B(new_n800), .C1(new_n611), .C2(new_n689), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(KEYINPUT23), .B2(new_n800), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT93), .B(G1956), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n785), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n761), .A2(new_n773), .A3(new_n775), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n720), .A2(new_n806), .ZN(G311));
  INV_X1    g382(.A(G311), .ZN(G150));
  NOR2_X1   g383(.A1(new_n601), .A2(new_n614), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n506), .A2(new_n508), .A3(G56), .ZN(new_n812));
  NAND2_X1  g387(.A1(G68), .A2(G543), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI22_X1  g389(.A1(G43), .A2(new_n572), .B1(new_n814), .B2(G651), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n496), .A2(G93), .A3(new_n501), .A4(new_n503), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n501), .A2(new_n503), .A3(G55), .A4(G543), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n496), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n816), .B(new_n817), .C1(new_n818), .C2(new_n498), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n815), .A2(new_n819), .A3(new_n535), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n506), .A2(new_n508), .A3(G67), .ZN(new_n821));
  NAND2_X1  g396(.A1(G80), .A2(G543), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n498), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n817), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n538), .A2(new_n825), .A3(new_n816), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n820), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(G860), .B1(new_n811), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n828), .B2(new_n811), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n819), .A2(G860), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT37), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(G145));
  NAND2_X1  g408(.A1(new_n492), .A2(new_n494), .ZN(new_n834));
  INV_X1    g409(.A(new_n490), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n781), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n726), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n797), .ZN(new_n839));
  AOI22_X1  g414(.A1(G130), .A2(new_n477), .B1(new_n479), .B2(G142), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT94), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n841), .A2(new_n462), .A3(G118), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n462), .B2(G118), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n843), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n840), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n622), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n714), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n839), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n839), .A2(new_n847), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n629), .B(G160), .ZN(new_n850));
  XNOR2_X1  g425(.A(G162), .B(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n847), .A2(KEYINPUT95), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n851), .B1(new_n839), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n839), .B2(new_n853), .ZN(new_n855));
  INV_X1    g430(.A(G37), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g433(.A(KEYINPUT96), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n601), .B2(new_n611), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n498), .B1(new_n585), .B2(KEYINPUT78), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n861), .A2(new_n588), .B1(new_n596), .B2(new_n599), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n862), .A2(G299), .A3(KEYINPUT96), .A4(new_n595), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT97), .B1(new_n601), .B2(new_n611), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n601), .A2(KEYINPUT97), .A3(new_n611), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n864), .A2(new_n866), .A3(KEYINPUT41), .A4(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n601), .A2(KEYINPUT97), .A3(new_n611), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(new_n865), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT41), .B1(new_n871), .B2(new_n864), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n616), .B(new_n828), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n871), .A2(KEYINPUT98), .A3(new_n864), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT98), .B1(new_n871), .B2(new_n864), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI22_X1  g453(.A1(new_n875), .A2(KEYINPUT99), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n873), .A2(new_n874), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n694), .A2(G290), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n506), .A2(new_n508), .A3(G60), .ZN(new_n884));
  NAND2_X1  g459(.A1(G72), .A2(G543), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n498), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n579), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(G288), .B1(new_n888), .B2(new_n578), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT100), .B1(new_n883), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(G305), .A2(G166), .ZN(new_n891));
  AOI22_X1  g466(.A1(G651), .A2(new_n569), .B1(new_n572), .B2(G48), .ZN(new_n892));
  NAND4_X1  g467(.A1(G303), .A2(new_n566), .A3(new_n892), .A4(new_n576), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n694), .A2(G290), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n888), .A2(G288), .A3(new_n578), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n890), .A2(new_n891), .A3(new_n893), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n893), .A2(new_n891), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(KEYINPUT42), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n898), .A2(new_n905), .A3(new_n901), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n905), .B1(new_n898), .B2(new_n901), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n904), .B1(KEYINPUT42), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n879), .A2(new_n882), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n882), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n878), .A2(new_n874), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(new_n880), .B2(new_n881), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n909), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT103), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n879), .A2(KEYINPUT102), .A3(new_n882), .A4(new_n910), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n920), .B(new_n909), .C1(new_n914), .C2(new_n916), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n913), .A2(new_n918), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  MUX2_X1   g497(.A(new_n819), .B(new_n922), .S(G868), .Z(G295));
  MUX2_X1   g498(.A(new_n819), .B(new_n922), .S(G868), .Z(G331));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n926), .B1(new_n820), .B2(new_n826), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n526), .B(new_n929), .C1(new_n530), .C2(new_n532), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(G168), .ZN(new_n931));
  INV_X1    g506(.A(new_n530), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(G651), .A3(new_n531), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n929), .B1(new_n933), .B2(new_n526), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(G301), .A2(KEYINPUT104), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(G168), .A3(new_n930), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n820), .A2(new_n826), .A3(new_n926), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n928), .A2(new_n935), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n931), .A2(new_n934), .ZN(new_n940));
  AND3_X1   g515(.A1(G286), .A2(KEYINPUT104), .A3(G301), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n820), .A2(new_n826), .A3(new_n926), .ZN(new_n942));
  OAI22_X1  g517(.A1(new_n940), .A2(new_n941), .B1(new_n942), .B2(new_n927), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n939), .B(new_n943), .C1(new_n876), .C2(new_n877), .ZN(new_n944));
  OR2_X1    g519(.A1(new_n906), .A2(new_n907), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n868), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n864), .A2(new_n866), .A3(new_n867), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT41), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n943), .A2(new_n939), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n871), .A2(KEYINPUT107), .A3(KEYINPUT41), .A4(new_n864), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n947), .A2(new_n950), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n944), .A2(new_n945), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n951), .B1(new_n869), .B2(new_n872), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n948), .A2(new_n943), .A3(new_n939), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n908), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n957), .A3(new_n856), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n925), .B1(new_n958), .B2(KEYINPUT43), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n908), .B1(new_n955), .B2(new_n956), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n960), .B1(new_n961), .B2(G37), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n948), .A2(new_n943), .A3(new_n939), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n950), .A2(new_n868), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n951), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT106), .B(new_n856), .C1(new_n965), .C2(new_n908), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n966), .A3(new_n957), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n959), .B1(new_n967), .B2(KEYINPUT43), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n970));
  AND4_X1   g545(.A1(new_n970), .A2(new_n954), .A3(new_n957), .A4(new_n856), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT108), .B1(new_n973), .B2(new_n925), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n971), .B1(new_n967), .B2(KEYINPUT43), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT44), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n968), .B1(new_n974), .B2(new_n977), .ZN(G397));
  INV_X1    g553(.A(G2067), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n781), .B(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT110), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n726), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(G164), .B2(G1384), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G40), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n466), .A2(new_n471), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n988), .A2(G1996), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(KEYINPUT46), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n992), .B1(KEYINPUT46), .B2(new_n991), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n991), .A2(new_n726), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n997), .A2(KEYINPUT109), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(KEYINPUT109), .ZN(new_n999));
  INV_X1    g574(.A(G1996), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n981), .A2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n998), .B(new_n999), .C1(new_n990), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n714), .A2(new_n716), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n714), .A2(new_n716), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n988), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n988), .A2(G1986), .A3(G290), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT48), .ZN(new_n1008));
  OAI22_X1  g583(.A1(new_n995), .A2(new_n996), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  OAI22_X1  g584(.A1(new_n1002), .A2(new_n1003), .B1(G2067), .B2(new_n781), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n989), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT127), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1011), .A2(KEYINPUT127), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1009), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1384), .B1(new_n834), .B2(new_n835), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n987), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G8), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT114), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n694), .A2(G1976), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1017), .A2(KEYINPUT114), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(new_n1016), .B2(G8), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1019), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n892), .B1(new_n575), .B2(new_n509), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(G1981), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n892), .A2(new_n1030), .A3(new_n566), .A4(new_n576), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT49), .B1(new_n1032), .B2(KEYINPUT115), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT49), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n1034), .B(new_n1035), .C1(new_n1029), .C2(new_n1031), .ZN(new_n1036));
  OAI22_X1  g611(.A1(new_n1033), .A2(new_n1036), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1022), .A2(new_n1027), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G8), .ZN(new_n1039));
  INV_X1    g614(.A(G1384), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n836), .A2(KEYINPUT45), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n984), .A2(new_n1041), .A3(new_n987), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT111), .B(G1971), .Z(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n836), .A2(new_n1046), .A3(new_n1040), .ZN(new_n1047));
  INV_X1    g622(.A(G2090), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .A4(new_n987), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1039), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G303), .A2(G8), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  NAND4_X1  g630(.A1(G303), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1050), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT113), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1050), .A2(new_n1060), .A3(new_n1057), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1045), .A2(new_n987), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT116), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1045), .A2(new_n1065), .A3(new_n987), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1064), .A2(new_n1047), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1044), .B1(new_n1067), .B2(G2090), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G8), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1057), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1038), .A2(new_n1062), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  OR3_X1    g648(.A1(new_n1042), .A2(new_n1073), .A3(G2078), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1073), .B1(new_n1042), .B2(G2078), .ZN(new_n1075));
  INV_X1    g650(.A(G1961), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1047), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1076), .B1(new_n1063), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1074), .A2(new_n1075), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(G171), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1072), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(G168), .A2(new_n1039), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1045), .A2(new_n1047), .A3(new_n987), .ZN(new_n1084));
  INV_X1    g659(.A(G2084), .ZN(new_n1085));
  INV_X1    g660(.A(G1966), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1084), .A2(new_n1085), .B1(new_n1042), .B2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(KEYINPUT51), .B(new_n1083), .C1(new_n1087), .C2(new_n1039), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1042), .A2(new_n1086), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1045), .A2(new_n1047), .A3(new_n1085), .A4(new_n987), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1089), .B(G8), .C1(new_n1092), .C2(G286), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT122), .B1(new_n1092), .B2(new_n1082), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n1095));
  AOI211_X1 g670(.A(new_n1095), .B(new_n1083), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1088), .B(new_n1093), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT123), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1095), .B1(new_n1087), .B2(new_n1083), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1092), .A2(KEYINPUT122), .A3(new_n1082), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1101), .A2(new_n1102), .A3(new_n1088), .A4(new_n1093), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1098), .A2(KEYINPUT62), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT62), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1081), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1022), .A2(new_n1027), .A3(new_n1037), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT63), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1087), .A2(new_n1039), .A3(G286), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1071), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1107), .B1(new_n1110), .B2(new_n1062), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1109), .B1(new_n1057), .B2(new_n1050), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT63), .B1(new_n1112), .B2(new_n1107), .ZN(new_n1113));
  NOR4_X1   g688(.A1(new_n1033), .A2(new_n1036), .A3(G1976), .A4(G288), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1031), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1018), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1111), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1106), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n464), .A2(new_n465), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT124), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1121), .A2(KEYINPUT124), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(G2105), .A3(new_n1123), .ZN(new_n1124));
  NOR4_X1   g699(.A1(new_n471), .A2(new_n1073), .A3(new_n986), .A4(G2078), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n984), .A3(new_n1041), .A4(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1075), .A2(new_n1078), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1120), .B1(new_n1127), .B2(G171), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1079), .B2(G171), .ZN(new_n1129));
  AND4_X1   g704(.A1(new_n1071), .A2(new_n1038), .A3(new_n1129), .A4(new_n1062), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT125), .B1(new_n1127), .B2(G171), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1080), .A2(new_n1131), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1127), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1120), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1130), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(G2072), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1042), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(G1956), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n1067), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT57), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n607), .B2(KEYINPUT117), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(G299), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT119), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1077), .B1(new_n1063), .B2(KEYINPUT116), .ZN(new_n1151));
  AOI21_X1  g726(.A(G1956), .B1(new_n1151), .B2(new_n1066), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1146), .B1(new_n1152), .B2(new_n1141), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1143), .A2(KEYINPUT119), .A3(new_n1147), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1150), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1016), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n987), .A2(new_n1015), .A3(KEYINPUT120), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n979), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n770), .B1(new_n1063), .B2(new_n1077), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n602), .ZN(new_n1165));
  NOR2_X1   g740(.A1(KEYINPUT121), .A2(G1996), .ZN(new_n1166));
  AND2_X1   g741(.A1(KEYINPUT121), .A2(G1996), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1042), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(KEYINPUT58), .B(G1341), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1169), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n539), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT59), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1173), .B(new_n539), .C1(new_n1168), .C2(new_n1170), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1165), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1148), .A2(KEYINPUT61), .A3(new_n1153), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n601), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1177), .B1(new_n1164), .B2(new_n1163), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1157), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1163), .A2(new_n602), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1153), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1150), .A2(new_n1182), .A3(new_n1154), .ZN(new_n1183));
  AOI22_X1  g758(.A1(new_n1136), .A2(new_n1137), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1119), .B1(new_n1138), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1006), .ZN(new_n1186));
  XOR2_X1   g761(.A(G290), .B(G1986), .Z(new_n1187));
  OAI21_X1  g762(.A(new_n1186), .B1(new_n988), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1014), .B1(new_n1185), .B2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g764(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1191));
  AND3_X1   g765(.A1(new_n1191), .A2(new_n857), .A3(new_n973), .ZN(G308));
  NAND3_X1  g766(.A1(new_n1191), .A2(new_n857), .A3(new_n973), .ZN(G225));
endmodule


