

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594;

  XNOR2_X1 U326 ( .A(n308), .B(n307), .ZN(n309) );
  INV_X1 U327 ( .A(KEYINPUT10), .ZN(n307) );
  AND2_X1 U328 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U329 ( .A(n493), .B(KEYINPUT99), .Z(n295) );
  NOR2_X1 U330 ( .A1(n480), .A2(n465), .ZN(n466) );
  INV_X1 U331 ( .A(KEYINPUT94), .ZN(n467) );
  XNOR2_X1 U332 ( .A(n398), .B(n294), .ZN(n302) );
  XOR2_X1 U333 ( .A(G197GAT), .B(KEYINPUT21), .Z(n415) );
  XNOR2_X1 U334 ( .A(n302), .B(n378), .ZN(n303) );
  XNOR2_X1 U335 ( .A(KEYINPUT116), .B(KEYINPUT47), .ZN(n368) );
  INV_X1 U336 ( .A(n380), .ZN(n381) );
  XNOR2_X1 U337 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U338 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n435) );
  XNOR2_X1 U339 ( .A(n369), .B(n368), .ZN(n375) );
  XNOR2_X1 U340 ( .A(n382), .B(n381), .ZN(n386) );
  XNOR2_X1 U341 ( .A(n332), .B(n331), .ZN(n336) );
  INV_X1 U342 ( .A(KEYINPUT96), .ZN(n488) );
  XNOR2_X1 U343 ( .A(n386), .B(n385), .ZN(n392) );
  XNOR2_X1 U344 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U345 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U346 ( .A(KEYINPUT97), .B(n491), .Z(n500) );
  XNOR2_X1 U347 ( .A(n342), .B(n341), .ZN(n584) );
  XNOR2_X1 U348 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U349 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XOR2_X1 U350 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n297) );
  XNOR2_X1 U351 ( .A(G92GAT), .B(KEYINPUT77), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n312) );
  XOR2_X1 U353 ( .A(KEYINPUT76), .B(KEYINPUT66), .Z(n299) );
  XOR2_X1 U354 ( .A(G99GAT), .B(G85GAT), .Z(n327) );
  XOR2_X1 U355 ( .A(G50GAT), .B(KEYINPUT75), .Z(n420) );
  XNOR2_X1 U356 ( .A(n327), .B(n420), .ZN(n298) );
  XNOR2_X1 U357 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U358 ( .A(n300), .B(G106GAT), .Z(n305) );
  XOR2_X1 U359 ( .A(G29GAT), .B(G134GAT), .Z(n398) );
  XNOR2_X1 U360 ( .A(G36GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n301), .B(G218GAT), .ZN(n378) );
  XNOR2_X1 U362 ( .A(G162GAT), .B(n303), .ZN(n304) );
  XNOR2_X1 U363 ( .A(n305), .B(n304), .ZN(n310) );
  XNOR2_X1 U364 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n306) );
  XNOR2_X1 U365 ( .A(n306), .B(KEYINPUT7), .ZN(n351) );
  XNOR2_X1 U366 ( .A(n351), .B(KEYINPUT78), .ZN(n308) );
  XNOR2_X1 U367 ( .A(n312), .B(n311), .ZN(n570) );
  XOR2_X1 U368 ( .A(G22GAT), .B(G15GAT), .Z(n348) );
  XNOR2_X1 U369 ( .A(n348), .B(G64GAT), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n313), .B(KEYINPUT79), .ZN(n326) );
  XNOR2_X1 U371 ( .A(G8GAT), .B(G183GAT), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n314), .B(G211GAT), .ZN(n379) );
  XOR2_X1 U373 ( .A(KEYINPUT14), .B(n379), .Z(n316) );
  NAND2_X1 U374 ( .A1(G231GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U376 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n318) );
  XNOR2_X1 U377 ( .A(G78GAT), .B(KEYINPUT15), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U379 ( .A(n320), .B(n319), .Z(n324) );
  XNOR2_X1 U380 ( .A(G1GAT), .B(G127GAT), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n321), .B(G155GAT), .ZN(n397) );
  XNOR2_X1 U382 ( .A(G71GAT), .B(G57GAT), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n322), .B(KEYINPUT13), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n397), .B(n328), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U386 ( .A(n326), .B(n325), .Z(n485) );
  XOR2_X1 U387 ( .A(KEYINPUT114), .B(n485), .Z(n574) );
  XOR2_X1 U388 ( .A(n328), .B(n327), .Z(n332) );
  NAND2_X1 U389 ( .A1(G230GAT), .A2(G233GAT), .ZN(n330) );
  INV_X1 U390 ( .A(KEYINPUT32), .ZN(n329) );
  XOR2_X1 U391 ( .A(G64GAT), .B(G204GAT), .Z(n334) );
  XNOR2_X1 U392 ( .A(G176GAT), .B(G92GAT), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n380) );
  XNOR2_X1 U394 ( .A(n380), .B(KEYINPUT31), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n342) );
  XOR2_X1 U396 ( .A(G120GAT), .B(G148GAT), .Z(n399) );
  XOR2_X1 U397 ( .A(G106GAT), .B(G78GAT), .Z(n416) );
  XNOR2_X1 U398 ( .A(n399), .B(n416), .ZN(n340) );
  XOR2_X1 U399 ( .A(KEYINPUT74), .B(KEYINPUT72), .Z(n338) );
  XNOR2_X1 U400 ( .A(KEYINPUT33), .B(KEYINPUT73), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n584), .B(KEYINPUT64), .ZN(n344) );
  INV_X1 U403 ( .A(KEYINPUT41), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n460) );
  XOR2_X1 U405 ( .A(G8GAT), .B(G197GAT), .Z(n346) );
  XNOR2_X1 U406 ( .A(G29GAT), .B(G50GAT), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U408 ( .A(n347), .B(G36GAT), .Z(n350) );
  XNOR2_X1 U409 ( .A(G169GAT), .B(n348), .ZN(n349) );
  XNOR2_X1 U410 ( .A(n350), .B(n349), .ZN(n355) );
  XOR2_X1 U411 ( .A(n351), .B(KEYINPUT70), .Z(n353) );
  NAND2_X1 U412 ( .A1(G229GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U414 ( .A(n355), .B(n354), .Z(n363) );
  XOR2_X1 U415 ( .A(KEYINPUT71), .B(KEYINPUT68), .Z(n357) );
  XNOR2_X1 U416 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U418 ( .A(G141GAT), .B(G113GAT), .Z(n359) );
  XNOR2_X1 U419 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U422 ( .A(n363), .B(n362), .Z(n548) );
  INV_X1 U423 ( .A(n548), .ZN(n580) );
  NAND2_X1 U424 ( .A1(n460), .A2(n580), .ZN(n364) );
  XOR2_X1 U425 ( .A(n364), .B(KEYINPUT46), .Z(n365) );
  NOR2_X1 U426 ( .A1(n574), .A2(n365), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n366), .B(KEYINPUT115), .ZN(n367) );
  NOR2_X1 U428 ( .A1(n570), .A2(n367), .ZN(n369) );
  INV_X1 U429 ( .A(n584), .ZN(n490) );
  XNOR2_X1 U430 ( .A(KEYINPUT36), .B(n570), .ZN(n589) );
  INV_X1 U431 ( .A(n485), .ZN(n587) );
  NAND2_X1 U432 ( .A1(n589), .A2(n587), .ZN(n371) );
  XOR2_X1 U433 ( .A(KEYINPUT45), .B(KEYINPUT117), .Z(n370) );
  XNOR2_X1 U434 ( .A(n371), .B(n370), .ZN(n372) );
  NOR2_X1 U435 ( .A1(n580), .A2(n372), .ZN(n373) );
  NAND2_X1 U436 ( .A1(n490), .A2(n373), .ZN(n374) );
  NAND2_X1 U437 ( .A1(n375), .A2(n374), .ZN(n377) );
  INV_X1 U438 ( .A(KEYINPUT48), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n562) );
  XNOR2_X1 U440 ( .A(n379), .B(n378), .ZN(n382) );
  XOR2_X1 U441 ( .A(KEYINPUT90), .B(n415), .Z(n384) );
  NAND2_X1 U442 ( .A1(G226GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U444 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n387), .B(KEYINPUT17), .ZN(n388) );
  XOR2_X1 U446 ( .A(n388), .B(KEYINPUT82), .Z(n390) );
  XNOR2_X1 U447 ( .A(G169GAT), .B(KEYINPUT83), .ZN(n389) );
  XOR2_X1 U448 ( .A(n390), .B(n389), .Z(n450) );
  INV_X1 U449 ( .A(n450), .ZN(n391) );
  XOR2_X1 U450 ( .A(n392), .B(n391), .Z(n469) );
  NOR2_X1 U451 ( .A1(n562), .A2(n469), .ZN(n394) );
  INV_X1 U452 ( .A(KEYINPUT54), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n413) );
  XOR2_X1 U454 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n396) );
  XNOR2_X1 U455 ( .A(G141GAT), .B(G162GAT), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n419) );
  XNOR2_X1 U457 ( .A(n397), .B(n419), .ZN(n412) );
  XOR2_X1 U458 ( .A(n399), .B(n398), .Z(n401) );
  NAND2_X1 U459 ( .A1(G225GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U461 ( .A(KEYINPUT6), .B(KEYINPUT87), .Z(n403) );
  XNOR2_X1 U462 ( .A(KEYINPUT88), .B(KEYINPUT1), .ZN(n402) );
  XNOR2_X1 U463 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U464 ( .A(n405), .B(n404), .Z(n410) );
  XOR2_X1 U465 ( .A(G113GAT), .B(KEYINPUT0), .Z(n440) );
  XOR2_X1 U466 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n407) );
  XNOR2_X1 U467 ( .A(G85GAT), .B(G57GAT), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n440), .B(n408), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n475) );
  XNOR2_X1 U472 ( .A(KEYINPUT89), .B(n475), .ZN(n534) );
  NOR2_X1 U473 ( .A1(n413), .A2(n534), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n414), .B(KEYINPUT65), .ZN(n577) );
  XOR2_X1 U475 ( .A(n416), .B(n415), .Z(n418) );
  XNOR2_X1 U476 ( .A(G218GAT), .B(G204GAT), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n424) );
  XOR2_X1 U478 ( .A(n420), .B(n419), .Z(n422) );
  NAND2_X1 U479 ( .A1(G228GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U481 ( .A(n424), .B(n423), .Z(n426) );
  XNOR2_X1 U482 ( .A(G22GAT), .B(G211GAT), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n434) );
  XOR2_X1 U484 ( .A(KEYINPUT86), .B(KEYINPUT23), .Z(n428) );
  XNOR2_X1 U485 ( .A(G155GAT), .B(G148GAT), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U487 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n430) );
  XNOR2_X1 U488 ( .A(KEYINPUT84), .B(KEYINPUT24), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U490 ( .A(n432), .B(n431), .Z(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n480) );
  NOR2_X1 U492 ( .A1(n577), .A2(n480), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n453) );
  XOR2_X1 U494 ( .A(G190GAT), .B(G99GAT), .Z(n438) );
  XNOR2_X1 U495 ( .A(G43GAT), .B(G134GAT), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U497 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U500 ( .A(KEYINPUT81), .B(KEYINPUT20), .Z(n444) );
  XNOR2_X1 U501 ( .A(G127GAT), .B(G120GAT), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U503 ( .A(n446), .B(n445), .Z(n452) );
  XOR2_X1 U504 ( .A(G71GAT), .B(G183GAT), .Z(n448) );
  XNOR2_X1 U505 ( .A(G15GAT), .B(G176GAT), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U507 ( .A(n450), .B(n449), .Z(n451) );
  XOR2_X1 U508 ( .A(n452), .B(n451), .Z(n470) );
  INV_X1 U509 ( .A(n470), .ZN(n547) );
  NAND2_X1 U510 ( .A1(n453), .A2(n547), .ZN(n455) );
  INV_X1 U511 ( .A(KEYINPUT122), .ZN(n454) );
  XNOR2_X2 U512 ( .A(n455), .B(n454), .ZN(n575) );
  NAND2_X1 U513 ( .A1(n575), .A2(n570), .ZN(n459) );
  XOR2_X1 U514 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n457) );
  XNOR2_X1 U515 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n456) );
  NAND2_X1 U516 ( .A1(n575), .A2(n460), .ZN(n463) );
  XOR2_X1 U517 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n461) );
  XNOR2_X1 U518 ( .A(n461), .B(G176GAT), .ZN(n462) );
  XNOR2_X1 U519 ( .A(n463), .B(n462), .ZN(G1349GAT) );
  NOR2_X1 U520 ( .A1(n469), .A2(n470), .ZN(n464) );
  XOR2_X1 U521 ( .A(KEYINPUT93), .B(n464), .Z(n465) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n466), .Z(n468) );
  XNOR2_X1 U523 ( .A(n468), .B(n467), .ZN(n474) );
  INV_X1 U524 ( .A(n469), .ZN(n537) );
  XNOR2_X1 U525 ( .A(n537), .B(KEYINPUT27), .ZN(n478) );
  NAND2_X1 U526 ( .A1(n480), .A2(n470), .ZN(n471) );
  XNOR2_X1 U527 ( .A(n471), .B(KEYINPUT26), .ZN(n472) );
  XOR2_X1 U528 ( .A(KEYINPUT92), .B(n472), .Z(n578) );
  NAND2_X1 U529 ( .A1(n478), .A2(n578), .ZN(n473) );
  NAND2_X1 U530 ( .A1(n474), .A2(n473), .ZN(n476) );
  NAND2_X1 U531 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U532 ( .A(n477), .B(KEYINPUT95), .ZN(n484) );
  NAND2_X1 U533 ( .A1(n534), .A2(n478), .ZN(n479) );
  XNOR2_X1 U534 ( .A(n479), .B(KEYINPUT91), .ZN(n560) );
  XNOR2_X1 U535 ( .A(KEYINPUT67), .B(KEYINPUT28), .ZN(n481) );
  XOR2_X1 U536 ( .A(n481), .B(n480), .Z(n541) );
  INV_X1 U537 ( .A(n541), .ZN(n482) );
  NAND2_X1 U538 ( .A1(n560), .A2(n482), .ZN(n545) );
  NOR2_X1 U539 ( .A1(n545), .A2(n547), .ZN(n483) );
  NOR2_X1 U540 ( .A1(n484), .A2(n483), .ZN(n503) );
  NOR2_X1 U541 ( .A1(n485), .A2(n570), .ZN(n486) );
  XOR2_X1 U542 ( .A(KEYINPUT16), .B(n486), .Z(n487) );
  NOR2_X1 U543 ( .A1(n503), .A2(n487), .ZN(n489) );
  XNOR2_X1 U544 ( .A(n489), .B(n488), .ZN(n518) );
  NAND2_X1 U545 ( .A1(n580), .A2(n490), .ZN(n507) );
  NOR2_X1 U546 ( .A1(n518), .A2(n507), .ZN(n491) );
  NAND2_X1 U547 ( .A1(n534), .A2(n500), .ZN(n492) );
  XNOR2_X1 U548 ( .A(n492), .B(KEYINPUT34), .ZN(n493) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n494) );
  XNOR2_X1 U550 ( .A(n295), .B(n494), .ZN(G1324GAT) );
  NAND2_X1 U551 ( .A1(n537), .A2(n500), .ZN(n495) );
  XNOR2_X1 U552 ( .A(n495), .B(KEYINPUT100), .ZN(n496) );
  XNOR2_X1 U553 ( .A(G8GAT), .B(n496), .ZN(G1325GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n498) );
  NAND2_X1 U555 ( .A1(n500), .A2(n547), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U557 ( .A(G15GAT), .B(n499), .Z(G1326GAT) );
  NAND2_X1 U558 ( .A1(n500), .A2(n541), .ZN(n501) );
  XNOR2_X1 U559 ( .A(n501), .B(KEYINPUT102), .ZN(n502) );
  XNOR2_X1 U560 ( .A(G22GAT), .B(n502), .ZN(G1327GAT) );
  NOR2_X1 U561 ( .A1(n503), .A2(n587), .ZN(n504) );
  XOR2_X1 U562 ( .A(KEYINPUT103), .B(n504), .Z(n505) );
  NAND2_X1 U563 ( .A1(n589), .A2(n505), .ZN(n506) );
  XOR2_X1 U564 ( .A(KEYINPUT37), .B(n506), .Z(n533) );
  NOR2_X1 U565 ( .A1(n533), .A2(n507), .ZN(n509) );
  XNOR2_X1 U566 ( .A(KEYINPUT38), .B(KEYINPUT104), .ZN(n508) );
  XNOR2_X1 U567 ( .A(n509), .B(n508), .ZN(n515) );
  NAND2_X1 U568 ( .A1(n515), .A2(n534), .ZN(n511) );
  XOR2_X1 U569 ( .A(G29GAT), .B(KEYINPUT39), .Z(n510) );
  XNOR2_X1 U570 ( .A(n511), .B(n510), .ZN(G1328GAT) );
  NAND2_X1 U571 ( .A1(n515), .A2(n537), .ZN(n512) );
  XNOR2_X1 U572 ( .A(G36GAT), .B(n512), .ZN(G1329GAT) );
  NAND2_X1 U573 ( .A1(n515), .A2(n547), .ZN(n513) );
  XNOR2_X1 U574 ( .A(n513), .B(KEYINPUT40), .ZN(n514) );
  XNOR2_X1 U575 ( .A(G43GAT), .B(n514), .ZN(G1330GAT) );
  XOR2_X1 U576 ( .A(G50GAT), .B(KEYINPUT105), .Z(n517) );
  NAND2_X1 U577 ( .A1(n515), .A2(n541), .ZN(n516) );
  XNOR2_X1 U578 ( .A(n517), .B(n516), .ZN(G1331GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n520) );
  NAND2_X1 U580 ( .A1(n460), .A2(n548), .ZN(n532) );
  NOR2_X1 U581 ( .A1(n518), .A2(n532), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n527), .A2(n534), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U584 ( .A(G57GAT), .B(n521), .Z(G1332GAT) );
  XOR2_X1 U585 ( .A(G64GAT), .B(KEYINPUT107), .Z(n523) );
  NAND2_X1 U586 ( .A1(n527), .A2(n537), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(G1333GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n525) );
  NAND2_X1 U589 ( .A1(n527), .A2(n547), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G71GAT), .B(n526), .ZN(G1334GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n529) );
  NAND2_X1 U593 ( .A1(n527), .A2(n541), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(n531) );
  XOR2_X1 U595 ( .A(G78GAT), .B(KEYINPUT111), .Z(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(G1335GAT) );
  XNOR2_X1 U597 ( .A(G85GAT), .B(KEYINPUT112), .ZN(n536) );
  NOR2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n542), .A2(n534), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1336GAT) );
  NAND2_X1 U601 ( .A1(n537), .A2(n542), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n538), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U603 ( .A(G99GAT), .B(KEYINPUT113), .Z(n540) );
  NAND2_X1 U604 ( .A1(n542), .A2(n547), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1338GAT) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n543), .B(KEYINPUT44), .ZN(n544) );
  XNOR2_X1 U608 ( .A(G106GAT), .B(n544), .ZN(G1339GAT) );
  NOR2_X1 U609 ( .A1(n562), .A2(n545), .ZN(n546) );
  NAND2_X1 U610 ( .A1(n547), .A2(n546), .ZN(n550) );
  NOR2_X1 U611 ( .A1(n548), .A2(n550), .ZN(n549) );
  XOR2_X1 U612 ( .A(G113GAT), .B(n549), .Z(G1340GAT) );
  INV_X1 U613 ( .A(n550), .ZN(n556) );
  AND2_X1 U614 ( .A1(n460), .A2(n556), .ZN(n552) );
  XNOR2_X1 U615 ( .A(KEYINPUT118), .B(KEYINPUT49), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U617 ( .A(G120GAT), .B(n553), .ZN(G1341GAT) );
  NAND2_X1 U618 ( .A1(n556), .A2(n574), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(KEYINPUT50), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G127GAT), .B(n555), .ZN(G1342GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n558) );
  NAND2_X1 U622 ( .A1(n556), .A2(n570), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U624 ( .A(G134GAT), .B(n559), .Z(G1343GAT) );
  NAND2_X1 U625 ( .A1(n578), .A2(n560), .ZN(n561) );
  NOR2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n569) );
  NAND2_X1 U627 ( .A1(n569), .A2(n580), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n565) );
  NAND2_X1 U630 ( .A1(n569), .A2(n460), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G148GAT), .B(n566), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n587), .A2(n569), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT120), .ZN(n568) );
  XNOR2_X1 U635 ( .A(G155GAT), .B(n568), .ZN(G1346GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U638 ( .A(G169GAT), .B(KEYINPUT123), .Z(n573) );
  NAND2_X1 U639 ( .A1(n580), .A2(n575), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(G1348GAT) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n576), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n582) );
  INV_X1 U644 ( .A(n578), .ZN(n579) );
  NOR2_X1 U645 ( .A1(n577), .A2(n579), .ZN(n590) );
  NAND2_X1 U646 ( .A1(n590), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U650 ( .A1(n590), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n590), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n594) );
  XOR2_X1 U655 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n592) );
  NAND2_X1 U656 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n594), .B(n593), .ZN(G1355GAT) );
endmodule

