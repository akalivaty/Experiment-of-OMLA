

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U548 ( .A1(n680), .A2(n770), .ZN(n732) );
  XNOR2_X1 U549 ( .A(KEYINPUT17), .B(KEYINPUT69), .ZN(n514) );
  NOR2_X1 U550 ( .A1(G2105), .A2(G2104), .ZN(n513) );
  XNOR2_X1 U551 ( .A(n514), .B(n513), .ZN(n874) );
  NAND2_X1 U552 ( .A1(G137), .A2(n874), .ZN(n516) );
  AND2_X1 U553 ( .A1(G2105), .A2(G2104), .ZN(n868) );
  NAND2_X1 U554 ( .A1(G113), .A2(n868), .ZN(n515) );
  AND2_X1 U555 ( .A1(n516), .A2(n515), .ZN(n673) );
  INV_X1 U556 ( .A(KEYINPUT23), .ZN(n519) );
  INV_X1 U557 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U558 ( .A1(n521), .A2(G2104), .ZN(n517) );
  XNOR2_X2 U559 ( .A(n517), .B(KEYINPUT67), .ZN(n872) );
  NAND2_X1 U560 ( .A1(G101), .A2(n872), .ZN(n518) );
  XNOR2_X1 U561 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U562 ( .A(n520), .B(KEYINPUT68), .ZN(n524) );
  NOR2_X1 U563 ( .A1(n521), .A2(G2104), .ZN(n522) );
  XNOR2_X1 U564 ( .A(n522), .B(KEYINPUT66), .ZN(n869) );
  NAND2_X1 U565 ( .A1(G125), .A2(n869), .ZN(n523) );
  AND2_X1 U566 ( .A1(n524), .A2(n523), .ZN(n675) );
  AND2_X1 U567 ( .A1(n673), .A2(n675), .ZN(G160) );
  AND2_X1 U568 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U569 ( .A(G132), .ZN(G219) );
  INV_X1 U570 ( .A(G82), .ZN(G220) );
  INV_X1 U571 ( .A(G651), .ZN(n530) );
  NOR2_X1 U572 ( .A1(G543), .A2(n530), .ZN(n525) );
  XOR2_X1 U573 ( .A(KEYINPUT1), .B(n525), .Z(n629) );
  NAND2_X1 U574 ( .A1(G64), .A2(n629), .ZN(n528) );
  XOR2_X1 U575 ( .A(G543), .B(KEYINPUT0), .Z(n623) );
  NOR2_X1 U576 ( .A1(G651), .A2(n623), .ZN(n526) );
  XOR2_X1 U577 ( .A(KEYINPUT65), .B(n526), .Z(n628) );
  NAND2_X1 U578 ( .A1(G52), .A2(n628), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U580 ( .A(KEYINPUT71), .B(n529), .Z(n536) );
  NOR2_X1 U581 ( .A1(n623), .A2(n530), .ZN(n634) );
  NAND2_X1 U582 ( .A1(n634), .A2(G77), .ZN(n533) );
  NOR2_X1 U583 ( .A1(G543), .A2(G651), .ZN(n531) );
  XNOR2_X1 U584 ( .A(n531), .B(KEYINPUT64), .ZN(n633) );
  NAND2_X1 U585 ( .A1(G90), .A2(n633), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U587 ( .A(KEYINPUT9), .B(n534), .Z(n535) );
  NOR2_X1 U588 ( .A1(n536), .A2(n535), .ZN(G171) );
  XOR2_X1 U589 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n538) );
  NAND2_X1 U590 ( .A1(G7), .A2(G661), .ZN(n537) );
  XNOR2_X1 U591 ( .A(n538), .B(n537), .ZN(G223) );
  XOR2_X1 U592 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n540) );
  INV_X1 U593 ( .A(G223), .ZN(n816) );
  NAND2_X1 U594 ( .A1(G567), .A2(n816), .ZN(n539) );
  XNOR2_X1 U595 ( .A(n540), .B(n539), .ZN(G234) );
  NAND2_X1 U596 ( .A1(G56), .A2(n629), .ZN(n541) );
  XOR2_X1 U597 ( .A(KEYINPUT14), .B(n541), .Z(n548) );
  NAND2_X1 U598 ( .A1(n633), .A2(G81), .ZN(n542) );
  XOR2_X1 U599 ( .A(KEYINPUT12), .B(n542), .Z(n543) );
  XNOR2_X1 U600 ( .A(n543), .B(KEYINPUT75), .ZN(n545) );
  NAND2_X1 U601 ( .A1(G68), .A2(n634), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U603 ( .A(KEYINPUT13), .B(n546), .Z(n547) );
  NOR2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n628), .A2(G43), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n940) );
  INV_X1 U607 ( .A(G860), .ZN(n582) );
  OR2_X1 U608 ( .A1(n940), .A2(n582), .ZN(G153) );
  INV_X1 U609 ( .A(G171), .ZN(G301) );
  NAND2_X1 U610 ( .A1(G66), .A2(n629), .ZN(n552) );
  NAND2_X1 U611 ( .A1(G92), .A2(n633), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U613 ( .A1(G54), .A2(n628), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G79), .A2(n634), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U616 ( .A1(n556), .A2(n555), .ZN(n558) );
  XNOR2_X1 U617 ( .A(KEYINPUT76), .B(KEYINPUT15), .ZN(n557) );
  XNOR2_X1 U618 ( .A(n558), .B(n557), .ZN(n888) );
  NOR2_X1 U619 ( .A1(n888), .A2(G868), .ZN(n560) );
  INV_X1 U620 ( .A(G868), .ZN(n649) );
  NOR2_X1 U621 ( .A1(n649), .A2(G301), .ZN(n559) );
  NOR2_X1 U622 ( .A1(n560), .A2(n559), .ZN(G284) );
  NAND2_X1 U623 ( .A1(G89), .A2(n633), .ZN(n561) );
  XNOR2_X1 U624 ( .A(n561), .B(KEYINPUT4), .ZN(n563) );
  NAND2_X1 U625 ( .A1(G76), .A2(n634), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U627 ( .A(n564), .B(KEYINPUT5), .ZN(n570) );
  XNOR2_X1 U628 ( .A(KEYINPUT77), .B(KEYINPUT6), .ZN(n568) );
  NAND2_X1 U629 ( .A1(G63), .A2(n629), .ZN(n566) );
  NAND2_X1 U630 ( .A1(G51), .A2(n628), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U634 ( .A(KEYINPUT7), .B(n571), .ZN(G168) );
  XOR2_X1 U635 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U636 ( .A1(G65), .A2(n629), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G53), .A2(n628), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n634), .A2(G78), .ZN(n575) );
  NAND2_X1 U640 ( .A1(G91), .A2(n633), .ZN(n574) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n713) );
  INV_X1 U643 ( .A(n713), .ZN(G299) );
  NOR2_X1 U644 ( .A1(G286), .A2(n649), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n578), .B(KEYINPUT78), .ZN(n580) );
  NOR2_X1 U646 ( .A1(G299), .A2(G868), .ZN(n579) );
  NOR2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U648 ( .A(KEYINPUT79), .B(n581), .Z(G297) );
  NAND2_X1 U649 ( .A1(G559), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n583), .B(KEYINPUT80), .ZN(n584) );
  INV_X1 U651 ( .A(n888), .ZN(n947) );
  NAND2_X1 U652 ( .A1(n584), .A2(n947), .ZN(n585) );
  XNOR2_X1 U653 ( .A(KEYINPUT16), .B(n585), .ZN(G148) );
  NOR2_X1 U654 ( .A1(G868), .A2(n940), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n947), .A2(G868), .ZN(n586) );
  NOR2_X1 U656 ( .A1(G559), .A2(n586), .ZN(n587) );
  NOR2_X1 U657 ( .A1(n588), .A2(n587), .ZN(G282) );
  XNOR2_X1 U658 ( .A(G2100), .B(KEYINPUT81), .ZN(n597) );
  NAND2_X1 U659 ( .A1(n869), .A2(G123), .ZN(n589) );
  XNOR2_X1 U660 ( .A(n589), .B(KEYINPUT18), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n868), .A2(G111), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G135), .A2(n874), .ZN(n593) );
  NAND2_X1 U664 ( .A1(G99), .A2(n872), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n921) );
  XNOR2_X1 U667 ( .A(n921), .B(G2096), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(G156) );
  NAND2_X1 U669 ( .A1(G559), .A2(n947), .ZN(n646) );
  XNOR2_X1 U670 ( .A(n940), .B(n646), .ZN(n598) );
  NOR2_X1 U671 ( .A1(G860), .A2(n598), .ZN(n606) );
  NAND2_X1 U672 ( .A1(G67), .A2(n629), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G93), .A2(n633), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U675 ( .A1(G55), .A2(n628), .ZN(n602) );
  NAND2_X1 U676 ( .A1(G80), .A2(n634), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n603) );
  OR2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n648) );
  XOR2_X1 U679 ( .A(n648), .B(KEYINPUT82), .Z(n605) );
  XNOR2_X1 U680 ( .A(n606), .B(n605), .ZN(G145) );
  NAND2_X1 U681 ( .A1(n634), .A2(G75), .ZN(n608) );
  NAND2_X1 U682 ( .A1(G88), .A2(n633), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U684 ( .A1(G62), .A2(n629), .ZN(n610) );
  NAND2_X1 U685 ( .A1(G50), .A2(n628), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U687 ( .A1(n612), .A2(n611), .ZN(G166) );
  NAND2_X1 U688 ( .A1(G61), .A2(n629), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G86), .A2(n633), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n634), .A2(G73), .ZN(n615) );
  XOR2_X1 U692 ( .A(KEYINPUT2), .B(n615), .Z(n616) );
  NOR2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n628), .A2(G48), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(G305) );
  NAND2_X1 U696 ( .A1(G49), .A2(n628), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G74), .A2(G651), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U699 ( .A1(n629), .A2(n622), .ZN(n626) );
  NAND2_X1 U700 ( .A1(G87), .A2(n623), .ZN(n624) );
  XOR2_X1 U701 ( .A(KEYINPUT83), .B(n624), .Z(n625) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U703 ( .A(KEYINPUT84), .B(n627), .ZN(G288) );
  NAND2_X1 U704 ( .A1(n628), .A2(G47), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n629), .A2(G60), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U707 ( .A(KEYINPUT70), .B(n632), .Z(n638) );
  NAND2_X1 U708 ( .A1(n633), .A2(G85), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n634), .A2(G72), .ZN(n635) );
  AND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n638), .A2(n637), .ZN(G290) );
  XOR2_X1 U712 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n640) );
  XNOR2_X1 U713 ( .A(n713), .B(G166), .ZN(n639) );
  XNOR2_X1 U714 ( .A(n640), .B(n639), .ZN(n641) );
  XOR2_X1 U715 ( .A(n648), .B(n641), .Z(n643) );
  XNOR2_X1 U716 ( .A(G305), .B(G288), .ZN(n642) );
  XNOR2_X1 U717 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U718 ( .A(n644), .B(G290), .ZN(n645) );
  XNOR2_X1 U719 ( .A(n645), .B(n940), .ZN(n889) );
  XNOR2_X1 U720 ( .A(n646), .B(n889), .ZN(n647) );
  NAND2_X1 U721 ( .A1(n647), .A2(G868), .ZN(n651) );
  NAND2_X1 U722 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n651), .A2(n650), .ZN(G295) );
  NAND2_X1 U724 ( .A1(G2078), .A2(G2084), .ZN(n653) );
  XOR2_X1 U725 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n652) );
  XNOR2_X1 U726 ( .A(n653), .B(n652), .ZN(n654) );
  NAND2_X1 U727 ( .A1(G2090), .A2(n654), .ZN(n655) );
  XNOR2_X1 U728 ( .A(KEYINPUT21), .B(n655), .ZN(n656) );
  NAND2_X1 U729 ( .A1(n656), .A2(G2072), .ZN(G158) );
  XOR2_X1 U730 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U731 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U732 ( .A1(G120), .A2(G108), .ZN(n657) );
  NOR2_X1 U733 ( .A1(G237), .A2(n657), .ZN(n658) );
  NAND2_X1 U734 ( .A1(G69), .A2(n658), .ZN(n820) );
  NAND2_X1 U735 ( .A1(n820), .A2(G567), .ZN(n663) );
  NOR2_X1 U736 ( .A1(G220), .A2(G219), .ZN(n659) );
  XOR2_X1 U737 ( .A(KEYINPUT22), .B(n659), .Z(n660) );
  NOR2_X1 U738 ( .A1(G218), .A2(n660), .ZN(n661) );
  NAND2_X1 U739 ( .A1(G96), .A2(n661), .ZN(n821) );
  NAND2_X1 U740 ( .A1(n821), .A2(G2106), .ZN(n662) );
  NAND2_X1 U741 ( .A1(n663), .A2(n662), .ZN(n822) );
  NAND2_X1 U742 ( .A1(G661), .A2(G483), .ZN(n664) );
  XOR2_X1 U743 ( .A(KEYINPUT87), .B(n664), .Z(n665) );
  NOR2_X1 U744 ( .A1(n822), .A2(n665), .ZN(n819) );
  NAND2_X1 U745 ( .A1(n819), .A2(G36), .ZN(G176) );
  NAND2_X1 U746 ( .A1(G138), .A2(n874), .ZN(n667) );
  NAND2_X1 U747 ( .A1(G126), .A2(n869), .ZN(n666) );
  NAND2_X1 U748 ( .A1(n667), .A2(n666), .ZN(n672) );
  NAND2_X1 U749 ( .A1(G102), .A2(n872), .ZN(n668) );
  XNOR2_X1 U750 ( .A(n668), .B(KEYINPUT88), .ZN(n670) );
  NAND2_X1 U751 ( .A1(n868), .A2(G114), .ZN(n669) );
  NAND2_X1 U752 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U753 ( .A1(n672), .A2(n671), .ZN(G164) );
  INV_X1 U754 ( .A(G166), .ZN(G303) );
  AND2_X1 U755 ( .A1(n673), .A2(G40), .ZN(n674) );
  NAND2_X1 U756 ( .A1(n675), .A2(n674), .ZN(n769) );
  INV_X1 U757 ( .A(n769), .ZN(n677) );
  INV_X1 U758 ( .A(KEYINPUT95), .ZN(n676) );
  NAND2_X1 U759 ( .A1(n677), .A2(n676), .ZN(n679) );
  NAND2_X1 U760 ( .A1(KEYINPUT95), .A2(n769), .ZN(n678) );
  NAND2_X1 U761 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U762 ( .A1(G164), .A2(G1384), .ZN(n770) );
  NAND2_X1 U763 ( .A1(G8), .A2(n732), .ZN(n757) );
  NOR2_X1 U764 ( .A1(G1976), .A2(G288), .ZN(n744) );
  NAND2_X1 U765 ( .A1(n744), .A2(KEYINPUT33), .ZN(n681) );
  NOR2_X1 U766 ( .A1(n757), .A2(n681), .ZN(n749) );
  NAND2_X1 U767 ( .A1(G1976), .A2(G288), .ZN(n944) );
  INV_X1 U768 ( .A(n944), .ZN(n682) );
  OR2_X1 U769 ( .A1(n682), .A2(n757), .ZN(n683) );
  INV_X1 U770 ( .A(n683), .ZN(n746) );
  NOR2_X1 U771 ( .A1(G1966), .A2(n757), .ZN(n685) );
  INV_X1 U772 ( .A(n685), .ZN(n726) );
  NOR2_X1 U773 ( .A1(G2084), .A2(n732), .ZN(n684) );
  XOR2_X1 U774 ( .A(n684), .B(KEYINPUT96), .Z(n727) );
  INV_X1 U775 ( .A(G8), .ZN(n686) );
  NOR2_X1 U776 ( .A1(n686), .A2(n685), .ZN(n687) );
  AND2_X1 U777 ( .A1(n727), .A2(n687), .ZN(n688) );
  XOR2_X1 U778 ( .A(n688), .B(KEYINPUT30), .Z(n689) );
  NOR2_X1 U779 ( .A1(G168), .A2(n689), .ZN(n693) );
  XOR2_X1 U780 ( .A(KEYINPUT25), .B(G2078), .Z(n965) );
  NOR2_X1 U781 ( .A1(n965), .A2(n732), .ZN(n691) );
  INV_X1 U782 ( .A(n732), .ZN(n708) );
  NOR2_X1 U783 ( .A1(n708), .A2(G1961), .ZN(n690) );
  NOR2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n720) );
  AND2_X1 U785 ( .A1(G301), .A2(n720), .ZN(n692) );
  NOR2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U787 ( .A(n694), .B(KEYINPUT31), .ZN(n724) );
  INV_X1 U788 ( .A(G1996), .ZN(n841) );
  NOR2_X1 U789 ( .A1(n732), .A2(n841), .ZN(n695) );
  XNOR2_X1 U790 ( .A(n695), .B(KEYINPUT26), .ZN(n697) );
  AND2_X1 U791 ( .A1(n732), .A2(G1341), .ZN(n696) );
  OR2_X1 U792 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U793 ( .A1(n940), .A2(n698), .ZN(n703) );
  NAND2_X1 U794 ( .A1(n703), .A2(n947), .ZN(n702) );
  NAND2_X1 U795 ( .A1(G1348), .A2(n732), .ZN(n700) );
  NAND2_X1 U796 ( .A1(G2067), .A2(n708), .ZN(n699) );
  NAND2_X1 U797 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U798 ( .A1(n702), .A2(n701), .ZN(n705) );
  OR2_X1 U799 ( .A1(n703), .A2(n947), .ZN(n704) );
  NAND2_X1 U800 ( .A1(n705), .A2(n704), .ZN(n712) );
  XOR2_X1 U801 ( .A(KEYINPUT97), .B(KEYINPUT27), .Z(n707) );
  NAND2_X1 U802 ( .A1(G2072), .A2(n708), .ZN(n706) );
  XNOR2_X1 U803 ( .A(n707), .B(n706), .ZN(n710) );
  INV_X1 U804 ( .A(G1956), .ZN(n999) );
  NOR2_X1 U805 ( .A1(n708), .A2(n999), .ZN(n709) );
  NOR2_X1 U806 ( .A1(n710), .A2(n709), .ZN(n714) );
  NAND2_X1 U807 ( .A1(n714), .A2(n713), .ZN(n711) );
  NAND2_X1 U808 ( .A1(n712), .A2(n711), .ZN(n718) );
  NOR2_X1 U809 ( .A1(n714), .A2(n713), .ZN(n716) );
  XOR2_X1 U810 ( .A(KEYINPUT28), .B(KEYINPUT98), .Z(n715) );
  XNOR2_X1 U811 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U813 ( .A(n719), .B(KEYINPUT29), .ZN(n722) );
  NOR2_X1 U814 ( .A1(G301), .A2(n720), .ZN(n721) );
  NOR2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U816 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U817 ( .A(KEYINPUT99), .B(n725), .ZN(n736) );
  AND2_X1 U818 ( .A1(n726), .A2(n736), .ZN(n730) );
  INV_X1 U819 ( .A(n727), .ZN(n728) );
  NAND2_X1 U820 ( .A1(G8), .A2(n728), .ZN(n729) );
  NAND2_X1 U821 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U822 ( .A(KEYINPUT100), .B(n731), .ZN(n742) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n757), .ZN(n734) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U826 ( .A1(n735), .A2(G303), .ZN(n738) );
  NAND2_X1 U827 ( .A1(G286), .A2(n736), .ZN(n737) );
  NAND2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U829 ( .A1(G8), .A2(n739), .ZN(n740) );
  XNOR2_X1 U830 ( .A(KEYINPUT32), .B(n740), .ZN(n741) );
  NAND2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n753) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n743) );
  NOR2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n948) );
  NAND2_X1 U834 ( .A1(n753), .A2(n948), .ZN(n745) );
  AND2_X1 U835 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U836 ( .A1(KEYINPUT33), .A2(n747), .ZN(n748) );
  NOR2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U838 ( .A(G1981), .B(G305), .Z(n936) );
  AND2_X1 U839 ( .A1(n750), .A2(n936), .ZN(n805) );
  NOR2_X1 U840 ( .A1(G2090), .A2(G303), .ZN(n751) );
  NAND2_X1 U841 ( .A1(G8), .A2(n751), .ZN(n752) );
  NAND2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n754), .A2(n757), .ZN(n759) );
  NOR2_X1 U844 ( .A1(G1981), .A2(G305), .ZN(n755) );
  XOR2_X1 U845 ( .A(n755), .B(KEYINPUT24), .Z(n756) );
  OR2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U847 ( .A1(n759), .A2(n758), .ZN(n803) );
  NAND2_X1 U848 ( .A1(n872), .A2(G105), .ZN(n761) );
  XNOR2_X1 U849 ( .A(KEYINPUT38), .B(KEYINPUT92), .ZN(n760) );
  XNOR2_X1 U850 ( .A(n761), .B(n760), .ZN(n768) );
  NAND2_X1 U851 ( .A1(G117), .A2(n868), .ZN(n763) );
  NAND2_X1 U852 ( .A1(G129), .A2(n869), .ZN(n762) );
  NAND2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n766) );
  NAND2_X1 U854 ( .A1(G141), .A2(n874), .ZN(n764) );
  XNOR2_X1 U855 ( .A(KEYINPUT93), .B(n764), .ZN(n765) );
  NOR2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n881) );
  NOR2_X1 U858 ( .A1(G1996), .A2(n881), .ZN(n918) );
  NOR2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n806) );
  NAND2_X1 U860 ( .A1(G1996), .A2(n881), .ZN(n779) );
  NAND2_X1 U861 ( .A1(G131), .A2(n874), .ZN(n772) );
  NAND2_X1 U862 ( .A1(G107), .A2(n868), .ZN(n771) );
  NAND2_X1 U863 ( .A1(n772), .A2(n771), .ZN(n775) );
  NAND2_X1 U864 ( .A1(G119), .A2(n869), .ZN(n773) );
  XNOR2_X1 U865 ( .A(KEYINPUT91), .B(n773), .ZN(n774) );
  NOR2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U867 ( .A1(n872), .A2(G95), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n861) );
  NAND2_X1 U869 ( .A1(G1991), .A2(n861), .ZN(n778) );
  NAND2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U871 ( .A(KEYINPUT94), .B(n780), .Z(n925) );
  INV_X1 U872 ( .A(n925), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n806), .A2(n781), .ZN(n807) );
  INV_X1 U874 ( .A(n807), .ZN(n784) );
  NOR2_X1 U875 ( .A1(G1991), .A2(n861), .ZN(n922) );
  NOR2_X1 U876 ( .A1(G1986), .A2(G290), .ZN(n782) );
  NOR2_X1 U877 ( .A1(n922), .A2(n782), .ZN(n783) );
  NOR2_X1 U878 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U879 ( .A1(n918), .A2(n785), .ZN(n786) );
  XNOR2_X1 U880 ( .A(KEYINPUT39), .B(n786), .ZN(n798) );
  XOR2_X1 U881 ( .A(G2067), .B(KEYINPUT37), .Z(n799) );
  NAND2_X1 U882 ( .A1(G140), .A2(n874), .ZN(n788) );
  NAND2_X1 U883 ( .A1(G104), .A2(n872), .ZN(n787) );
  NAND2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U885 ( .A(KEYINPUT34), .B(n789), .ZN(n795) );
  NAND2_X1 U886 ( .A1(G128), .A2(n869), .ZN(n790) );
  XOR2_X1 U887 ( .A(KEYINPUT89), .B(n790), .Z(n792) );
  NAND2_X1 U888 ( .A1(n868), .A2(G116), .ZN(n791) );
  NAND2_X1 U889 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U890 ( .A(KEYINPUT35), .B(n793), .Z(n794) );
  NOR2_X1 U891 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U892 ( .A(KEYINPUT36), .B(n796), .Z(n864) );
  NAND2_X1 U893 ( .A1(n799), .A2(n864), .ZN(n797) );
  XOR2_X1 U894 ( .A(KEYINPUT90), .B(n797), .Z(n916) );
  NAND2_X1 U895 ( .A1(n806), .A2(n916), .ZN(n808) );
  NAND2_X1 U896 ( .A1(n798), .A2(n808), .ZN(n800) );
  OR2_X1 U897 ( .A1(n799), .A2(n864), .ZN(n913) );
  NAND2_X1 U898 ( .A1(n800), .A2(n913), .ZN(n801) );
  NAND2_X1 U899 ( .A1(n801), .A2(n806), .ZN(n812) );
  INV_X1 U900 ( .A(n812), .ZN(n802) );
  OR2_X1 U901 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U902 ( .A1(n805), .A2(n804), .ZN(n814) );
  XNOR2_X1 U903 ( .A(G1986), .B(G290), .ZN(n955) );
  AND2_X1 U904 ( .A1(n955), .A2(n806), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n809) );
  OR2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n811) );
  AND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U909 ( .A(n815), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n816), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U912 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(G188) );
  XOR2_X1 U915 ( .A(G108), .B(KEYINPUT110), .Z(G238) );
  INV_X1 U917 ( .A(G120), .ZN(G236) );
  INV_X1 U918 ( .A(G96), .ZN(G221) );
  INV_X1 U919 ( .A(G69), .ZN(G235) );
  NOR2_X1 U920 ( .A1(n821), .A2(n820), .ZN(G325) );
  INV_X1 U921 ( .A(G325), .ZN(G261) );
  INV_X1 U922 ( .A(n822), .ZN(G319) );
  XOR2_X1 U923 ( .A(G2100), .B(KEYINPUT43), .Z(n824) );
  XNOR2_X1 U924 ( .A(G2090), .B(G2678), .ZN(n823) );
  XNOR2_X1 U925 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U926 ( .A(n825), .B(KEYINPUT102), .Z(n827) );
  XNOR2_X1 U927 ( .A(G2067), .B(G2072), .ZN(n826) );
  XNOR2_X1 U928 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U929 ( .A(KEYINPUT42), .B(G2096), .Z(n829) );
  XNOR2_X1 U930 ( .A(G2078), .B(G2084), .ZN(n828) );
  XNOR2_X1 U931 ( .A(n829), .B(n828), .ZN(n830) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(G227) );
  XOR2_X1 U933 ( .A(G1976), .B(G1971), .Z(n833) );
  XNOR2_X1 U934 ( .A(G1991), .B(G1986), .ZN(n832) );
  XNOR2_X1 U935 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U936 ( .A(G1981), .B(G1956), .Z(n835) );
  XNOR2_X1 U937 ( .A(G1966), .B(G1961), .ZN(n834) );
  XNOR2_X1 U938 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U939 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U940 ( .A(G2474), .B(KEYINPUT41), .ZN(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U942 ( .A(KEYINPUT103), .B(n840), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(G229) );
  NAND2_X1 U944 ( .A1(n869), .A2(G124), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n843), .B(KEYINPUT44), .ZN(n844) );
  XNOR2_X1 U946 ( .A(KEYINPUT104), .B(n844), .ZN(n847) );
  NAND2_X1 U947 ( .A1(G136), .A2(n874), .ZN(n845) );
  XOR2_X1 U948 ( .A(KEYINPUT105), .B(n845), .Z(n846) );
  NAND2_X1 U949 ( .A1(n847), .A2(n846), .ZN(n851) );
  NAND2_X1 U950 ( .A1(G112), .A2(n868), .ZN(n849) );
  NAND2_X1 U951 ( .A1(G100), .A2(n872), .ZN(n848) );
  NAND2_X1 U952 ( .A1(n849), .A2(n848), .ZN(n850) );
  NOR2_X1 U953 ( .A1(n851), .A2(n850), .ZN(G162) );
  NAND2_X1 U954 ( .A1(G139), .A2(n874), .ZN(n853) );
  NAND2_X1 U955 ( .A1(G103), .A2(n872), .ZN(n852) );
  NAND2_X1 U956 ( .A1(n853), .A2(n852), .ZN(n859) );
  NAND2_X1 U957 ( .A1(G115), .A2(n868), .ZN(n855) );
  NAND2_X1 U958 ( .A1(G127), .A2(n869), .ZN(n854) );
  NAND2_X1 U959 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U960 ( .A(KEYINPUT47), .B(n856), .ZN(n857) );
  XNOR2_X1 U961 ( .A(KEYINPUT107), .B(n857), .ZN(n858) );
  NOR2_X1 U962 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U963 ( .A(KEYINPUT108), .B(n860), .Z(n909) );
  XNOR2_X1 U964 ( .A(n909), .B(n921), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n864), .B(n863), .ZN(n886) );
  XOR2_X1 U967 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n866) );
  XNOR2_X1 U968 ( .A(G162), .B(KEYINPUT109), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U970 ( .A(G164), .B(n867), .ZN(n884) );
  NAND2_X1 U971 ( .A1(G118), .A2(n868), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G130), .A2(n869), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n879) );
  NAND2_X1 U974 ( .A1(n872), .A2(G106), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n873), .B(KEYINPUT106), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G142), .A2(n874), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U978 ( .A(KEYINPUT45), .B(n877), .Z(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U980 ( .A(G160), .B(n880), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n886), .B(n885), .ZN(n887) );
  NOR2_X1 U984 ( .A1(G37), .A2(n887), .ZN(G395) );
  XNOR2_X1 U985 ( .A(n888), .B(G286), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n891), .B(G171), .ZN(n892) );
  NOR2_X1 U988 ( .A1(G37), .A2(n892), .ZN(G397) );
  XOR2_X1 U989 ( .A(G2454), .B(G2435), .Z(n894) );
  XNOR2_X1 U990 ( .A(G2438), .B(G2427), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n901) );
  XOR2_X1 U992 ( .A(KEYINPUT101), .B(G2446), .Z(n896) );
  XNOR2_X1 U993 ( .A(G2443), .B(G2430), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U995 ( .A(n897), .B(G2451), .Z(n899) );
  XNOR2_X1 U996 ( .A(G1348), .B(G1341), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  NAND2_X1 U999 ( .A1(n902), .A2(G14), .ZN(n908) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n908), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n903), .ZN(n904) );
  NOR2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(n908), .ZN(G401) );
  XNOR2_X1 U1008 ( .A(KEYINPUT55), .B(KEYINPUT113), .ZN(n982) );
  XOR2_X1 U1009 ( .A(G164), .B(G2078), .Z(n911) );
  XNOR2_X1 U1010 ( .A(G2072), .B(n909), .ZN(n910) );
  NOR2_X1 U1011 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n912), .B(KEYINPUT50), .ZN(n914) );
  NAND2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(n930) );
  XOR2_X1 U1015 ( .A(G2090), .B(G162), .Z(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(KEYINPUT51), .B(n919), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(n920), .B(KEYINPUT111), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n928) );
  XNOR2_X1 U1021 ( .A(G2084), .B(G160), .ZN(n926) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1024 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1025 ( .A(KEYINPUT52), .B(n931), .ZN(n932) );
  XOR2_X1 U1026 ( .A(KEYINPUT112), .B(n932), .Z(n933) );
  NAND2_X1 U1027 ( .A1(n982), .A2(n933), .ZN(n934) );
  NAND2_X1 U1028 ( .A1(n934), .A2(G29), .ZN(n990) );
  XOR2_X1 U1029 ( .A(G16), .B(KEYINPUT118), .Z(n935) );
  XNOR2_X1 U1030 ( .A(KEYINPUT56), .B(n935), .ZN(n961) );
  XNOR2_X1 U1031 ( .A(G1966), .B(G168), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(n938), .B(KEYINPUT57), .ZN(n942) );
  XOR2_X1 U1034 ( .A(G1341), .B(KEYINPUT120), .Z(n939) );
  XNOR2_X1 U1035 ( .A(n940), .B(n939), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n958) );
  NAND2_X1 U1037 ( .A1(G1971), .A2(G303), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n946) );
  XNOR2_X1 U1039 ( .A(G1956), .B(G299), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n953) );
  XNOR2_X1 U1041 ( .A(G1348), .B(n947), .ZN(n949) );
  NAND2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(G1961), .B(G301), .ZN(n950) );
  NOR2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(n956), .B(KEYINPUT119), .ZN(n957) );
  NOR2_X1 U1048 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1049 ( .A(KEYINPUT121), .B(n959), .Z(n960) );
  NOR2_X1 U1050 ( .A1(n961), .A2(n960), .ZN(n988) );
  XNOR2_X1 U1051 ( .A(KEYINPUT54), .B(KEYINPUT115), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(n962), .B(G34), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(G2084), .B(n963), .ZN(n979) );
  XNOR2_X1 U1054 ( .A(G2090), .B(G35), .ZN(n977) );
  XOR2_X1 U1055 ( .A(G1991), .B(G25), .Z(n964) );
  NAND2_X1 U1056 ( .A1(n964), .A2(G28), .ZN(n974) );
  XNOR2_X1 U1057 ( .A(G1996), .B(G32), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(n965), .B(G27), .ZN(n966) );
  NOR2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(KEYINPUT114), .B(n968), .ZN(n972) );
  XNOR2_X1 U1061 ( .A(G2067), .B(G26), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(G33), .B(G2072), .ZN(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(KEYINPUT53), .B(n975), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(n980), .B(KEYINPUT116), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(n982), .B(n981), .ZN(n984) );
  INV_X1 U1071 ( .A(G29), .ZN(n983) );
  NAND2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1073 ( .A1(n985), .A2(G11), .ZN(n986) );
  XOR2_X1 U1074 ( .A(KEYINPUT117), .B(n986), .Z(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1076 ( .A1(n990), .A2(n989), .ZN(n1020) );
  XNOR2_X1 U1077 ( .A(G1986), .B(G24), .ZN(n995) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G22), .ZN(n992) );
  XNOR2_X1 U1079 ( .A(G1976), .B(G23), .ZN(n991) );
  NOR2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(KEYINPUT127), .B(n993), .ZN(n994) );
  NOR2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1083 ( .A(KEYINPUT58), .B(n996), .Z(n1016) );
  XNOR2_X1 U1084 ( .A(G1961), .B(G5), .ZN(n1013) );
  XOR2_X1 U1085 ( .A(KEYINPUT124), .B(G4), .Z(n998) );
  XNOR2_X1 U1086 ( .A(G1348), .B(KEYINPUT59), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n998), .B(n997), .ZN(n1007) );
  XNOR2_X1 U1088 ( .A(G20), .B(n999), .ZN(n1002) );
  XOR2_X1 U1089 ( .A(G1341), .B(G19), .Z(n1000) );
  XNOR2_X1 U1090 ( .A(KEYINPUT122), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G6), .B(G1981), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1005), .B(KEYINPUT123), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1096 ( .A(KEYINPUT60), .B(n1008), .Z(n1010) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G21), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(KEYINPUT125), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1101 ( .A(KEYINPUT126), .B(n1014), .Z(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1017), .Z(n1018) );
  NOR2_X1 U1104 ( .A1(G16), .A2(n1018), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(n1021), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

