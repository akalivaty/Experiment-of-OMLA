//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049;
  XOR2_X1   g000(.A(KEYINPUT75), .B(KEYINPUT27), .Z(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G101), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT2), .B(G113), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G116), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT71), .B(G119), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G116), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT70), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n194), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(KEYINPUT71), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT71), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G119), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n203), .A3(G116), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(G116), .B2(new_n195), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT70), .A3(new_n193), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n200), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G137), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT11), .A3(G134), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G131), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n211), .A2(new_n213), .A3(new_n217), .A4(new_n214), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G143), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT0), .A2(G128), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n220), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G143), .B(G146), .ZN(new_n228));
  INV_X1    g042(.A(new_n226), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(KEYINPUT64), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n227), .A2(new_n230), .B1(new_n225), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n219), .B1(new_n233), .B2(KEYINPUT65), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n225), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT64), .B1(new_n228), .B2(new_n229), .ZN(new_n236));
  AND4_X1   g050(.A1(KEYINPUT64), .A2(new_n229), .A3(new_n222), .A4(new_n224), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT66), .B1(new_n234), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n222), .A2(new_n224), .A3(G128), .ZN(new_n242));
  OR2_X1    g056(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT68), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n247));
  NOR2_X1   g061(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n249), .A2(new_n228), .A3(new_n250), .A4(G128), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n223), .B(G146), .C1(new_n247), .C2(new_n248), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n253), .B(new_n254), .C1(G128), .C2(new_n228), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n223), .A2(G146), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(new_n243), .B2(new_n244), .ZN(new_n257));
  AOI21_X1  g071(.A(G128), .B1(new_n222), .B2(new_n224), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT69), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n252), .A2(new_n255), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n214), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n210), .A2(G137), .ZN(new_n262));
  OAI21_X1  g076(.A(G131), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n263), .A2(new_n218), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n238), .A2(new_n239), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n227), .A2(new_n230), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT65), .A3(new_n235), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT66), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n266), .A2(new_n268), .A3(new_n269), .A4(new_n219), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n241), .A2(new_n265), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT30), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n208), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n260), .A2(new_n274), .A3(new_n264), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n274), .B1(new_n260), .B2(new_n264), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n238), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n267), .A2(KEYINPUT72), .A3(new_n235), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n280), .A3(new_n219), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT30), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT74), .B1(new_n277), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n285));
  NOR4_X1   g099(.A1(new_n282), .A2(new_n275), .A3(new_n276), .A4(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n273), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n265), .A2(KEYINPUT73), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n260), .A2(new_n274), .A3(new_n264), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n208), .A3(new_n281), .A4(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n192), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n271), .A2(new_n207), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n290), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n192), .B(KEYINPUT76), .Z(new_n296));
  NAND3_X1  g110(.A1(new_n281), .A2(new_n265), .A3(new_n208), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n293), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n292), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT77), .B1(new_n291), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n266), .A2(new_n268), .A3(new_n219), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n302), .A2(KEYINPUT66), .B1(new_n260), .B2(new_n264), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n208), .B1(new_n303), .B2(new_n270), .ZN(new_n304));
  AND4_X1   g118(.A1(new_n208), .A2(new_n288), .A3(new_n281), .A4(new_n289), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT28), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n298), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n192), .B(KEYINPUT76), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT29), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n288), .A2(new_n289), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n285), .B1(new_n312), .B2(new_n282), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n277), .A2(new_n283), .A3(KEYINPUT74), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n305), .B1(new_n315), .B2(new_n273), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n310), .B(new_n311), .C1(new_n192), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n277), .A2(new_n281), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n207), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n290), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n307), .B1(new_n320), .B2(KEYINPUT28), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n192), .A2(KEYINPUT29), .ZN(new_n322));
  AOI21_X1  g136(.A(G902), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n301), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G472), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n290), .A2(new_n192), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n287), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT31), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n287), .A2(KEYINPUT31), .A3(new_n329), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n306), .A2(new_n298), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n332), .A2(new_n333), .B1(new_n308), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(G472), .A2(G902), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT32), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n308), .ZN(new_n339));
  AOI211_X1 g153(.A(new_n331), .B(new_n328), .C1(new_n315), .C2(new_n273), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT31), .B1(new_n287), .B2(new_n329), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT32), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n343), .A3(new_n336), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n324), .A2(KEYINPUT78), .A3(G472), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n327), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT82), .B(KEYINPUT25), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n197), .A2(G128), .ZN(new_n350));
  INV_X1    g164(.A(G128), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G119), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT24), .B(G110), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(KEYINPUT23), .A3(G119), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(KEYINPUT79), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n197), .A2(G128), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n357), .B(new_n350), .C1(KEYINPUT23), .C2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n355), .B1(new_n359), .B2(G110), .ZN(new_n360));
  INV_X1    g174(.A(G140), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G125), .ZN(new_n362));
  INV_X1    g176(.A(G125), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G140), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n364), .A3(KEYINPUT80), .ZN(new_n365));
  OR3_X1    g179(.A1(new_n361), .A2(KEYINPUT80), .A3(G125), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(KEYINPUT16), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT16), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G146), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n367), .A2(new_n221), .A3(new_n369), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(KEYINPUT81), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT81), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(new_n374), .A3(G146), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n360), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n353), .A2(new_n354), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n377), .B1(new_n359), .B2(G110), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n362), .A2(new_n364), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n221), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n371), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT22), .B(G137), .ZN(new_n382));
  INV_X1    g196(.A(G953), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(G221), .A3(G234), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n382), .B(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n376), .A2(new_n381), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n385), .B1(new_n376), .B2(new_n381), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G902), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n349), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n376), .A2(new_n381), .ZN(new_n392));
  INV_X1    g206(.A(new_n385), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT25), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n394), .A2(new_n395), .A3(new_n390), .A4(new_n386), .ZN(new_n396));
  INV_X1    g210(.A(G217), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(G234), .B2(new_n390), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT83), .B1(new_n391), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n394), .A2(new_n386), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n348), .B1(new_n401), .B2(G902), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n396), .A4(new_n398), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n398), .A2(G902), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n389), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n400), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G214), .B1(G237), .B2(G902), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT90), .B1(new_n233), .B2(new_n363), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n252), .A2(new_n363), .A3(new_n255), .A4(new_n259), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT90), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n238), .A2(new_n413), .A3(G125), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G224), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(G953), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n415), .B(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G104), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT3), .B1(new_n419), .B2(G107), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT3), .ZN(new_n421));
  INV_X1    g235(.A(G107), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n422), .A3(G104), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n419), .A2(G107), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n420), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n425), .A2(G101), .ZN(new_n426));
  INV_X1    g240(.A(G101), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n420), .A2(new_n423), .A3(new_n427), .A4(new_n424), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT4), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT85), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(G101), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT4), .A4(new_n428), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT86), .B(KEYINPUT4), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n200), .A2(new_n206), .B1(new_n426), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT5), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n197), .A2(new_n438), .A3(G116), .ZN(new_n439));
  OAI211_X1 g253(.A(G113), .B(new_n439), .C1(new_n205), .C2(new_n438), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT87), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n205), .A2(new_n193), .ZN(new_n443));
  INV_X1    g257(.A(new_n424), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n419), .A2(G107), .ZN(new_n445));
  OAI21_X1  g259(.A(G101), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n428), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n198), .A2(KEYINPUT5), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n449), .A2(KEYINPUT87), .A3(G113), .A4(new_n439), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n442), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n437), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n453));
  XNOR2_X1  g267(.A(G110), .B(G122), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT89), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n452), .A2(new_n458), .A3(new_n453), .A4(new_n455), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT88), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n452), .A2(new_n455), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n437), .A2(new_n451), .A3(new_n454), .ZN(new_n463));
  AND4_X1   g277(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT6), .A4(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n453), .B1(new_n452), .B2(new_n455), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n461), .B1(new_n465), .B2(new_n463), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n418), .B(new_n460), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n415), .A2(new_n417), .ZN(new_n468));
  INV_X1    g282(.A(new_n417), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT91), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT7), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n470), .B2(new_n469), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n411), .A2(new_n412), .A3(new_n414), .A4(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT7), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n415), .A2(new_n474), .ZN(new_n475));
  AND4_X1   g289(.A1(new_n468), .A2(new_n463), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n442), .A2(new_n450), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n447), .B1(new_n477), .B2(new_n443), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n448), .A2(new_n440), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n454), .B(KEYINPUT8), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(G902), .B1(new_n476), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n467), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G210), .B1(G237), .B2(G902), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n467), .A2(new_n485), .A3(new_n483), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n410), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G113), .B(G122), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(new_n419), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n495));
  OAI21_X1  g309(.A(G131), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT17), .ZN(new_n497));
  INV_X1    g311(.A(G237), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n383), .A3(G214), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n223), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n217), .A3(new_n493), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n496), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT93), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT93), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n496), .A2(new_n504), .A3(new_n497), .A4(new_n501), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n493), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT17), .A3(G131), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(new_n375), .B2(new_n373), .ZN(new_n509));
  NAND2_X1  g323(.A1(KEYINPUT18), .A2(G131), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n506), .B(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n365), .A2(G146), .A3(new_n366), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n380), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n492), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT94), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n503), .A2(new_n505), .A3(new_n507), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n373), .A2(new_n375), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n491), .A3(new_n514), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n516), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n390), .B1(new_n516), .B2(new_n517), .ZN(new_n523));
  OAI21_X1  g337(.A(G475), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(G475), .A2(G902), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n492), .B(new_n515), .C1(new_n518), .C2(new_n519), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT92), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n370), .A2(G146), .B1(new_n496), .B2(new_n501), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT19), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n365), .B2(new_n366), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n379), .A2(KEYINPUT19), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n221), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n528), .A2(new_n532), .B1(new_n511), .B2(new_n513), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n527), .B1(new_n533), .B2(new_n491), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n496), .A2(new_n501), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n371), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n514), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT92), .A3(new_n492), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n525), .B1(new_n526), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT20), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n521), .A2(new_n538), .A3(new_n534), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(new_n525), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n524), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n351), .B2(G143), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n223), .A2(KEYINPUT95), .A3(G128), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(G128), .B2(new_n223), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G134), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n550), .B(new_n210), .C1(G128), .C2(new_n223), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G116), .B(G122), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G122), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G116), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n422), .B1(new_n558), .B2(KEYINPUT14), .ZN(new_n559));
  OR2_X1    g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n556), .A2(new_n559), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n554), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT9), .B(G234), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n563), .A2(new_n397), .A3(G953), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n223), .A2(G128), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT13), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n565), .B1(new_n550), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT96), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n548), .A2(KEYINPUT13), .A3(new_n549), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT13), .B1(new_n548), .B2(new_n549), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT96), .B1(new_n571), .B2(new_n565), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n573), .A2(G134), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n555), .A2(G107), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n556), .A2(new_n422), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n553), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n562), .B(new_n564), .C1(new_n574), .C2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n564), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n577), .B1(new_n573), .B2(G134), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n554), .A2(new_n560), .A3(new_n561), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n390), .ZN(new_n584));
  INV_X1    g398(.A(G478), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(KEYINPUT15), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n584), .B(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n383), .A2(G952), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(G234), .B2(G237), .ZN(new_n591));
  AOI211_X1 g405(.A(new_n390), .B(new_n383), .C1(G234), .C2(G237), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT21), .B(G898), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n546), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(G221), .B1(new_n563), .B2(G902), .ZN(new_n596));
  XOR2_X1   g410(.A(new_n596), .B(KEYINPUT84), .Z(new_n597));
  INV_X1    g411(.A(G469), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n390), .ZN(new_n599));
  XNOR2_X1  g413(.A(G110), .B(G140), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n383), .A2(G227), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n224), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n258), .B1(KEYINPUT1), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n252), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n447), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n447), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n607), .A2(new_n608), .B1(new_n260), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n426), .A2(new_n435), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n434), .A2(new_n279), .A3(new_n280), .A4(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n219), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n613), .B1(new_n610), .B2(new_n612), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n602), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n617));
  INV_X1    g431(.A(new_n602), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n252), .A2(new_n255), .A3(new_n259), .A4(new_n447), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n613), .B1(new_n607), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(KEYINPUT12), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT12), .ZN(new_n622));
  AOI211_X1 g436(.A(new_n622), .B(new_n613), .C1(new_n607), .C2(new_n619), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n617), .B(new_n618), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(G902), .B1(new_n616), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n599), .B1(new_n625), .B2(new_n598), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n621), .A2(new_n623), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n602), .B1(new_n627), .B2(new_n614), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n610), .A2(new_n612), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n219), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(new_n617), .A3(new_n618), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n628), .A2(G469), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n597), .B1(new_n626), .B2(new_n632), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n489), .A2(new_n595), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n347), .A2(new_n408), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  NAND2_X1  g450(.A1(new_n408), .A2(new_n633), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n342), .A2(new_n336), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(G472), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n342), .B2(new_n390), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n637), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n546), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT97), .B1(new_n580), .B2(new_n581), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT33), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n583), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n578), .A2(new_n582), .A3(new_n644), .A4(KEYINPUT33), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n585), .A2(G902), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT98), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n646), .A2(KEYINPUT98), .A3(new_n647), .A4(new_n648), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT99), .B(G478), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n651), .A2(new_n652), .B1(new_n584), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n643), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n594), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n489), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n642), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G104), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  NOR2_X1   g475(.A1(new_n546), .A2(new_n588), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n489), .A2(new_n656), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n642), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT101), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT35), .B(G107), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  OAI21_X1  g481(.A(G472), .B1(new_n335), .B2(G902), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n393), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT102), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n392), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n405), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n400), .A2(new_n404), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n668), .A2(new_n638), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT103), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n668), .A2(new_n676), .A3(new_n638), .A4(new_n673), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n675), .A2(new_n634), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  INV_X1    g494(.A(G900), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n591), .B1(new_n592), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n662), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n626), .A2(new_n632), .ZN(new_n685));
  INV_X1    g499(.A(new_n597), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n673), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n467), .A2(new_n485), .A3(new_n483), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n485), .B1(new_n467), .B2(new_n483), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n409), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n684), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n347), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  XNOR2_X1  g507(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n682), .B(new_n694), .Z(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n633), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT40), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n487), .A2(new_n488), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT38), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n487), .A2(KEYINPUT38), .A3(new_n488), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n320), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n330), .B1(new_n706), .B2(new_n296), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n390), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(G472), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n342), .A2(new_n343), .A3(new_n336), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n343), .B1(new_n342), .B2(new_n336), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n400), .A2(new_n404), .A3(new_n672), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n588), .B1(new_n524), .B2(new_n545), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n713), .A2(new_n409), .A3(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n699), .A2(new_n705), .A3(new_n712), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  NAND2_X1  g531(.A1(new_n651), .A2(new_n652), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n584), .A2(new_n653), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n546), .A3(new_n683), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n687), .A2(new_n690), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n347), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G146), .ZN(G48));
  OAI21_X1  g538(.A(new_n346), .B1(new_n711), .B2(new_n710), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT78), .B1(new_n324), .B2(G472), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n625), .A2(new_n598), .ZN(new_n728));
  AOI211_X1 g542(.A(G469), .B(G902), .C1(new_n616), .C2(new_n624), .ZN(new_n729));
  INV_X1    g543(.A(new_n596), .ZN(new_n730));
  OR3_X1    g544(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n407), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n489), .A3(new_n655), .A4(new_n656), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT41), .B(G113), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  NAND4_X1  g550(.A1(new_n732), .A2(new_n489), .A3(new_n656), .A4(new_n662), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n727), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g552(.A(new_n738), .B(G116), .Z(G18));
  NOR3_X1   g553(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n740));
  AND4_X1   g554(.A1(new_n489), .A2(new_n595), .A3(new_n673), .A4(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n725), .B2(new_n726), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  NAND2_X1  g557(.A1(new_n342), .A2(new_n390), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT106), .B1(new_n744), .B2(G472), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  AOI211_X1 g560(.A(new_n746), .B(new_n640), .C1(new_n342), .C2(new_n390), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  OAI22_X1  g562(.A1(new_n340), .A2(new_n341), .B1(new_n321), .B2(new_n296), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n336), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(KEYINPUT105), .A3(new_n336), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n714), .B(new_n409), .C1(new_n688), .C2(new_n689), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n740), .A2(new_n656), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n748), .A2(new_n408), .A3(new_n754), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  NOR3_X1   g573(.A1(new_n690), .A2(new_n721), .A3(new_n731), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n748), .A2(new_n760), .A3(new_n673), .A4(new_n754), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  NAND3_X1  g576(.A1(new_n487), .A2(new_n409), .A3(new_n488), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n617), .A2(new_n618), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT107), .B1(new_n764), .B2(new_n615), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n630), .A2(new_n766), .A3(new_n617), .A4(new_n618), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(G469), .A3(new_n628), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n626), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n596), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n763), .A2(new_n721), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n347), .A2(new_n408), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n347), .A2(KEYINPUT42), .A3(new_n408), .A4(new_n772), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G131), .ZN(G33));
  NOR3_X1   g592(.A1(new_n684), .A2(new_n763), .A3(new_n771), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n408), .B(new_n779), .C1(new_n725), .C2(new_n726), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  INV_X1    g595(.A(KEYINPUT43), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(new_n654), .B2(new_n546), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT111), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n785), .B(new_n782), .C1(new_n654), .C2(new_n546), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n524), .A2(new_n545), .A3(KEYINPUT112), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT112), .B1(new_n524), .B2(new_n545), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n654), .A2(new_n782), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n784), .A2(new_n786), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n673), .B1(new_n639), .B2(new_n641), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT113), .B1(new_n794), .B2(new_n763), .ZN(new_n795));
  INV_X1    g609(.A(new_n793), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n784), .A2(new_n786), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n789), .A2(new_n790), .ZN(new_n798));
  OAI211_X1 g612(.A(KEYINPUT44), .B(new_n796), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n800));
  INV_X1    g614(.A(new_n763), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n795), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n768), .A2(KEYINPUT45), .A3(new_n628), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT109), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n632), .B(KEYINPUT108), .C1(new_n806), .C2(new_n598), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT109), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n768), .A2(new_n808), .A3(KEYINPUT45), .A4(new_n628), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n620), .B(KEYINPUT12), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n618), .B1(new_n810), .B2(new_n617), .ZN(new_n811));
  OAI21_X1  g625(.A(G469), .B1(new_n764), .B2(new_n615), .ZN(new_n812));
  OAI22_X1  g626(.A1(new_n811), .A2(new_n812), .B1(new_n806), .B2(new_n598), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT108), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n805), .A2(new_n807), .A3(new_n809), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n599), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT46), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT110), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n816), .A2(KEYINPUT46), .A3(new_n817), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n625), .A2(new_n598), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n818), .A2(KEYINPUT110), .A3(new_n819), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n822), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n792), .B1(new_n791), .B2(new_n793), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n596), .A4(new_n696), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n803), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(KEYINPUT114), .B(G137), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n830), .B(new_n831), .ZN(G39));
  NOR3_X1   g646(.A1(new_n763), .A2(new_n721), .A3(new_n408), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n727), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n727), .A2(KEYINPUT115), .A3(new_n833), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n827), .A2(KEYINPUT47), .A3(new_n596), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT47), .B1(new_n827), .B2(new_n596), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(G140), .ZN(G42));
  NAND2_X1  g657(.A1(new_n668), .A2(new_n746), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n641), .A2(KEYINPUT106), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n754), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n846), .A2(new_n408), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  INV_X1    g662(.A(new_n591), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n791), .A2(new_n849), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n409), .B(new_n731), .C1(new_n702), .C2(new_n703), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n847), .A2(new_n848), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n791), .A2(new_n849), .A3(new_n731), .A4(new_n763), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n748), .A2(new_n673), .A3(new_n754), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n801), .A2(new_n408), .A3(new_n591), .A4(new_n740), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n712), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n720), .A2(new_n546), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n853), .A2(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n850), .A2(new_n408), .A3(new_n846), .A4(new_n851), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT50), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n852), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n827), .A2(new_n596), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT47), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n728), .A2(new_n729), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n597), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n839), .A3(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n850), .A2(new_n408), .A3(new_n846), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n870), .A2(new_n801), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n861), .A2(new_n862), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT51), .B1(new_n863), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n727), .A2(new_n407), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n853), .A2(new_n874), .A3(KEYINPUT121), .A4(KEYINPUT48), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n870), .A2(new_n489), .A3(new_n740), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n853), .A2(new_n874), .ZN(new_n877));
  XOR2_X1   g691(.A(KEYINPUT121), .B(KEYINPUT48), .Z(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n590), .B1(new_n856), .B2(new_n655), .ZN(new_n880));
  AND4_X1   g694(.A1(new_n875), .A2(new_n876), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n869), .A2(new_n871), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n852), .A2(new_n858), .A3(new_n860), .A4(KEYINPUT51), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n873), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n642), .B1(new_n657), .B2(new_n663), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n635), .A2(new_n678), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n748), .A2(new_n772), .A3(new_n673), .A4(new_n754), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n643), .A2(new_n588), .A3(new_n683), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n889), .A2(new_n687), .A3(new_n763), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n725), .B2(new_n726), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n780), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n758), .A2(new_n742), .ZN(new_n895));
  INV_X1    g709(.A(new_n725), .ZN(new_n896));
  AOI22_X1  g710(.A1(new_n896), .A2(new_n327), .B1(new_n733), .B2(new_n737), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n894), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n347), .B(new_n732), .C1(new_n657), .C2(new_n663), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n899), .A2(KEYINPUT117), .A3(new_n742), .A4(new_n758), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n893), .A2(new_n777), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT53), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT52), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n730), .B1(new_n626), .B2(new_n769), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n713), .A2(new_n906), .A3(new_n683), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n755), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n908), .A2(new_n712), .A3(KEYINPUT118), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT118), .B1(new_n908), .B2(new_n712), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n723), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n692), .A2(new_n761), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n904), .B(new_n905), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n905), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n692), .A2(new_n761), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT118), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n338), .A2(new_n344), .B1(G472), .B2(new_n708), .ZN(new_n917));
  AOI211_X1 g731(.A(new_n730), .B(new_n682), .C1(new_n626), .C2(new_n769), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n489), .A2(new_n918), .A3(new_n713), .A4(new_n714), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n908), .A2(new_n712), .A3(KEYINPUT118), .ZN(new_n921));
  AOI22_X1  g735(.A1(new_n920), .A2(new_n921), .B1(new_n347), .B2(new_n722), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n915), .A2(KEYINPUT52), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n914), .A2(new_n923), .A3(KEYINPUT119), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n902), .A2(new_n903), .A3(new_n913), .A4(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n914), .A2(new_n923), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT53), .B1(new_n926), .B2(new_n901), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n925), .A2(KEYINPUT54), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n903), .B1(new_n926), .B2(new_n901), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT54), .ZN(new_n930));
  INV_X1    g744(.A(new_n892), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n635), .A2(new_n678), .A3(new_n886), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n777), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n895), .A2(new_n897), .A3(new_n903), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n924), .A2(new_n933), .A3(new_n913), .A4(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n929), .A2(new_n930), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n928), .A2(new_n936), .ZN(new_n937));
  OAI22_X1  g751(.A1(new_n885), .A2(new_n937), .B1(G952), .B2(G953), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n867), .B(KEYINPUT49), .Z(new_n939));
  NOR4_X1   g753(.A1(new_n939), .A2(new_n410), .A3(new_n597), .A4(new_n654), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n408), .A3(new_n789), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n941), .A2(new_n712), .A3(new_n705), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT116), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n938), .A2(new_n943), .ZN(G75));
  OAI21_X1  g758(.A(new_n460), .B1(new_n464), .B2(new_n466), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(new_n418), .Z(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT55), .ZN(new_n947));
  INV_X1    g761(.A(G210), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n948), .B(new_n390), .C1(new_n929), .C2(new_n935), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n949), .B2(KEYINPUT56), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT56), .ZN(new_n951));
  INV_X1    g765(.A(new_n947), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n929), .A2(new_n935), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(G902), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n951), .B(new_n952), .C1(new_n954), .C2(new_n948), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n383), .A2(G952), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n950), .A2(new_n955), .A3(new_n957), .ZN(G51));
  XNOR2_X1  g772(.A(new_n599), .B(KEYINPUT57), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n929), .A2(new_n930), .A3(new_n935), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n930), .B1(new_n929), .B2(new_n935), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n616), .A2(new_n624), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n954), .A2(new_n816), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n956), .B1(new_n964), .B2(new_n965), .ZN(G54));
  INV_X1    g780(.A(KEYINPUT122), .ZN(new_n967));
  NAND2_X1  g781(.A1(KEYINPUT58), .A2(G475), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n390), .B(new_n968), .C1(new_n929), .C2(new_n935), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n967), .B1(new_n969), .B2(new_n542), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n956), .B1(new_n969), .B2(new_n542), .ZN(new_n971));
  INV_X1    g785(.A(new_n542), .ZN(new_n972));
  OAI211_X1 g786(.A(KEYINPUT122), .B(new_n972), .C1(new_n954), .C2(new_n968), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(G60));
  AND2_X1   g788(.A1(new_n646), .A2(new_n647), .ZN(new_n975));
  NAND2_X1  g789(.A1(G478), .A2(G902), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT59), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n975), .B(new_n977), .C1(new_n960), .C2(new_n961), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n957), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n975), .B1(new_n937), .B2(new_n977), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(G63));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g796(.A1(G217), .A2(G902), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT60), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n929), .B2(new_n935), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n671), .B(KEYINPUT123), .Z(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n957), .B1(new_n985), .B2(new_n389), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n982), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n929), .A2(new_n935), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n401), .B1(new_n991), .B2(new_n984), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n992), .A2(KEYINPUT61), .A3(new_n957), .A4(new_n987), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n990), .A2(new_n993), .ZN(G66));
  OAI21_X1  g808(.A(G953), .B1(new_n593), .B2(new_n416), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n898), .A2(new_n932), .A3(new_n900), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n995), .B1(new_n996), .B2(G953), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n945), .B1(G898), .B2(new_n383), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(G69));
  AOI21_X1  g813(.A(new_n383), .B1(G227), .B2(G900), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n271), .A2(new_n272), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n315), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT124), .Z(new_n1003));
  NOR2_X1   g817(.A1(new_n530), .A2(new_n531), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n716), .A2(new_n692), .A3(new_n723), .A4(new_n761), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT62), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n842), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n697), .A2(new_n763), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n874), .B(new_n1011), .C1(new_n655), .C2(new_n662), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1012), .B1(new_n803), .B2(new_n829), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(KEYINPUT125), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT125), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n1015), .B(new_n1012), .C1(new_n803), .C2(new_n829), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1010), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1005), .B1(new_n1018), .B2(new_n383), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n912), .B1(new_n347), .B2(new_n722), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n727), .A2(new_n407), .A3(new_n755), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1021), .A2(new_n596), .A3(new_n696), .A4(new_n827), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1020), .A2(new_n1022), .A3(new_n777), .A4(new_n780), .ZN(new_n1023));
  AOI22_X1  g837(.A1(new_n866), .A2(new_n839), .B1(new_n836), .B2(new_n837), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n1023), .A2(new_n830), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n383), .ZN(new_n1026));
  NAND2_X1  g840(.A1(G900), .A2(G953), .ZN(new_n1027));
  AND3_X1   g841(.A1(new_n1026), .A2(new_n1005), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1000), .B1(new_n1019), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1026), .A2(new_n1005), .A3(new_n1027), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1000), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1017), .A2(G953), .ZN(new_n1032));
  OAI211_X1 g846(.A(new_n1030), .B(new_n1031), .C1(new_n1032), .C2(new_n1005), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1029), .A2(new_n1033), .ZN(G72));
  INV_X1    g848(.A(new_n316), .ZN(new_n1035));
  OR2_X1    g849(.A1(new_n1035), .A2(new_n192), .ZN(new_n1036));
  NAND2_X1  g850(.A1(G472), .A2(G902), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT63), .Z(new_n1038));
  NAND2_X1  g852(.A1(new_n1035), .A2(new_n192), .ZN(new_n1039));
  AND3_X1   g853(.A1(new_n1036), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n925), .A2(new_n927), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g855(.A(new_n1038), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1042), .B1(new_n1017), .B2(new_n996), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1041), .B1(new_n1043), .B2(new_n1039), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1042), .B1(new_n1025), .B2(new_n996), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n957), .B1(new_n1045), .B2(new_n1036), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT126), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g862(.A(KEYINPUT126), .B(new_n957), .C1(new_n1045), .C2(new_n1036), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1044), .B1(new_n1048), .B2(new_n1049), .ZN(G57));
endmodule


