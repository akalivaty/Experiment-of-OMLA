//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n550, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n617, new_n619,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  OR2_X1    g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT69), .Z(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(G2106), .B2(new_n454), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(KEYINPUT71), .A3(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G125), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT70), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G125), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n472), .B1(new_n481), .B2(G2105), .ZN(G160));
  INV_X1    g057(.A(new_n470), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n466), .A2(new_n468), .A3(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND4_X1  g065(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n469), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n467), .A2(new_n462), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(new_n473), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n491), .A2(KEYINPUT4), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n466), .A2(new_n468), .A3(G126), .A4(G2105), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n496), .A2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT72), .B1(new_n502), .B2(KEYINPUT6), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(new_n505), .A3(G651), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n503), .A2(new_n506), .B1(KEYINPUT6), .B2(new_n502), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G88), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n503), .A2(new_n506), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(G543), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G62), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n512), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n515), .A2(new_n520), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND2_X1  g101(.A1(new_n514), .A2(G89), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n519), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT7), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI211_X1 g108(.A(new_n531), .B(new_n532), .C1(new_n513), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n527), .A2(new_n528), .A3(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n502), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n514), .A2(G90), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n519), .A2(G52), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n502), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n514), .A2(G81), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n519), .A2(G43), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n518), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n507), .A2(KEYINPUT73), .A3(G53), .A4(G543), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n557), .A2(KEYINPUT9), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n512), .A2(KEYINPUT74), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n509), .B2(new_n511), .ZN(new_n562));
  XOR2_X1   g137(.A(KEYINPUT75), .B(G65), .Z(new_n563));
  NOR3_X1   g138(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AND2_X1   g139(.A1(G78), .A2(G543), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n555), .B(new_n567), .C1(new_n518), .C2(new_n556), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n514), .A2(G91), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n559), .A2(new_n566), .A3(new_n568), .A4(new_n569), .ZN(G299));
  NAND2_X1  g145(.A1(G168), .A2(KEYINPUT76), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT76), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n535), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(G286));
  NAND2_X1  g149(.A1(new_n514), .A2(G87), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n519), .A2(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n512), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n519), .A2(G48), .B1(G651), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n514), .A2(new_n583), .A3(G86), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n507), .A2(new_n513), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT77), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n582), .A2(new_n584), .A3(new_n587), .ZN(G305));
  XNOR2_X1  g163(.A(KEYINPUT78), .B(G47), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n519), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  XOR2_X1   g166(.A(KEYINPUT79), .B(G85), .Z(new_n592));
  OAI221_X1 g167(.A(new_n590), .B1(new_n502), .B2(new_n591), .C1(new_n585), .C2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n514), .A2(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n560), .A2(new_n562), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n519), .A2(G54), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n597), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT80), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n594), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n594), .B1(new_n606), .B2(G868), .ZN(G321));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n609));
  INV_X1    g184(.A(G286), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n611), .B2(G299), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n612), .B1(new_n614), .B2(new_n609), .ZN(G297));
  OAI21_X1  g190(.A(new_n612), .B1(new_n614), .B2(new_n609), .ZN(G280));
  NOR2_X1   g191(.A1(new_n605), .A2(G559), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(G860), .B2(new_n606), .ZN(G148));
  NAND2_X1  g193(.A1(new_n547), .A2(new_n611), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n617), .B2(new_n611), .ZN(G323));
  XOR2_X1   g195(.A(KEYINPUT82), .B(KEYINPUT11), .Z(new_n621));
  XNOR2_X1  g196(.A(G323), .B(new_n621), .ZN(G282));
  NAND2_X1  g197(.A1(new_n483), .A2(G135), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n485), .A2(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n469), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n493), .A2(new_n463), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT83), .B(G2100), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n630), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n628), .A2(new_n633), .ZN(G156));
  XOR2_X1   g209(.A(KEYINPUT84), .B(KEYINPUT14), .Z(new_n635));
  XOR2_X1   g210(.A(KEYINPUT15), .B(G2435), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2438), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2430), .Z(new_n638));
  AOI21_X1  g213(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n637), .B2(new_n638), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT16), .B(G1341), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  AND2_X1   g221(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(G14), .B1(new_n640), .B2(new_n646), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2072), .B(G2078), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT18), .Z(new_n654));
  XOR2_X1   g229(.A(new_n652), .B(KEYINPUT85), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(new_n650), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n650), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n651), .B(KEYINPUT17), .Z(new_n658));
  OAI21_X1  g233(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR3_X1   g234(.A1(new_n655), .A2(new_n651), .A3(new_n650), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n654), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2096), .B(G2100), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G227));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n666), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n666), .A2(new_n671), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n670), .B(new_n672), .C1(new_n673), .C2(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n673), .B2(new_n675), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1991), .ZN(new_n678));
  INV_X1    g253(.A(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(G229));
  MUX2_X1   g261(.A(G6), .B(G305), .S(G16), .Z(new_n687));
  XOR2_X1   g262(.A(KEYINPUT32), .B(G1981), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G22), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G166), .B2(new_n690), .ZN(new_n692));
  INV_X1    g267(.A(G1971), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n690), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT33), .B(G1976), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT88), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n697), .B(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n689), .A2(new_n694), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT34), .Z(new_n702));
  INV_X1    g277(.A(KEYINPUT36), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(KEYINPUT89), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G25), .ZN(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n707));
  INV_X1    g282(.A(G107), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G2105), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT87), .Z(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G131), .B2(new_n483), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n485), .A2(G119), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n706), .B1(new_n714), .B2(new_n705), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT35), .B(G1991), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  MUX2_X1   g292(.A(G24), .B(G290), .S(G16), .Z(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(G1986), .Z(new_n719));
  NAND4_X1  g294(.A1(new_n702), .A2(new_n704), .A3(new_n717), .A4(new_n719), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n703), .A2(KEYINPUT89), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n463), .A2(G103), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT91), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT25), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(new_n469), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G139), .B2(new_n483), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT92), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(KEYINPUT92), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n705), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n705), .B2(G33), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G2072), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n483), .A2(G141), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n485), .A2(G129), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n463), .A2(G105), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT26), .Z(new_n740));
  NAND4_X1  g315(.A1(new_n736), .A2(new_n737), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(new_n705), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n742), .A2(KEYINPUT93), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(KEYINPUT93), .ZN(new_n744));
  OAI22_X1  g319(.A1(new_n743), .A2(new_n744), .B1(G29), .B2(G32), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT27), .B(G1996), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(G171), .A2(G16), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G5), .B2(G16), .ZN(new_n749));
  INV_X1    g324(.A(G1961), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT24), .ZN(new_n752));
  INV_X1    g327(.A(G34), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n752), .B2(new_n753), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G160), .B2(new_n705), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n751), .B1(G2084), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n749), .A2(new_n750), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n548), .A2(G16), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G16), .B2(G19), .ZN(new_n760));
  INV_X1    g335(.A(G1341), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n757), .A2(new_n758), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(G168), .A2(G16), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G16), .B2(G21), .ZN(new_n765));
  INV_X1    g340(.A(G1966), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT94), .Z(new_n768));
  NAND4_X1  g343(.A1(new_n735), .A2(new_n747), .A3(new_n763), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G4), .A2(G16), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n606), .B2(G16), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1348), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n705), .A2(G35), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G162), .B2(new_n705), .ZN(new_n774));
  MUX2_X1   g349(.A(new_n773), .B(new_n774), .S(KEYINPUT96), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT29), .ZN(new_n776));
  INV_X1    g351(.A(G2090), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n705), .A2(G26), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n485), .A2(G128), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT90), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n483), .A2(G140), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n469), .A2(G116), .ZN(new_n784));
  OAI21_X1  g359(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n782), .B(new_n783), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n780), .A2(new_n781), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n779), .B1(new_n788), .B2(new_n705), .ZN(new_n789));
  MUX2_X1   g364(.A(new_n779), .B(new_n789), .S(KEYINPUT28), .Z(new_n790));
  INV_X1    g365(.A(G2067), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT30), .B(G28), .ZN(new_n793));
  OR2_X1    g368(.A1(KEYINPUT31), .A2(G11), .ZN(new_n794));
  NAND2_X1  g369(.A1(KEYINPUT31), .A2(G11), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n793), .A2(new_n705), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n627), .B2(new_n705), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n705), .A2(G27), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G164), .B2(new_n705), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT95), .B(G2078), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n756), .A2(G2084), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n801), .B(new_n802), .C1(new_n765), .C2(new_n766), .ZN(new_n803));
  AOI211_X1 g378(.A(new_n797), .B(new_n803), .C1(new_n761), .C2(new_n760), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n778), .A2(new_n792), .A3(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n769), .A2(new_n772), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT23), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n690), .A2(G20), .ZN(new_n808));
  AOI211_X1 g383(.A(new_n807), .B(new_n808), .C1(G299), .C2(G16), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n807), .B2(new_n808), .ZN(new_n810));
  INV_X1    g385(.A(G1956), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n722), .A2(new_n723), .A3(new_n806), .A4(new_n812), .ZN(G150));
  INV_X1    g388(.A(G150), .ZN(G311));
  NAND2_X1  g389(.A1(new_n606), .A2(G559), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT38), .Z(new_n816));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  INV_X1    g392(.A(G67), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n512), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G651), .ZN(new_n820));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  INV_X1    g396(.A(G93), .ZN(new_n822));
  OAI221_X1 g397(.A(new_n820), .B1(new_n518), .B2(new_n821), .C1(new_n822), .C2(new_n585), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT97), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(new_n547), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n548), .A2(new_n823), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT39), .Z(new_n829));
  AOI21_X1  g404(.A(G860), .B1(new_n816), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n816), .B2(new_n829), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT98), .Z(new_n832));
  INV_X1    g407(.A(new_n825), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G860), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT37), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n832), .A2(new_n835), .ZN(G145));
  NAND2_X1  g411(.A1(new_n483), .A2(G142), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n485), .A2(G130), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n469), .A2(G118), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n837), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n630), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n500), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n845));
  AOI221_X4 g420(.A(new_n845), .B1(new_n493), .B2(new_n495), .C1(new_n491), .C2(KEYINPUT4), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n493), .A2(new_n495), .ZN(new_n848));
  AOI21_X1  g423(.A(KEYINPUT100), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n844), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT101), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT101), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n852), .B(new_n844), .C1(new_n846), .C2(new_n849), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n788), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n854), .A2(new_n788), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n741), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n847), .A2(new_n848), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n845), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n496), .A2(KEYINPUT100), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n852), .B1(new_n862), .B2(new_n844), .ZN(new_n863));
  INV_X1    g438(.A(new_n853), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n788), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n741), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n855), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n858), .A2(KEYINPUT102), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n730), .B1(new_n870), .B2(KEYINPUT92), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n858), .A2(new_n869), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n732), .A2(KEYINPUT102), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n713), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n875), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n877), .A2(new_n871), .A3(new_n714), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n843), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n872), .A2(new_n875), .A3(new_n713), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n714), .B1(new_n877), .B2(new_n871), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(new_n842), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n489), .B(KEYINPUT99), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(G160), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(new_n627), .Z(new_n886));
  AOI21_X1  g461(.A(G37), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n888));
  INV_X1    g463(.A(new_n886), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n879), .A2(new_n888), .A3(new_n889), .A4(new_n882), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n879), .A2(new_n889), .A3(new_n882), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT103), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT40), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n887), .A2(new_n892), .A3(new_n895), .A4(new_n890), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(G395));
  XOR2_X1   g472(.A(new_n617), .B(new_n828), .Z(new_n898));
  XNOR2_X1  g473(.A(new_n604), .B(G299), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT41), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n899), .A2(KEYINPUT41), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n898), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n900), .B1(KEYINPUT104), .B2(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n906), .A2(KEYINPUT104), .ZN(new_n908));
  XNOR2_X1  g483(.A(G166), .B(G290), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n696), .B(G305), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n911), .B(KEYINPUT42), .Z(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n907), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n907), .B2(new_n908), .ZN(new_n915));
  OAI21_X1  g490(.A(G868), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(G868), .B2(new_n825), .ZN(G295));
  OAI21_X1  g492(.A(new_n916), .B1(G868), .B2(new_n825), .ZN(G331));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  NOR2_X1   g494(.A1(G171), .A2(new_n535), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n920), .B1(G286), .B2(G171), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n828), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n828), .A2(new_n921), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n901), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n911), .A2(KEYINPUT105), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n899), .B(new_n902), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n925), .B(new_n926), .C1(new_n927), .C2(new_n924), .ZN(new_n928));
  INV_X1    g503(.A(G37), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n899), .B1(new_n922), .B2(new_n923), .ZN(new_n931));
  INV_X1    g506(.A(new_n924), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n932), .B2(new_n905), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n933), .A2(new_n926), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n919), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n899), .A2(KEYINPUT107), .A3(KEYINPUT41), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n936), .A2(new_n922), .A3(new_n923), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n903), .A2(new_n938), .A3(new_n904), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n931), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT108), .B1(new_n940), .B2(new_n911), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  INV_X1    g517(.A(new_n911), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n936), .A2(new_n922), .A3(new_n923), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n944), .B1(new_n927), .B2(new_n938), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n942), .B(new_n943), .C1(new_n945), .C2(new_n931), .ZN(new_n946));
  AOI21_X1  g521(.A(G37), .B1(new_n933), .B2(new_n911), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n941), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n935), .B1(new_n948), .B2(new_n919), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT44), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT43), .B1(new_n930), .B2(new_n934), .ZN(new_n951));
  OAI211_X1 g526(.A(KEYINPUT106), .B(new_n951), .C1(new_n948), .C2(KEYINPUT43), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n951), .A2(KEYINPUT106), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n950), .B1(new_n954), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g530(.A(G8), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n957));
  AOI211_X1 g532(.A(new_n957), .B(G1384), .C1(new_n851), .C2(new_n853), .ZN(new_n958));
  INV_X1    g533(.A(G40), .ZN(new_n959));
  AOI211_X1 g534(.A(new_n959), .B(new_n472), .C1(new_n481), .C2(G2105), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n496), .B2(new_n500), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n957), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n693), .B1(new_n958), .B2(new_n964), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n962), .A2(KEYINPUT50), .ZN(new_n966));
  AOI21_X1  g541(.A(G1384), .B1(new_n862), .B2(new_n844), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n960), .B(new_n966), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n969), .A2(G2090), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n956), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(G303), .A2(G8), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT55), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT112), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n956), .B1(new_n967), .B2(new_n960), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n696), .A2(G1976), .ZN(new_n977));
  INV_X1    g552(.A(G1976), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT52), .B1(G288), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n960), .A2(new_n850), .A3(new_n961), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n981), .A3(G8), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT52), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT49), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n581), .A2(G651), .ZN(new_n986));
  INV_X1    g561(.A(G48), .ZN(new_n987));
  XNOR2_X1  g562(.A(KEYINPUT110), .B(G86), .ZN(new_n988));
  OAI221_X1 g563(.A(new_n986), .B1(new_n518), .B2(new_n987), .C1(new_n585), .C2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(G1981), .ZN(new_n990));
  INV_X1    g565(.A(G1981), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n582), .A2(new_n584), .A3(new_n991), .A4(new_n587), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n985), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n976), .B1(new_n984), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n993), .A2(new_n984), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n980), .B(new_n983), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G125), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n492), .B2(new_n473), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n480), .B1(new_n998), .B2(new_n478), .ZN(new_n999));
  INV_X1    g574(.A(new_n479), .ZN(new_n1000));
  OAI21_X1  g575(.A(G2105), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n472), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(G40), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n962), .A2(KEYINPUT50), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n850), .A2(new_n968), .A3(new_n961), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n962), .A2(KEYINPUT109), .A3(KEYINPUT50), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1009), .A2(G2090), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n956), .B1(new_n965), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n996), .B1(new_n1011), .B2(new_n974), .ZN(new_n1012));
  OAI211_X1 g587(.A(KEYINPUT45), .B(new_n961), .C1(new_n863), .C2(new_n864), .ZN(new_n1013));
  INV_X1    g588(.A(new_n964), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1971), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n969), .A2(G2090), .ZN(new_n1016));
  OAI21_X1  g591(.A(G8), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n973), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n967), .A2(KEYINPUT45), .ZN(new_n1021));
  OAI211_X1 g596(.A(G160), .B(G40), .C1(new_n962), .C2(new_n957), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1020), .B(new_n766), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n850), .A2(new_n961), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1022), .B1(new_n1024), .B2(new_n957), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT113), .B1(new_n1025), .B2(G1966), .ZN(new_n1026));
  INV_X1    g601(.A(G2084), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1006), .A2(new_n1007), .A3(new_n1027), .A4(new_n1008), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1023), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1029), .A2(G8), .A3(new_n610), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n975), .A2(new_n1012), .A3(new_n1019), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT63), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1009), .A2(G2090), .ZN(new_n1034));
  OAI21_X1  g609(.A(G8), .B1(new_n1015), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n973), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1012), .A2(KEYINPUT63), .A3(new_n1030), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1029), .A2(G8), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1040), .A2(new_n1032), .A3(G286), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1041), .A2(KEYINPUT114), .A3(new_n1012), .A4(new_n1036), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1033), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1035), .A2(new_n996), .A3(new_n973), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n978), .B(new_n696), .C1(new_n994), .C2(new_n995), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n992), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1044), .B1(new_n976), .B2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT56), .B(G2072), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1013), .A2(new_n1014), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n969), .A2(new_n811), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1052), .A2(KEYINPUT115), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(KEYINPUT115), .ZN(new_n1054));
  XOR2_X1   g629(.A(new_n1054), .B(KEYINPUT116), .Z(new_n1055));
  AND3_X1   g630(.A1(G299), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1055), .B1(G299), .B2(new_n1053), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT117), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OR3_X1    g633(.A1(new_n1056), .A2(new_n1057), .A3(KEYINPUT117), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1051), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AND4_X1   g635(.A1(new_n961), .A2(new_n960), .A3(new_n850), .A4(new_n791), .ZN(new_n1061));
  INV_X1    g636(.A(G1348), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1061), .B1(new_n1009), .B2(new_n1062), .ZN(new_n1063));
  OR2_X1    g638(.A1(new_n1063), .A2(new_n604), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1049), .A2(new_n1050), .A3(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1066), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1051), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1049), .A2(new_n1066), .A3(new_n1050), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT61), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT120), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1063), .A2(KEYINPUT60), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1009), .A2(new_n1062), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1061), .ZN(new_n1077));
  AND4_X1   g652(.A1(KEYINPUT60), .A2(new_n1076), .A3(new_n604), .A4(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n604), .B1(new_n1063), .B2(KEYINPUT60), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1075), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n547), .B1(KEYINPUT119), .B2(KEYINPUT59), .ZN(new_n1081));
  AOI21_X1  g656(.A(G1384), .B1(new_n851), .B2(new_n853), .ZN(new_n1082));
  AOI211_X1 g657(.A(G1996), .B(new_n964), .C1(new_n1082), .C2(KEYINPUT45), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT58), .B(G1341), .Z(new_n1084));
  NAND2_X1  g659(.A1(new_n981), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT118), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n981), .A2(new_n1087), .A3(new_n1084), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1081), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI221_X1 g667(.A(new_n1081), .B1(KEYINPUT119), .B2(KEYINPUT59), .C1(new_n1083), .C2(new_n1089), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1080), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1074), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1071), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1049), .A2(new_n1066), .A3(new_n1050), .A4(KEYINPUT121), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1097), .A2(new_n1060), .A3(KEYINPUT61), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1066), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1100));
  OAI211_X1 g675(.A(KEYINPUT120), .B(new_n1073), .C1(new_n1067), .C2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1068), .B1(new_n1095), .B2(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n975), .A2(new_n1012), .A3(new_n1019), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n535), .A2(G8), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1029), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n1106), .B2(KEYINPUT122), .ZN(new_n1110));
  OAI211_X1 g685(.A(G8), .B(new_n1110), .C1(new_n1029), .C2(new_n535), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI211_X1 g687(.A(new_n1107), .B(new_n1110), .C1(new_n1029), .C2(G8), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1108), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(G301), .B(KEYINPUT54), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1082), .A2(KEYINPUT45), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n1117));
  NOR4_X1   g692(.A1(new_n1116), .A2(new_n1117), .A3(G2078), .A4(new_n1003), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1115), .B1(new_n1118), .B2(new_n1013), .ZN(new_n1119));
  INV_X1    g694(.A(G2078), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1013), .A2(new_n1120), .A3(new_n1014), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1121), .A2(new_n1117), .B1(new_n750), .B2(new_n1009), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1025), .A2(KEYINPUT53), .A3(new_n1120), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1119), .A2(new_n1122), .B1(new_n1124), .B2(new_n1115), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1105), .A2(new_n1114), .A3(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1043), .B(new_n1047), .C1(new_n1104), .C2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT123), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1073), .B1(new_n1067), .B2(new_n1100), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1131), .A2(new_n1080), .A3(new_n1093), .A4(new_n1092), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1132), .A2(new_n1102), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1105), .A2(new_n1114), .A3(new_n1125), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1135), .A2(new_n1136), .A3(new_n1043), .A4(new_n1047), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1138), .B(new_n1108), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1139));
  AOI21_X1  g714(.A(G301), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(new_n1105), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT124), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1139), .A2(new_n1105), .A3(new_n1143), .A4(new_n1140), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1114), .A2(KEYINPUT62), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1142), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1128), .A2(new_n1137), .A3(new_n1146), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1082), .A2(KEYINPUT45), .A3(new_n1003), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n714), .A2(new_n716), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n788), .B(G2067), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n741), .B(new_n679), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n714), .A2(new_n716), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(G290), .B(G1986), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1148), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1147), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1148), .A2(new_n679), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT46), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1150), .A2(new_n868), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1157), .A2(new_n1158), .B1(new_n1148), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n1158), .B2(new_n1157), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT47), .ZN(new_n1162));
  XOR2_X1   g737(.A(new_n1152), .B(KEYINPUT125), .Z(new_n1163));
  NAND2_X1  g738(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1163), .A2(new_n1164), .B1(G2067), .B2(new_n866), .ZN(new_n1165));
  NOR2_X1   g740(.A1(G290), .A2(G1986), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1148), .A2(KEYINPUT48), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT48), .B1(new_n1148), .B2(new_n1166), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1168), .B1(new_n1148), .B2(new_n1153), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1165), .A2(new_n1148), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1162), .A2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT126), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1156), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g748(.A1(new_n663), .A2(G319), .ZN(new_n1175));
  XNOR2_X1  g749(.A(new_n1175), .B(KEYINPUT127), .ZN(new_n1176));
  OAI21_X1  g750(.A(new_n1176), .B1(new_n647), .B2(new_n648), .ZN(new_n1177));
  NOR3_X1   g751(.A1(new_n684), .A2(new_n685), .A3(new_n1177), .ZN(new_n1178));
  AND3_X1   g752(.A1(new_n952), .A2(new_n953), .A3(new_n1178), .ZN(new_n1179));
  AND2_X1   g753(.A1(new_n1179), .A2(new_n893), .ZN(G308));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n893), .ZN(G225));
endmodule


