

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U553 ( .A(n691), .ZN(n674) );
  NOR2_X2 U554 ( .A1(n679), .A2(n678), .ZN(n681) );
  AND2_X2 U555 ( .A1(n526), .A2(G2104), .ZN(n852) );
  NOR2_X2 U556 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  OR2_X1 U557 ( .A1(n659), .A2(n948), .ZN(n520) );
  OR2_X1 U558 ( .A1(n943), .A2(n660), .ZN(n521) );
  INV_X1 U559 ( .A(KEYINPUT26), .ZN(n644) );
  INV_X1 U560 ( .A(KEYINPUT94), .ZN(n680) );
  INV_X1 U561 ( .A(KEYINPUT32), .ZN(n699) );
  XNOR2_X1 U562 ( .A(n700), .B(n699), .ZN(n708) );
  INV_X1 U563 ( .A(KEYINPUT97), .ZN(n720) );
  OR2_X1 U564 ( .A1(n752), .A2(n596), .ZN(n628) );
  NAND2_X1 U565 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U566 ( .A(KEYINPUT0), .B(G543), .Z(n576) );
  NOR2_X2 U567 ( .A1(G2104), .A2(n526), .ZN(n848) );
  NOR2_X1 U568 ( .A1(G651), .A2(n576), .ZN(n787) );
  XOR2_X1 U569 ( .A(KEYINPUT1), .B(n535), .Z(n786) );
  BUF_X1 U570 ( .A(n589), .Z(G164) );
  INV_X1 U571 ( .A(G2105), .ZN(n526) );
  NAND2_X1 U572 ( .A1(G126), .A2(n848), .ZN(n523) );
  AND2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n849) );
  NAND2_X1 U574 ( .A1(G114), .A2(n849), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U576 ( .A(KEYINPUT84), .B(n524), .ZN(n530) );
  XOR2_X2 U577 ( .A(KEYINPUT17), .B(n525), .Z(n854) );
  NAND2_X1 U578 ( .A1(G138), .A2(n854), .ZN(n528) );
  NAND2_X1 U579 ( .A1(G102), .A2(n852), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U581 ( .A1(n530), .A2(n529), .ZN(n589) );
  XOR2_X1 U582 ( .A(KEYINPUT80), .B(KEYINPUT2), .Z(n533) );
  INV_X1 U583 ( .A(G651), .ZN(n534) );
  NOR2_X1 U584 ( .A1(n534), .A2(n576), .ZN(n531) );
  XNOR2_X2 U585 ( .A(n531), .B(KEYINPUT64), .ZN(n783) );
  NAND2_X1 U586 ( .A1(G73), .A2(n783), .ZN(n532) );
  XNOR2_X1 U587 ( .A(n533), .B(n532), .ZN(n540) );
  NOR2_X1 U588 ( .A1(G543), .A2(n534), .ZN(n535) );
  NAND2_X1 U589 ( .A1(G61), .A2(n786), .ZN(n537) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n782) );
  NAND2_X1 U591 ( .A1(G86), .A2(n782), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U593 ( .A(KEYINPUT79), .B(n538), .Z(n539) );
  NOR2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n787), .A2(G48), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n542), .A2(n541), .ZN(G305) );
  NAND2_X1 U597 ( .A1(G91), .A2(n782), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G53), .A2(n787), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U600 ( .A1(G65), .A2(n786), .ZN(n546) );
  NAND2_X1 U601 ( .A1(G78), .A2(n783), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U604 ( .A(n549), .B(KEYINPUT67), .ZN(G299) );
  NAND2_X1 U605 ( .A1(G77), .A2(n783), .ZN(n550) );
  XNOR2_X1 U606 ( .A(n550), .B(KEYINPUT66), .ZN(n552) );
  NAND2_X1 U607 ( .A1(G90), .A2(n782), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U609 ( .A(KEYINPUT9), .B(n553), .ZN(n557) );
  NAND2_X1 U610 ( .A1(G64), .A2(n786), .ZN(n555) );
  NAND2_X1 U611 ( .A1(G52), .A2(n787), .ZN(n554) );
  AND2_X1 U612 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n557), .A2(n556), .ZN(G301) );
  INV_X1 U614 ( .A(G301), .ZN(G171) );
  NAND2_X1 U615 ( .A1(n782), .A2(G89), .ZN(n558) );
  XNOR2_X1 U616 ( .A(KEYINPUT4), .B(n558), .ZN(n561) );
  NAND2_X1 U617 ( .A1(G76), .A2(n783), .ZN(n559) );
  XOR2_X1 U618 ( .A(KEYINPUT73), .B(n559), .Z(n560) );
  NAND2_X1 U619 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U620 ( .A(n562), .B(KEYINPUT5), .ZN(n567) );
  NAND2_X1 U621 ( .A1(G63), .A2(n786), .ZN(n564) );
  NAND2_X1 U622 ( .A1(G51), .A2(n787), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U624 ( .A(KEYINPUT6), .B(n565), .Z(n566) );
  NAND2_X1 U625 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U626 ( .A(n568), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(n782), .A2(G88), .ZN(n570) );
  NAND2_X1 U629 ( .A1(G75), .A2(n783), .ZN(n569) );
  NAND2_X1 U630 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U631 ( .A1(G62), .A2(n786), .ZN(n572) );
  NAND2_X1 U632 ( .A1(G50), .A2(n787), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U634 ( .A1(n574), .A2(n573), .ZN(G166) );
  XNOR2_X1 U635 ( .A(KEYINPUT85), .B(G166), .ZN(G303) );
  NAND2_X1 U636 ( .A1(G49), .A2(n787), .ZN(n575) );
  XNOR2_X1 U637 ( .A(n575), .B(KEYINPUT78), .ZN(n581) );
  NAND2_X1 U638 ( .A1(G87), .A2(n576), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G74), .A2(G651), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U641 ( .A1(n786), .A2(n579), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n581), .A2(n580), .ZN(G288) );
  NAND2_X1 U643 ( .A1(G72), .A2(n783), .ZN(n583) );
  NAND2_X1 U644 ( .A1(n786), .A2(G60), .ZN(n582) );
  NAND2_X1 U645 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U646 ( .A1(G85), .A2(n782), .ZN(n585) );
  NAND2_X1 U647 ( .A1(G47), .A2(n787), .ZN(n584) );
  NAND2_X1 U648 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U649 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U650 ( .A(KEYINPUT65), .B(n588), .ZN(G290) );
  NOR2_X2 U651 ( .A1(n589), .A2(G1384), .ZN(n629) );
  NAND2_X1 U652 ( .A1(n854), .A2(G137), .ZN(n592) );
  NAND2_X1 U653 ( .A1(G101), .A2(n852), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT23), .B(n590), .Z(n591) );
  NAND2_X1 U655 ( .A1(n592), .A2(n591), .ZN(n752) );
  NAND2_X1 U656 ( .A1(G125), .A2(n848), .ZN(n594) );
  NAND2_X1 U657 ( .A1(G113), .A2(n849), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n751) );
  INV_X1 U659 ( .A(G40), .ZN(n595) );
  OR2_X1 U660 ( .A1(n751), .A2(n595), .ZN(n596) );
  NOR2_X1 U661 ( .A1(n629), .A2(n628), .ZN(n746) );
  XNOR2_X1 U662 ( .A(KEYINPUT37), .B(G2067), .ZN(n744) );
  NAND2_X1 U663 ( .A1(G140), .A2(n854), .ZN(n598) );
  NAND2_X1 U664 ( .A1(G104), .A2(n852), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U666 ( .A(KEYINPUT34), .B(n599), .ZN(n604) );
  NAND2_X1 U667 ( .A1(G128), .A2(n848), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G116), .A2(n849), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U670 ( .A(KEYINPUT35), .B(n602), .Z(n603) );
  NOR2_X1 U671 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U672 ( .A(KEYINPUT36), .B(n605), .ZN(n862) );
  NOR2_X1 U673 ( .A1(n744), .A2(n862), .ZN(n1007) );
  NAND2_X1 U674 ( .A1(n746), .A2(n1007), .ZN(n742) );
  NAND2_X1 U675 ( .A1(G129), .A2(n848), .ZN(n607) );
  NAND2_X1 U676 ( .A1(G141), .A2(n854), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U678 ( .A1(G105), .A2(n852), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n608), .B(KEYINPUT89), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n609), .B(KEYINPUT38), .ZN(n610) );
  NOR2_X1 U681 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U682 ( .A1(n849), .A2(G117), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n613), .A2(n612), .ZN(n833) );
  NAND2_X1 U684 ( .A1(G1996), .A2(n833), .ZN(n614) );
  XOR2_X1 U685 ( .A(KEYINPUT90), .B(n614), .Z(n625) );
  NAND2_X1 U686 ( .A1(n852), .A2(G95), .ZN(n615) );
  XOR2_X1 U687 ( .A(KEYINPUT87), .B(n615), .Z(n617) );
  NAND2_X1 U688 ( .A1(n854), .A2(G131), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U690 ( .A(KEYINPUT88), .B(n618), .ZN(n621) );
  NAND2_X1 U691 ( .A1(n849), .A2(G107), .ZN(n619) );
  XOR2_X1 U692 ( .A(KEYINPUT86), .B(n619), .Z(n620) );
  NOR2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U694 ( .A1(n848), .A2(G119), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n845) );
  AND2_X1 U696 ( .A1(n845), .A2(G1991), .ZN(n624) );
  NOR2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n1005) );
  XNOR2_X1 U698 ( .A(KEYINPUT91), .B(n746), .ZN(n626) );
  NOR2_X1 U699 ( .A1(n1005), .A2(n626), .ZN(n739) );
  INV_X1 U700 ( .A(n739), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n742), .A2(n627), .ZN(n734) );
  INV_X1 U702 ( .A(n628), .ZN(n630) );
  NAND2_X2 U703 ( .A1(n630), .A2(n629), .ZN(n691) );
  NAND2_X1 U704 ( .A1(G8), .A2(n691), .ZN(n727) );
  NOR2_X1 U705 ( .A1(G1981), .A2(G305), .ZN(n631) );
  XOR2_X1 U706 ( .A(n631), .B(KEYINPUT24), .Z(n632) );
  NOR2_X1 U707 ( .A1(n727), .A2(n632), .ZN(n732) );
  NAND2_X1 U708 ( .A1(n787), .A2(G54), .ZN(n639) );
  NAND2_X1 U709 ( .A1(G66), .A2(n786), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G79), .A2(n783), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G92), .A2(n782), .ZN(n635) );
  XNOR2_X1 U713 ( .A(KEYINPUT71), .B(n635), .ZN(n636) );
  NOR2_X1 U714 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X2 U715 ( .A(KEYINPUT15), .B(n640), .Z(n943) );
  NAND2_X1 U716 ( .A1(G1348), .A2(n691), .ZN(n642) );
  NAND2_X1 U717 ( .A1(G2067), .A2(n674), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n642), .A2(n641), .ZN(n660) );
  INV_X1 U719 ( .A(G1996), .ZN(n643) );
  NOR2_X1 U720 ( .A1(n691), .A2(n643), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n645), .B(n644), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n691), .A2(G1341), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n659) );
  NAND2_X1 U724 ( .A1(G56), .A2(n786), .ZN(n648) );
  XNOR2_X1 U725 ( .A(KEYINPUT14), .B(n648), .ZN(n650) );
  NAND2_X1 U726 ( .A1(n787), .A2(G43), .ZN(n649) );
  AND2_X1 U727 ( .A1(n650), .A2(n649), .ZN(n658) );
  NAND2_X1 U728 ( .A1(G68), .A2(n783), .ZN(n651) );
  XNOR2_X1 U729 ( .A(KEYINPUT70), .B(n651), .ZN(n655) );
  XOR2_X1 U730 ( .A(KEYINPUT12), .B(KEYINPUT69), .Z(n653) );
  NAND2_X1 U731 ( .A1(G81), .A2(n782), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n653), .B(n652), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U734 ( .A(n656), .B(KEYINPUT13), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n658), .A2(n657), .ZN(n948) );
  NAND2_X1 U736 ( .A1(n521), .A2(n520), .ZN(n662) );
  NAND2_X1 U737 ( .A1(n943), .A2(n660), .ZN(n661) );
  NAND2_X1 U738 ( .A1(n662), .A2(n661), .ZN(n667) );
  INV_X1 U739 ( .A(G299), .ZN(n940) );
  NAND2_X1 U740 ( .A1(n674), .A2(G2072), .ZN(n663) );
  XNOR2_X1 U741 ( .A(n663), .B(KEYINPUT27), .ZN(n665) );
  INV_X1 U742 ( .A(G1956), .ZN(n972) );
  NOR2_X1 U743 ( .A1(n972), .A2(n674), .ZN(n664) );
  NOR2_X1 U744 ( .A1(n665), .A2(n664), .ZN(n668) );
  NAND2_X1 U745 ( .A1(n940), .A2(n668), .ZN(n666) );
  NAND2_X1 U746 ( .A1(n667), .A2(n666), .ZN(n672) );
  NOR2_X1 U747 ( .A1(n940), .A2(n668), .ZN(n670) );
  XNOR2_X1 U748 ( .A(KEYINPUT28), .B(KEYINPUT93), .ZN(n669) );
  XNOR2_X1 U749 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U750 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U751 ( .A(n673), .B(KEYINPUT29), .ZN(n679) );
  NAND2_X1 U752 ( .A1(n691), .A2(G1961), .ZN(n676) );
  XOR2_X1 U753 ( .A(G2078), .B(KEYINPUT25), .Z(n915) );
  NAND2_X1 U754 ( .A1(n674), .A2(n915), .ZN(n675) );
  NAND2_X1 U755 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U756 ( .A(n677), .B(KEYINPUT92), .Z(n682) );
  AND2_X1 U757 ( .A1(G171), .A2(n682), .ZN(n678) );
  XNOR2_X1 U758 ( .A(n681), .B(n680), .ZN(n690) );
  NOR2_X1 U759 ( .A1(G171), .A2(n682), .ZN(n687) );
  NOR2_X1 U760 ( .A1(G1966), .A2(n727), .ZN(n704) );
  NOR2_X1 U761 ( .A1(G2084), .A2(n691), .ZN(n701) );
  NOR2_X1 U762 ( .A1(n704), .A2(n701), .ZN(n683) );
  NAND2_X1 U763 ( .A1(G8), .A2(n683), .ZN(n684) );
  XNOR2_X1 U764 ( .A(KEYINPUT30), .B(n684), .ZN(n685) );
  NOR2_X1 U765 ( .A1(G168), .A2(n685), .ZN(n686) );
  NOR2_X1 U766 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U767 ( .A(KEYINPUT31), .B(n688), .Z(n689) );
  NAND2_X1 U768 ( .A1(n690), .A2(n689), .ZN(n702) );
  NAND2_X1 U769 ( .A1(n702), .A2(G286), .ZN(n698) );
  INV_X1 U770 ( .A(G8), .ZN(n696) );
  NOR2_X1 U771 ( .A1(G1971), .A2(n727), .ZN(n693) );
  NOR2_X1 U772 ( .A1(G2090), .A2(n691), .ZN(n692) );
  NOR2_X1 U773 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U774 ( .A1(n694), .A2(G303), .ZN(n695) );
  OR2_X1 U775 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U776 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U777 ( .A1(G8), .A2(n701), .ZN(n706) );
  INV_X1 U778 ( .A(n702), .ZN(n703) );
  NOR2_X1 U779 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U780 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U781 ( .A1(n708), .A2(n707), .ZN(n723) );
  NOR2_X1 U782 ( .A1(G1976), .A2(G288), .ZN(n716) );
  NOR2_X1 U783 ( .A1(G1971), .A2(G303), .ZN(n709) );
  NOR2_X1 U784 ( .A1(n716), .A2(n709), .ZN(n939) );
  NAND2_X1 U785 ( .A1(n723), .A2(n939), .ZN(n710) );
  XNOR2_X1 U786 ( .A(KEYINPUT95), .B(n710), .ZN(n713) );
  NAND2_X1 U787 ( .A1(G1976), .A2(G288), .ZN(n946) );
  INV_X1 U788 ( .A(n727), .ZN(n711) );
  NAND2_X1 U789 ( .A1(n946), .A2(n711), .ZN(n712) );
  NOR2_X1 U790 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U791 ( .A1(n714), .A2(KEYINPUT33), .ZN(n715) );
  XNOR2_X1 U792 ( .A(n715), .B(KEYINPUT96), .ZN(n719) );
  NAND2_X1 U793 ( .A1(n716), .A2(KEYINPUT33), .ZN(n717) );
  NOR2_X1 U794 ( .A1(n727), .A2(n717), .ZN(n718) );
  NOR2_X1 U795 ( .A1(n719), .A2(n718), .ZN(n721) );
  XNOR2_X1 U796 ( .A(n721), .B(n720), .ZN(n722) );
  XOR2_X1 U797 ( .A(G1981), .B(G305), .Z(n958) );
  NAND2_X1 U798 ( .A1(n722), .A2(n958), .ZN(n730) );
  NOR2_X1 U799 ( .A1(G2090), .A2(G303), .ZN(n724) );
  NAND2_X1 U800 ( .A1(G8), .A2(n724), .ZN(n725) );
  NAND2_X1 U801 ( .A1(n723), .A2(n725), .ZN(n726) );
  XNOR2_X1 U802 ( .A(n726), .B(KEYINPUT98), .ZN(n728) );
  NAND2_X1 U803 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U804 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U806 ( .A1(n734), .A2(n733), .ZN(n736) );
  XNOR2_X1 U807 ( .A(G1986), .B(G290), .ZN(n937) );
  NAND2_X1 U808 ( .A1(n937), .A2(n746), .ZN(n735) );
  NAND2_X1 U809 ( .A1(n736), .A2(n735), .ZN(n749) );
  NOR2_X1 U810 ( .A1(G1996), .A2(n833), .ZN(n1003) );
  NOR2_X1 U811 ( .A1(G1991), .A2(n845), .ZN(n1011) );
  NOR2_X1 U812 ( .A1(G1986), .A2(G290), .ZN(n737) );
  NOR2_X1 U813 ( .A1(n1011), .A2(n737), .ZN(n738) );
  NOR2_X1 U814 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U815 ( .A1(n1003), .A2(n740), .ZN(n741) );
  XNOR2_X1 U816 ( .A(n741), .B(KEYINPUT39), .ZN(n743) );
  NAND2_X1 U817 ( .A1(n743), .A2(n742), .ZN(n745) );
  NAND2_X1 U818 ( .A1(n744), .A2(n862), .ZN(n1015) );
  NAND2_X1 U819 ( .A1(n745), .A2(n1015), .ZN(n747) );
  NAND2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U822 ( .A(n750), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U823 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U824 ( .A(G57), .ZN(G237) );
  INV_X1 U825 ( .A(G120), .ZN(G236) );
  INV_X1 U826 ( .A(G132), .ZN(G219) );
  INV_X1 U827 ( .A(G82), .ZN(G220) );
  NOR2_X1 U828 ( .A1(n752), .A2(n751), .ZN(G160) );
  NAND2_X1 U829 ( .A1(G7), .A2(G661), .ZN(n753) );
  XNOR2_X1 U830 ( .A(n753), .B(KEYINPUT10), .ZN(n754) );
  XNOR2_X1 U831 ( .A(KEYINPUT68), .B(n754), .ZN(G223) );
  INV_X1 U832 ( .A(G223), .ZN(n819) );
  NAND2_X1 U833 ( .A1(n819), .A2(G567), .ZN(n755) );
  XOR2_X1 U834 ( .A(KEYINPUT11), .B(n755), .Z(G234) );
  INV_X1 U835 ( .A(G860), .ZN(n781) );
  OR2_X1 U836 ( .A1(n948), .A2(n781), .ZN(G153) );
  INV_X1 U837 ( .A(G868), .ZN(n759) );
  NAND2_X1 U838 ( .A1(n943), .A2(n759), .ZN(n756) );
  XNOR2_X1 U839 ( .A(n756), .B(KEYINPUT72), .ZN(n758) );
  NAND2_X1 U840 ( .A1(G868), .A2(G301), .ZN(n757) );
  NAND2_X1 U841 ( .A1(n758), .A2(n757), .ZN(G284) );
  NOR2_X1 U842 ( .A1(G286), .A2(n759), .ZN(n760) );
  XNOR2_X1 U843 ( .A(n760), .B(KEYINPUT74), .ZN(n762) );
  NOR2_X1 U844 ( .A1(G299), .A2(G868), .ZN(n761) );
  NOR2_X1 U845 ( .A1(n762), .A2(n761), .ZN(G297) );
  NAND2_X1 U846 ( .A1(n781), .A2(G559), .ZN(n763) );
  INV_X1 U847 ( .A(n943), .ZN(n779) );
  NAND2_X1 U848 ( .A1(n763), .A2(n779), .ZN(n764) );
  XNOR2_X1 U849 ( .A(n764), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U850 ( .A1(G868), .A2(n948), .ZN(n765) );
  XOR2_X1 U851 ( .A(KEYINPUT75), .B(n765), .Z(n768) );
  NAND2_X1 U852 ( .A1(G868), .A2(n779), .ZN(n766) );
  NOR2_X1 U853 ( .A1(G559), .A2(n766), .ZN(n767) );
  NOR2_X1 U854 ( .A1(n768), .A2(n767), .ZN(G282) );
  NAND2_X1 U855 ( .A1(n848), .A2(G123), .ZN(n769) );
  XNOR2_X1 U856 ( .A(n769), .B(KEYINPUT18), .ZN(n771) );
  NAND2_X1 U857 ( .A1(G135), .A2(n854), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U859 ( .A(KEYINPUT76), .B(n772), .ZN(n776) );
  NAND2_X1 U860 ( .A1(G111), .A2(n849), .ZN(n774) );
  NAND2_X1 U861 ( .A1(G99), .A2(n852), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n1010) );
  XNOR2_X1 U864 ( .A(n1010), .B(G2096), .ZN(n778) );
  INV_X1 U865 ( .A(G2100), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(G156) );
  NAND2_X1 U867 ( .A1(G559), .A2(n779), .ZN(n780) );
  XOR2_X1 U868 ( .A(n948), .B(n780), .Z(n800) );
  NAND2_X1 U869 ( .A1(n781), .A2(n800), .ZN(n793) );
  NAND2_X1 U870 ( .A1(n782), .A2(G93), .ZN(n785) );
  NAND2_X1 U871 ( .A1(G80), .A2(n783), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n792) );
  NAND2_X1 U873 ( .A1(G67), .A2(n786), .ZN(n789) );
  NAND2_X1 U874 ( .A1(G55), .A2(n787), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U876 ( .A(KEYINPUT77), .B(n790), .Z(n791) );
  NOR2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n802) );
  XOR2_X1 U878 ( .A(n793), .B(n802), .Z(G145) );
  XOR2_X1 U879 ( .A(KEYINPUT19), .B(KEYINPUT81), .Z(n794) );
  XNOR2_X1 U880 ( .A(G288), .B(n794), .ZN(n795) );
  XNOR2_X1 U881 ( .A(n802), .B(n795), .ZN(n797) );
  XNOR2_X1 U882 ( .A(G290), .B(G166), .ZN(n796) );
  XNOR2_X1 U883 ( .A(n797), .B(n796), .ZN(n798) );
  XNOR2_X1 U884 ( .A(n798), .B(G299), .ZN(n799) );
  XNOR2_X1 U885 ( .A(n799), .B(G305), .ZN(n868) );
  XNOR2_X1 U886 ( .A(n800), .B(n868), .ZN(n801) );
  NAND2_X1 U887 ( .A1(n801), .A2(G868), .ZN(n804) );
  OR2_X1 U888 ( .A1(G868), .A2(n802), .ZN(n803) );
  NAND2_X1 U889 ( .A1(n804), .A2(n803), .ZN(G295) );
  NAND2_X1 U890 ( .A1(G2084), .A2(G2078), .ZN(n805) );
  XOR2_X1 U891 ( .A(KEYINPUT20), .B(n805), .Z(n806) );
  NAND2_X1 U892 ( .A1(G2090), .A2(n806), .ZN(n807) );
  XNOR2_X1 U893 ( .A(KEYINPUT21), .B(n807), .ZN(n808) );
  NAND2_X1 U894 ( .A1(n808), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U895 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U896 ( .A1(G220), .A2(G219), .ZN(n809) );
  XOR2_X1 U897 ( .A(KEYINPUT22), .B(n809), .Z(n810) );
  NOR2_X1 U898 ( .A1(G218), .A2(n810), .ZN(n811) );
  NAND2_X1 U899 ( .A1(G96), .A2(n811), .ZN(n823) );
  NAND2_X1 U900 ( .A1(G2106), .A2(n823), .ZN(n812) );
  XNOR2_X1 U901 ( .A(n812), .B(KEYINPUT82), .ZN(n817) );
  NOR2_X1 U902 ( .A1(G236), .A2(G237), .ZN(n813) );
  NAND2_X1 U903 ( .A1(G69), .A2(n813), .ZN(n814) );
  XNOR2_X1 U904 ( .A(KEYINPUT83), .B(n814), .ZN(n815) );
  NAND2_X1 U905 ( .A1(n815), .A2(G108), .ZN(n824) );
  NAND2_X1 U906 ( .A1(G567), .A2(n824), .ZN(n816) );
  NAND2_X1 U907 ( .A1(n817), .A2(n816), .ZN(n893) );
  NAND2_X1 U908 ( .A1(G661), .A2(G483), .ZN(n818) );
  NOR2_X1 U909 ( .A1(n893), .A2(n818), .ZN(n822) );
  NAND2_X1 U910 ( .A1(n822), .A2(G36), .ZN(G176) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n819), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U913 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(G188) );
  INV_X1 U917 ( .A(G108), .ZN(G238) );
  INV_X1 U918 ( .A(G96), .ZN(G221) );
  NOR2_X1 U919 ( .A1(n824), .A2(n823), .ZN(G325) );
  INV_X1 U920 ( .A(G325), .ZN(G261) );
  NAND2_X1 U921 ( .A1(n848), .A2(G124), .ZN(n825) );
  XNOR2_X1 U922 ( .A(n825), .B(KEYINPUT44), .ZN(n827) );
  NAND2_X1 U923 ( .A1(G112), .A2(n849), .ZN(n826) );
  NAND2_X1 U924 ( .A1(n827), .A2(n826), .ZN(n831) );
  NAND2_X1 U925 ( .A1(G136), .A2(n854), .ZN(n829) );
  NAND2_X1 U926 ( .A1(G100), .A2(n852), .ZN(n828) );
  NAND2_X1 U927 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U928 ( .A1(n831), .A2(n830), .ZN(G162) );
  XOR2_X1 U929 ( .A(G160), .B(G162), .Z(n832) );
  XNOR2_X1 U930 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U931 ( .A(n834), .B(KEYINPUT48), .Z(n836) );
  XNOR2_X1 U932 ( .A(KEYINPUT106), .B(KEYINPUT46), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n844) );
  NAND2_X1 U934 ( .A1(G139), .A2(n854), .ZN(n838) );
  NAND2_X1 U935 ( .A1(G103), .A2(n852), .ZN(n837) );
  NAND2_X1 U936 ( .A1(n838), .A2(n837), .ZN(n843) );
  NAND2_X1 U937 ( .A1(G127), .A2(n848), .ZN(n840) );
  NAND2_X1 U938 ( .A1(G115), .A2(n849), .ZN(n839) );
  NAND2_X1 U939 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U940 ( .A(KEYINPUT47), .B(n841), .Z(n842) );
  NOR2_X1 U941 ( .A1(n843), .A2(n842), .ZN(n998) );
  XOR2_X1 U942 ( .A(n844), .B(n998), .Z(n847) );
  XOR2_X1 U943 ( .A(G164), .B(n845), .Z(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n864) );
  NAND2_X1 U945 ( .A1(G130), .A2(n848), .ZN(n851) );
  NAND2_X1 U946 ( .A1(G118), .A2(n849), .ZN(n850) );
  NAND2_X1 U947 ( .A1(n851), .A2(n850), .ZN(n859) );
  NAND2_X1 U948 ( .A1(n852), .A2(G106), .ZN(n853) );
  XOR2_X1 U949 ( .A(KEYINPUT105), .B(n853), .Z(n856) );
  NAND2_X1 U950 ( .A1(n854), .A2(G142), .ZN(n855) );
  NAND2_X1 U951 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U952 ( .A(KEYINPUT45), .B(n857), .Z(n858) );
  NOR2_X1 U953 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U954 ( .A(n1010), .B(n860), .Z(n861) );
  XNOR2_X1 U955 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U956 ( .A(n864), .B(n863), .Z(n865) );
  NOR2_X1 U957 ( .A1(G37), .A2(n865), .ZN(n866) );
  XOR2_X1 U958 ( .A(KEYINPUT107), .B(n866), .Z(G395) );
  XNOR2_X1 U959 ( .A(KEYINPUT108), .B(n948), .ZN(n867) );
  XNOR2_X1 U960 ( .A(n867), .B(n943), .ZN(n869) );
  XOR2_X1 U961 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U962 ( .A(G171), .B(G286), .ZN(n870) );
  XNOR2_X1 U963 ( .A(n871), .B(n870), .ZN(n872) );
  NOR2_X1 U964 ( .A1(G37), .A2(n872), .ZN(G397) );
  XOR2_X1 U965 ( .A(G2100), .B(KEYINPUT43), .Z(n874) );
  XNOR2_X1 U966 ( .A(KEYINPUT42), .B(G2678), .ZN(n873) );
  XNOR2_X1 U967 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U968 ( .A(KEYINPUT102), .B(G2090), .Z(n876) );
  XNOR2_X1 U969 ( .A(G2067), .B(G2072), .ZN(n875) );
  XNOR2_X1 U970 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U971 ( .A(n878), .B(n877), .Z(n880) );
  XNOR2_X1 U972 ( .A(KEYINPUT103), .B(G2096), .ZN(n879) );
  XNOR2_X1 U973 ( .A(n880), .B(n879), .ZN(n882) );
  XOR2_X1 U974 ( .A(G2084), .B(G2078), .Z(n881) );
  XNOR2_X1 U975 ( .A(n882), .B(n881), .ZN(G227) );
  XNOR2_X1 U976 ( .A(G1981), .B(G2474), .ZN(n892) );
  XOR2_X1 U977 ( .A(G1976), .B(G1971), .Z(n884) );
  XNOR2_X1 U978 ( .A(G1966), .B(G1961), .ZN(n883) );
  XNOR2_X1 U979 ( .A(n884), .B(n883), .ZN(n888) );
  XOR2_X1 U980 ( .A(G1956), .B(G1986), .Z(n886) );
  XNOR2_X1 U981 ( .A(G1996), .B(G1991), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U983 ( .A(n888), .B(n887), .Z(n890) );
  XNOR2_X1 U984 ( .A(KEYINPUT104), .B(KEYINPUT41), .ZN(n889) );
  XNOR2_X1 U985 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U986 ( .A(n892), .B(n891), .ZN(G229) );
  XNOR2_X1 U987 ( .A(KEYINPUT101), .B(n893), .ZN(G319) );
  NOR2_X1 U988 ( .A1(G395), .A2(G397), .ZN(n894) );
  XNOR2_X1 U989 ( .A(KEYINPUT110), .B(n894), .ZN(n911) );
  NOR2_X1 U990 ( .A1(G227), .A2(G229), .ZN(n895) );
  XNOR2_X1 U991 ( .A(n895), .B(KEYINPUT49), .ZN(n909) );
  XNOR2_X1 U992 ( .A(G2451), .B(G2446), .ZN(n905) );
  XOR2_X1 U993 ( .A(G2430), .B(G2443), .Z(n897) );
  XNOR2_X1 U994 ( .A(G2454), .B(G2435), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n901) );
  XOR2_X1 U996 ( .A(G2438), .B(KEYINPUT99), .Z(n899) );
  XNOR2_X1 U997 ( .A(G1341), .B(G1348), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U999 ( .A(n901), .B(n900), .Z(n903) );
  XNOR2_X1 U1000 ( .A(KEYINPUT100), .B(G2427), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(n906), .A2(G14), .ZN(n912) );
  NAND2_X1 U1004 ( .A1(n912), .A2(G319), .ZN(n907) );
  XOR2_X1 U1005 ( .A(KEYINPUT109), .B(n907), .Z(n908) );
  NOR2_X1 U1006 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G69), .ZN(G235) );
  INV_X1 U1010 ( .A(n912), .ZN(G401) );
  XOR2_X1 U1011 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n1029) );
  XNOR2_X1 U1012 ( .A(KEYINPUT113), .B(G2090), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n913), .B(G35), .ZN(n928) );
  XOR2_X1 U1014 ( .A(G25), .B(G1991), .Z(n914) );
  NAND2_X1 U1015 ( .A1(n914), .A2(G28), .ZN(n924) );
  XNOR2_X1 U1016 ( .A(G1996), .B(G32), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(n915), .B(G27), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(KEYINPUT114), .B(n918), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(G2067), .B(G26), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(G33), .B(G2072), .ZN(n919) );
  NOR2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(KEYINPUT53), .B(KEYINPUT115), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(n926), .B(n925), .ZN(n927) );
  NAND2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(G34), .B(G2084), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(KEYINPUT54), .B(n929), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(KEYINPUT55), .B(n932), .ZN(n934) );
  INV_X1 U1032 ( .A(G29), .ZN(n933) );
  NAND2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n935), .A2(G11), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(KEYINPUT116), .B(n936), .ZN(n996) );
  XNOR2_X1 U1036 ( .A(G16), .B(KEYINPUT56), .ZN(n963) );
  INV_X1 U1037 ( .A(n937), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n954) );
  XNOR2_X1 U1039 ( .A(G171), .B(G1961), .ZN(n952) );
  XNOR2_X1 U1040 ( .A(n940), .B(G1956), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(G1971), .A2(G303), .ZN(n941) );
  NAND2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(G1348), .B(n943), .ZN(n944) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n947) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G1341), .B(n948), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(KEYINPUT118), .B(n955), .ZN(n961) );
  XOR2_X1 U1051 ( .A(G1966), .B(G168), .Z(n956) );
  XNOR2_X1 U1052 ( .A(KEYINPUT117), .B(n956), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(KEYINPUT57), .B(n959), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n994) );
  INV_X1 U1057 ( .A(G16), .ZN(n992) );
  XNOR2_X1 U1058 ( .A(G1986), .B(G24), .ZN(n970) );
  XNOR2_X1 U1059 ( .A(G1976), .B(KEYINPUT122), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n964), .B(G23), .ZN(n967) );
  XOR2_X1 U1061 ( .A(G1971), .B(G22), .Z(n965) );
  XNOR2_X1 U1062 ( .A(KEYINPUT121), .B(n965), .ZN(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(KEYINPUT123), .B(n968), .ZN(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(KEYINPUT58), .B(n971), .ZN(n988) );
  XNOR2_X1 U1067 ( .A(G20), .B(n972), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(G1341), .B(G19), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(G6), .B(G1981), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1071 ( .A(KEYINPUT119), .B(n975), .Z(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n980) );
  XOR2_X1 U1073 ( .A(KEYINPUT59), .B(G1348), .Z(n978) );
  XNOR2_X1 U1074 ( .A(G4), .B(n978), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1076 ( .A(KEYINPUT60), .B(n981), .Z(n983) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G21), .ZN(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1079 ( .A(KEYINPUT120), .B(n984), .Z(n986) );
  XNOR2_X1 U1080 ( .A(G1961), .B(G5), .ZN(n985) );
  NOR2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(n989), .B(KEYINPUT61), .ZN(n990) );
  XOR2_X1 U1084 ( .A(KEYINPUT124), .B(n990), .Z(n991) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1088 ( .A(KEYINPUT125), .B(n997), .Z(n1027) );
  XOR2_X1 U1089 ( .A(G2072), .B(n998), .Z(n1000) );
  XOR2_X1 U1090 ( .A(G164), .B(G2078), .Z(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1092 ( .A(KEYINPUT50), .B(n1001), .Z(n1021) );
  XOR2_X1 U1093 ( .A(G2090), .B(G162), .Z(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1095 ( .A(KEYINPUT51), .B(n1004), .Z(n1009) );
  INV_X1 U1096 ( .A(n1005), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1018) );
  XNOR2_X1 U1099 ( .A(G160), .B(G2084), .ZN(n1013) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(n1014), .B(KEYINPUT111), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1105 ( .A(KEYINPUT112), .B(n1019), .Z(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(KEYINPUT52), .B(n1022), .ZN(n1024) );
  INV_X1 U1108 ( .A(KEYINPUT55), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(G29), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(n1029), .B(n1028), .ZN(G311) );
  XNOR2_X1 U1113 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

