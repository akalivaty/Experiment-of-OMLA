//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974;
  INV_X1    g000(.A(KEYINPUT103), .ZN(new_n202));
  INV_X1    g001(.A(G218gat), .ZN(new_n203));
  AND2_X1   g002(.A1(G43gat), .A2(G50gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G43gat), .A2(G50gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT91), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G43gat), .ZN(new_n207));
  INV_X1    g006(.A(G50gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT91), .ZN(new_n210));
  NAND2_X1  g009(.A1(G43gat), .A2(G50gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n206), .A2(new_n212), .A3(KEYINPUT15), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  INV_X1    g013(.A(G36gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT14), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT14), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G29gat), .B2(G36gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT92), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n219), .A2(KEYINPUT92), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n213), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT95), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT15), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n211), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(KEYINPUT91), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT94), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n219), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT94), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n212), .A2(new_n227), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n209), .A2(new_n225), .A3(new_n211), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT93), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n209), .A2(KEYINPUT93), .A3(new_n225), .A4(new_n211), .ZN(new_n235));
  NAND2_X1  g034(.A1(G29gat), .A2(G36gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n224), .B1(new_n231), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT94), .B1(new_n216), .B2(new_n218), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT94), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n213), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n242), .A2(KEYINPUT95), .A3(new_n237), .ZN(new_n243));
  OAI211_X1 g042(.A(KEYINPUT17), .B(new_n223), .C1(new_n239), .C2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT101), .B(G92gat), .ZN(new_n245));
  INV_X1    g044(.A(G85gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n245), .A2(new_n246), .B1(KEYINPUT8), .B2(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(G99gat), .A2(G106gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(G99gat), .A2(G106gat), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT102), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OR2_X1    g050(.A1(G99gat), .A2(G106gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT102), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n253), .A3(new_n247), .ZN(new_n254));
  NAND2_X1  g053(.A1(G85gat), .A2(G92gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT7), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT7), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(G85gat), .A3(G92gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n248), .A2(new_n251), .A3(new_n254), .A4(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G92gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT101), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT101), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G92gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n264), .A3(new_n246), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n247), .A2(KEYINPUT8), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n259), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n254), .A2(new_n251), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n260), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n231), .A2(new_n238), .A3(new_n224), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT95), .B1(new_n242), .B2(new_n237), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n222), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT96), .B(KEYINPUT17), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n244), .B(new_n271), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G190gat), .ZN(new_n277));
  AND3_X1   g076(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n223), .B1(new_n239), .B2(new_n243), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(new_n270), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n276), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n277), .B1(new_n276), .B2(new_n280), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n203), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n244), .A2(new_n271), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n274), .A2(new_n275), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n280), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G190gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n276), .A2(new_n277), .A3(new_n280), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n287), .A2(G218gat), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT100), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n283), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G134gat), .B(G162gat), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n292), .B(new_n293), .Z(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n283), .A2(new_n289), .A3(new_n290), .A4(new_n294), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G57gat), .B(G64gat), .Z(new_n299));
  INV_X1    g098(.A(G71gat), .ZN(new_n300));
  INV_X1    g099(.A(G78gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G71gat), .A2(G78gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT9), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n299), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G57gat), .B(G64gat), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n303), .B(new_n302), .C1(new_n308), .C2(new_n305), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT21), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G231gat), .A2(G233gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G127gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G15gat), .B(G22gat), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n317), .A2(G1gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT16), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n319), .B2(G1gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(KEYINPUT97), .ZN(new_n322));
  INV_X1    g121(.A(G8gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n318), .B(new_n320), .C1(KEYINPUT97), .C2(G8gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(new_n311), .B2(new_n310), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n316), .B(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n329));
  INV_X1    g128(.A(G155gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(G183gat), .B(G211gat), .Z(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n328), .B(new_n333), .Z(new_n334));
  OAI21_X1  g133(.A(new_n202), .B1(new_n298), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n328), .B(new_n333), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n336), .A2(new_n296), .A3(KEYINPUT103), .A4(new_n297), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n244), .B(new_n326), .C1(new_n274), .C2(new_n275), .ZN(new_n340));
  NAND2_X1  g139(.A1(G229gat), .A2(G233gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n272), .A2(new_n273), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n326), .B1(new_n342), .B2(new_n223), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n340), .A2(KEYINPUT18), .A3(new_n341), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT98), .ZN(new_n346));
  INV_X1    g145(.A(new_n326), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n347), .B1(new_n274), .B2(KEYINPUT17), .ZN(new_n348));
  INV_X1    g147(.A(new_n275), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n279), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n343), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT98), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT18), .A4(new_n341), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n346), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G113gat), .B(G141gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(G197gat), .ZN(new_n356));
  XOR2_X1   g155(.A(KEYINPUT11), .B(G169gat), .Z(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(KEYINPUT90), .B(KEYINPUT12), .Z(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n341), .B(KEYINPUT13), .Z(new_n362));
  AND3_X1   g161(.A1(new_n342), .A2(new_n223), .A3(new_n326), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n362), .B1(new_n363), .B2(new_n343), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT99), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT99), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n366), .B(new_n362), .C1(new_n363), .C2(new_n343), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n340), .A2(new_n341), .A3(new_n344), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT18), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n365), .A2(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n354), .A2(new_n361), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n361), .B1(new_n354), .B2(new_n370), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n307), .A2(new_n309), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n248), .A2(new_n259), .B1(new_n251), .B2(new_n254), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n267), .A2(new_n268), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n260), .A2(new_n310), .A3(new_n269), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n270), .A2(KEYINPUT10), .A3(new_n375), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G230gat), .A2(G233gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n384), .B(KEYINPUT104), .Z(new_n385));
  OAI21_X1  g184(.A(KEYINPUT105), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n385), .B1(new_n381), .B2(new_n382), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT105), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n385), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n378), .B2(new_n380), .ZN(new_n391));
  XNOR2_X1  g190(.A(G120gat), .B(G148gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G176gat), .B(G204gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n386), .A2(new_n389), .A3(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n395), .B1(new_n387), .B2(new_n391), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT106), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n339), .A2(new_n374), .A3(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(G227gat), .A2(G233gat), .ZN(new_n403));
  INV_X1    g202(.A(G113gat), .ZN(new_n404));
  INV_X1    g203(.A(G120gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT1), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(G113gat), .B2(G120gat), .ZN(new_n408));
  OAI211_X1 g207(.A(KEYINPUT73), .B(G134gat), .C1(new_n406), .C2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT1), .B1(new_n404), .B2(new_n405), .ZN(new_n410));
  INV_X1    g209(.A(G134gat), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n410), .B(new_n411), .C1(new_n404), .C2(new_n405), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n409), .A2(new_n412), .A3(new_n315), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n315), .B1(new_n409), .B2(new_n412), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G169gat), .A2(G176gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(G169gat), .A2(G176gat), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(KEYINPUT23), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n419), .B1(KEYINPUT23), .B2(new_n418), .ZN(new_n420));
  NAND2_X1  g219(.A1(G183gat), .A2(G190gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT24), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(new_n423), .B(KEYINPUT66), .Z(new_n424));
  OAI21_X1  g223(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n425));
  NAND3_X1  g224(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n420), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT25), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n419), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G169gat), .ZN(new_n432));
  INV_X1    g231(.A(G176gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT67), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT67), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(KEYINPUT23), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT68), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n421), .A2(new_n439), .A3(new_n422), .ZN(new_n440));
  INV_X1    g239(.A(G183gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(new_n277), .A3(KEYINPUT69), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT69), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(G183gat), .B2(G190gat), .ZN(new_n444));
  OAI211_X1 g243(.A(G183gat), .B(G190gat), .C1(KEYINPUT68), .C2(KEYINPUT24), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n440), .A2(new_n442), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n438), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT70), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n431), .A2(new_n438), .A3(KEYINPUT70), .A4(new_n446), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n428), .A2(new_n429), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT27), .ZN(new_n452));
  AOI21_X1  g251(.A(G190gat), .B1(new_n452), .B2(G183gat), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT28), .B1(new_n453), .B2(KEYINPUT71), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n441), .A2(KEYINPUT27), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n453), .B(new_n455), .C1(KEYINPUT71), .C2(KEYINPUT28), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT72), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT72), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n461), .A3(new_n458), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT26), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n435), .A2(new_n463), .A3(new_n437), .ZN(new_n464));
  INV_X1    g263(.A(new_n417), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n465), .B1(KEYINPUT26), .B2(new_n434), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n464), .A2(new_n466), .B1(G183gat), .B2(G190gat), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n460), .A2(new_n462), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n416), .B1(new_n451), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n428), .A2(new_n429), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n449), .A2(new_n450), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n460), .A2(new_n462), .A3(new_n467), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n415), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n403), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT34), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI211_X1 g276(.A(KEYINPUT34), .B(new_n403), .C1(new_n469), .C2(new_n474), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(G15gat), .B(G43gat), .Z(new_n480));
  XNOR2_X1  g279(.A(G71gat), .B(G99gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n469), .A2(new_n403), .A3(new_n474), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT33), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n479), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n484), .A2(KEYINPUT32), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n486), .B1(new_n477), .B2(new_n478), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n490), .B1(new_n488), .B2(new_n491), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT36), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT36), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(new_n493), .B2(new_n494), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT31), .B(G50gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G141gat), .B(G148gat), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G162gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n330), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G155gat), .A2(G162gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(KEYINPUT2), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n503), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n506), .B(new_n505), .C1(new_n502), .C2(KEYINPUT2), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G197gat), .B(G204gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT22), .ZN(new_n513));
  INV_X1    g312(.A(G211gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(new_n203), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G211gat), .B(G218gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(KEYINPUT29), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n511), .B1(new_n519), .B2(KEYINPUT3), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(KEYINPUT74), .ZN(new_n521));
  INV_X1    g320(.A(new_n517), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n516), .B(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT74), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XOR2_X1   g324(.A(KEYINPUT80), .B(KEYINPUT3), .Z(new_n526));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n510), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT29), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n521), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n520), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(G228gat), .A3(G233gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(KEYINPUT88), .ZN(new_n533));
  NAND2_X1  g332(.A1(G228gat), .A2(G233gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n521), .A2(new_n525), .A3(new_n535), .A4(new_n529), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n526), .B1(new_n518), .B2(KEYINPUT29), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n511), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n533), .A2(new_n534), .A3(new_n536), .A4(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n501), .B1(new_n532), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G78gat), .B(G106gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G22gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n532), .A2(new_n539), .A3(new_n501), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n543), .ZN(new_n546));
  INV_X1    g345(.A(new_n544), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(new_n540), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G8gat), .B(G36gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT78), .ZN(new_n551));
  XNOR2_X1  g350(.A(G64gat), .B(G92gat), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n551), .B(new_n552), .Z(new_n553));
  NAND2_X1  g352(.A1(G226gat), .A2(G233gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT75), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT76), .B1(new_n451), .B2(new_n468), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT76), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n472), .A2(new_n558), .A3(new_n473), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n556), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n521), .A2(new_n525), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AOI211_X1 g361(.A(KEYINPUT29), .B(new_n555), .C1(new_n472), .C2(new_n473), .ZN(new_n563));
  OR3_X1    g362(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n557), .A2(new_n559), .A3(new_n528), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n556), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n556), .B1(new_n472), .B2(new_n473), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n562), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n553), .B1(new_n564), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT79), .B1(new_n570), .B2(KEYINPUT30), .ZN(new_n571));
  AOI211_X1 g370(.A(new_n561), .B(new_n567), .C1(new_n565), .C2(new_n556), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n560), .A2(new_n563), .A3(new_n562), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT77), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT77), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n564), .A2(new_n569), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n576), .A3(new_n553), .ZN(new_n577));
  INV_X1    g376(.A(new_n553), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n578), .B1(new_n572), .B2(new_n573), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT79), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT30), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n570), .A2(KEYINPUT30), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n571), .A2(new_n577), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT5), .ZN(new_n585));
  NAND2_X1  g384(.A1(G225gat), .A2(G233gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n409), .A2(new_n412), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(G127gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n409), .A2(new_n412), .A3(new_n315), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n589), .A2(new_n511), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n511), .B1(new_n589), .B2(new_n590), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT82), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT82), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n595), .B(new_n587), .C1(new_n591), .C2(new_n592), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n585), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n511), .A2(KEYINPUT3), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n415), .A2(new_n527), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT81), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n415), .A2(KEYINPUT81), .A3(new_n527), .A4(new_n598), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n587), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n510), .B(new_n509), .C1(new_n413), .C2(new_n414), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT4), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT4), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n592), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n597), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G57gat), .B(G85gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT84), .ZN(new_n612));
  XOR2_X1   g411(.A(KEYINPUT83), .B(KEYINPUT0), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G1gat), .B(G29gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n607), .A2(KEYINPUT85), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT86), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n592), .A2(new_n618), .A3(new_n606), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT86), .B1(new_n604), .B2(KEYINPUT4), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n618), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT85), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n623), .B1(new_n592), .B2(new_n606), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n604), .A2(KEYINPUT86), .A3(KEYINPUT4), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n621), .A2(new_n626), .A3(new_n603), .A4(new_n585), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n616), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT87), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n610), .A2(new_n627), .ZN(new_n631));
  INV_X1    g430(.A(new_n616), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT6), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n610), .A2(new_n627), .A3(KEYINPUT87), .A4(new_n616), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n630), .A2(new_n633), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n616), .B1(new_n610), .B2(new_n627), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT6), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n549), .B1(new_n584), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n499), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n601), .A2(new_n602), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n621), .A2(new_n626), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n587), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT89), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n645), .A2(KEYINPUT89), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n642), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n645), .A2(KEYINPUT89), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n591), .A2(new_n592), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n642), .B1(new_n651), .B2(new_n586), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n646), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n649), .A2(new_n653), .A3(new_n616), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n637), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n649), .A2(new_n653), .A3(KEYINPUT40), .A4(new_n616), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(new_n584), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n574), .A2(new_n576), .A3(KEYINPUT37), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT37), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(new_n572), .B2(new_n573), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n553), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT38), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT38), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n562), .B1(new_n560), .B2(new_n563), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n567), .B1(new_n565), .B2(new_n556), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n665), .B(KEYINPUT37), .C1(new_n666), .C2(new_n562), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n661), .A2(new_n664), .A3(new_n553), .A4(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n663), .A2(new_n639), .A3(new_n579), .A4(new_n668), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n545), .A2(new_n548), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n658), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n641), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n491), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n486), .A2(new_n477), .A3(new_n478), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n489), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(new_n670), .A3(new_n492), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n571), .A2(new_n582), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n636), .A2(new_n638), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n577), .A2(new_n583), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n677), .A2(new_n678), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT35), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n584), .A2(new_n676), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT35), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n684), .A3(new_n679), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n402), .B1(new_n672), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n639), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  AND3_X1   g489(.A1(new_n687), .A2(new_n584), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n323), .B1(new_n687), .B2(new_n584), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT42), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(KEYINPUT42), .B2(new_n691), .ZN(G1325gat));
  INV_X1    g493(.A(G15gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n687), .A2(new_n695), .A3(new_n495), .ZN(new_n696));
  INV_X1    g495(.A(new_n499), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n687), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n698), .B2(new_n695), .ZN(G1326gat));
  NAND2_X1  g498(.A1(new_n687), .A2(new_n549), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT43), .B(G22gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  INV_X1    g501(.A(new_n298), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n672), .B2(new_n686), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n373), .A2(new_n336), .A3(new_n400), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR4_X1   g505(.A1(new_n706), .A2(KEYINPUT107), .A3(G29gat), .A4(new_n679), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n704), .A2(new_n705), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n679), .A2(G29gat), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n712));
  OR3_X1    g511(.A1(new_n707), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n684), .B1(new_n683), .B2(new_n679), .ZN(new_n716));
  NOR4_X1   g515(.A1(new_n584), .A2(new_n639), .A3(new_n676), .A4(KEYINPUT35), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n682), .A2(KEYINPUT109), .A3(new_n685), .ZN(new_n719));
  AOI22_X1  g518(.A1(new_n718), .A2(new_n719), .B1(new_n671), .B2(new_n641), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n714), .B1(new_n720), .B2(new_n703), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n704), .A2(KEYINPUT44), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n705), .B(KEYINPUT108), .Z(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G29gat), .B1(new_n725), .B2(new_n679), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n712), .B1(new_n707), .B2(new_n711), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n713), .A2(new_n726), .A3(new_n727), .ZN(G1328gat));
  INV_X1    g527(.A(new_n584), .ZN(new_n729));
  OAI21_X1  g528(.A(G36gat), .B1(new_n725), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT110), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n584), .A2(new_n215), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n706), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n731), .A2(KEYINPUT110), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n730), .A2(new_n736), .ZN(G1329gat));
  NOR2_X1   g536(.A1(new_n499), .A2(new_n207), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n721), .A2(new_n722), .A3(new_n724), .A4(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n495), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n207), .B1(new_n706), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1330gat));
  NAND4_X1  g543(.A1(new_n721), .A2(new_n549), .A3(new_n722), .A4(new_n724), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G50gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT112), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n709), .A2(new_n208), .A3(new_n549), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT48), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n746), .B(new_n748), .C1(KEYINPUT112), .C2(KEYINPUT48), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(G1331gat));
  INV_X1    g552(.A(new_n719), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT109), .B1(new_n682), .B2(new_n685), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n672), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n374), .A2(new_n401), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n756), .A2(KEYINPUT113), .A3(new_n339), .A4(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n339), .A2(new_n757), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n720), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n639), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g564(.A(KEYINPUT49), .B(G64gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n763), .A2(new_n584), .A3(new_n766), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n762), .A2(new_n729), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(G1333gat));
  NAND3_X1  g568(.A1(new_n758), .A2(new_n761), .A3(new_n697), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G71gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n495), .A2(new_n300), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n762), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n771), .B(KEYINPUT50), .C1(new_n762), .C2(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(G1334gat));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n670), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(new_n301), .ZN(G1335gat));
  NOR2_X1   g578(.A1(new_n374), .A2(new_n336), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n756), .A2(new_n298), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT51), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n756), .A2(new_n783), .A3(new_n298), .A4(new_n780), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(new_n400), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(new_n246), .A3(new_n639), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n374), .A2(new_n336), .A3(new_n401), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n721), .A2(new_n639), .A3(new_n722), .A4(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n246), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n790), .B2(new_n789), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n787), .A2(new_n792), .ZN(G1336gat));
  NAND4_X1  g592(.A1(new_n721), .A2(new_n584), .A3(new_n722), .A4(new_n788), .ZN(new_n794));
  INV_X1    g593(.A(new_n245), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n584), .A2(new_n261), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n785), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT52), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n796), .B(new_n800), .C1(new_n785), .C2(new_n797), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(G1337gat));
  AND3_X1   g601(.A1(new_n723), .A2(new_n697), .A3(new_n788), .ZN(new_n803));
  INV_X1    g602(.A(G99gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n495), .A2(new_n804), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n803), .A2(new_n804), .B1(new_n785), .B2(new_n805), .ZN(G1338gat));
  NOR2_X1   g605(.A1(new_n670), .A2(G106gat), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n782), .A2(new_n400), .A3(new_n784), .A4(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n721), .A2(new_n549), .A3(new_n722), .A4(new_n788), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G106gat), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(KEYINPUT115), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(KEYINPUT115), .ZN(new_n814));
  AND4_X1   g613(.A1(new_n808), .A2(new_n810), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n812), .B1(new_n809), .B2(G106gat), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n816), .B2(new_n808), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n815), .A2(new_n817), .ZN(G1339gat));
  NAND3_X1  g617(.A1(new_n381), .A2(new_n382), .A3(new_n385), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n381), .A2(KEYINPUT116), .A3(new_n382), .A4(new_n385), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n823), .A2(new_n386), .A3(KEYINPUT54), .A4(new_n389), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n394), .B1(new_n387), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(new_n397), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n826), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n828), .B(new_n831), .C1(new_n371), .C2(new_n372), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n354), .A2(new_n370), .A3(new_n361), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n351), .A2(new_n341), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n363), .A2(new_n343), .A3(new_n362), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n358), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n400), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n298), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n831), .A2(new_n397), .A3(new_n827), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n833), .A2(new_n836), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n298), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n334), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n335), .A2(new_n373), .A3(new_n337), .A4(new_n401), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n639), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n683), .ZN(new_n847));
  OAI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n373), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n374), .A2(new_n404), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT117), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n848), .B1(new_n847), .B2(new_n850), .ZN(G1340gat));
  NOR2_X1   g650(.A1(new_n847), .A2(new_n401), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(new_n405), .ZN(G1341gat));
  NOR2_X1   g652(.A1(new_n847), .A2(new_n334), .ZN(new_n854));
  XOR2_X1   g653(.A(KEYINPUT73), .B(G127gat), .Z(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(G1342gat));
  NOR2_X1   g655(.A1(new_n847), .A2(new_n703), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n411), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n859), .B(new_n860), .C1(new_n411), .C2(new_n857), .ZN(G1343gat));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n832), .A2(new_n837), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n703), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n298), .A2(new_n840), .A3(new_n839), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n336), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND4_X1   g665(.A1(new_n373), .A2(new_n335), .A3(new_n337), .A4(new_n401), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n862), .B(new_n549), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n499), .A2(new_n729), .A3(new_n639), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n829), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n824), .A2(KEYINPUT118), .A3(new_n826), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n830), .A3(new_n873), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n874), .B(new_n828), .C1(new_n371), .C2(new_n372), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n298), .B1(new_n875), .B2(new_n837), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n334), .B1(new_n876), .B2(new_n841), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n670), .B1(new_n877), .B2(new_n843), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n868), .B(new_n870), .C1(new_n862), .C2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G141gat), .B1(new_n879), .B2(new_n373), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n697), .A2(new_n670), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(KEYINPUT119), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(KEYINPUT119), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n882), .A2(new_n729), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n846), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n373), .A2(G141gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n880), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g687(.A(G148gat), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(KEYINPUT59), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT120), .B(new_n890), .C1(new_n879), .C2(new_n401), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n843), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n549), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(KEYINPUT57), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n670), .B1(new_n842), .B2(new_n843), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n869), .B1(new_n896), .B2(new_n862), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n897), .A3(new_n400), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT120), .B1(new_n898), .B2(new_n890), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n893), .B2(new_n549), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n862), .B(new_n670), .C1(new_n842), .C2(new_n843), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n400), .B(new_n870), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n900), .B1(new_n903), .B2(G148gat), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n892), .A2(new_n899), .A3(new_n904), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n884), .A2(new_n889), .A3(new_n400), .A4(new_n846), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT121), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  INV_X1    g708(.A(new_n899), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n891), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n909), .B(new_n906), .C1(new_n911), .C2(new_n904), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n908), .A2(new_n912), .ZN(G1345gat));
  OAI21_X1  g712(.A(G155gat), .B1(new_n879), .B2(new_n334), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n336), .A2(new_n330), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n885), .B2(new_n915), .ZN(G1346gat));
  NOR3_X1   g715(.A1(new_n879), .A2(new_n504), .A3(new_n703), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n884), .A2(new_n298), .A3(new_n846), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n504), .ZN(G1347gat));
  AOI21_X1  g718(.A(new_n639), .B1(new_n842), .B2(new_n843), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n729), .A2(new_n676), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n373), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(new_n432), .ZN(G1348gat));
  NOR2_X1   g723(.A1(new_n922), .A2(new_n401), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(new_n433), .ZN(G1349gat));
  NOR2_X1   g725(.A1(new_n922), .A2(new_n334), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n452), .A2(G183gat), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n455), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(G183gat), .B2(new_n927), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n931), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g731(.A1(new_n920), .A2(new_n298), .A3(new_n921), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n933), .A2(G190gat), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(G190gat), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT61), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT122), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n938), .A3(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n941), .B1(new_n935), .B2(KEYINPUT61), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT61), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n933), .A2(KEYINPUT123), .A3(new_n943), .A4(G190gat), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n934), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT124), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n948), .B(new_n934), .C1(new_n940), .C2(new_n945), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1351gat));
  OR2_X1    g749(.A1(new_n901), .A2(new_n902), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n697), .A2(new_n639), .A3(new_n729), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(new_n374), .A3(new_n952), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n953), .A2(KEYINPUT126), .ZN(new_n954));
  XNOR2_X1  g753(.A(KEYINPUT125), .B(G197gat), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n956), .B1(new_n953), .B2(KEYINPUT126), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n920), .A2(new_n584), .A3(new_n881), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n374), .A2(new_n955), .ZN(new_n959));
  OAI22_X1  g758(.A1(new_n954), .A2(new_n957), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  NOR3_X1   g759(.A1(new_n958), .A2(G204gat), .A3(new_n401), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT62), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n951), .A2(new_n400), .A3(new_n952), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G204gat), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1353gat));
  NAND2_X1  g764(.A1(new_n951), .A2(new_n952), .ZN(new_n966));
  OAI21_X1  g765(.A(G211gat), .B1(new_n966), .B2(new_n334), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n336), .A2(new_n514), .ZN(new_n971));
  OAI22_X1  g770(.A1(new_n969), .A2(new_n970), .B1(new_n958), .B2(new_n971), .ZN(G1354gat));
  OAI21_X1  g771(.A(G218gat), .B1(new_n966), .B2(new_n703), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n298), .A2(new_n203), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n973), .B1(new_n958), .B2(new_n974), .ZN(G1355gat));
endmodule


