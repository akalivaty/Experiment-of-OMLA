

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583;

  NOR2_X1 U324 ( .A1(n491), .A2(n462), .ZN(n452) );
  INV_X1 U325 ( .A(n541), .ZN(n494) );
  XOR2_X1 U326 ( .A(n450), .B(n449), .Z(n569) );
  XNOR2_X1 U327 ( .A(KEYINPUT97), .B(n395), .ZN(n545) );
  XOR2_X1 U328 ( .A(n443), .B(n442), .Z(n292) );
  INV_X1 U329 ( .A(KEYINPUT47), .ZN(n504) );
  XNOR2_X1 U330 ( .A(n504), .B(KEYINPUT114), .ZN(n505) );
  XNOR2_X1 U331 ( .A(n506), .B(n505), .ZN(n514) );
  XNOR2_X1 U332 ( .A(n300), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U333 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U334 ( .A(n385), .B(n310), .ZN(n311) );
  XNOR2_X1 U335 ( .A(n312), .B(n311), .ZN(n313) );
  NOR2_X1 U336 ( .A1(n551), .A2(n313), .ZN(n562) );
  XNOR2_X1 U337 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U338 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  XOR2_X1 U339 ( .A(G120GAT), .B(KEYINPUT87), .Z(n294) );
  XNOR2_X1 U340 ( .A(G43GAT), .B(KEYINPUT20), .ZN(n293) );
  XNOR2_X1 U341 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U342 ( .A(KEYINPUT86), .B(KEYINPUT84), .Z(n296) );
  XNOR2_X1 U343 ( .A(G113GAT), .B(KEYINPUT85), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U345 ( .A(n298), .B(n297), .Z(n304) );
  XNOR2_X1 U346 ( .A(G134GAT), .B(G127GAT), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n299), .B(KEYINPUT0), .ZN(n351) );
  XOR2_X1 U348 ( .A(n351), .B(G99GAT), .Z(n302) );
  NAND2_X1 U349 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n312) );
  XOR2_X1 U351 ( .A(KEYINPUT88), .B(KEYINPUT17), .Z(n306) );
  XNOR2_X1 U352 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U354 ( .A(KEYINPUT19), .B(n307), .ZN(n385) );
  XOR2_X1 U355 ( .A(G71GAT), .B(G176GAT), .Z(n309) );
  XNOR2_X1 U356 ( .A(G169GAT), .B(G15GAT), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n310) );
  INV_X1 U358 ( .A(n313), .ZN(n550) );
  XOR2_X1 U359 ( .A(KEYINPUT76), .B(KEYINPUT78), .Z(n315) );
  XNOR2_X1 U360 ( .A(G162GAT), .B(KEYINPUT11), .ZN(n314) );
  XNOR2_X1 U361 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U362 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n317) );
  XNOR2_X1 U363 ( .A(KEYINPUT10), .B(KEYINPUT64), .ZN(n316) );
  XNOR2_X1 U364 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U365 ( .A(n319), .B(n318), .Z(n330) );
  XOR2_X1 U366 ( .A(G29GAT), .B(KEYINPUT7), .Z(n321) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(G36GAT), .ZN(n320) );
  XNOR2_X1 U368 ( .A(n321), .B(n320), .ZN(n323) );
  XOR2_X1 U369 ( .A(G50GAT), .B(KEYINPUT8), .Z(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n449) );
  INV_X1 U371 ( .A(n449), .ZN(n328) );
  XNOR2_X1 U372 ( .A(G99GAT), .B(G85GAT), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n324), .B(KEYINPUT73), .ZN(n423) );
  XOR2_X1 U374 ( .A(G190GAT), .B(KEYINPUT79), .Z(n374) );
  XOR2_X1 U375 ( .A(n423), .B(n374), .Z(n326) );
  XNOR2_X1 U376 ( .A(G134GAT), .B(G218GAT), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n330), .B(n329), .ZN(n335) );
  XOR2_X1 U380 ( .A(KEYINPUT75), .B(G92GAT), .Z(n332) );
  NAND2_X1 U381 ( .A1(G232GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U383 ( .A(G106GAT), .B(n333), .Z(n334) );
  XNOR2_X1 U384 ( .A(n335), .B(n334), .ZN(n563) );
  INV_X1 U385 ( .A(n563), .ZN(n457) );
  XNOR2_X1 U386 ( .A(n457), .B(KEYINPUT36), .ZN(n579) );
  XOR2_X1 U387 ( .A(KEYINPUT92), .B(KEYINPUT2), .Z(n337) );
  XNOR2_X1 U388 ( .A(G162GAT), .B(KEYINPUT91), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U390 ( .A(n338), .B(KEYINPUT3), .Z(n340) );
  XNOR2_X1 U391 ( .A(G141GAT), .B(G155GAT), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n373) );
  XOR2_X1 U393 ( .A(KEYINPUT95), .B(KEYINPUT6), .Z(n342) );
  XNOR2_X1 U394 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U396 ( .A(n343), .B(G85GAT), .Z(n345) );
  XOR2_X1 U397 ( .A(G113GAT), .B(G1GAT), .Z(n440) );
  XNOR2_X1 U398 ( .A(G29GAT), .B(n440), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n373), .B(n346), .ZN(n355) );
  XOR2_X1 U401 ( .A(KEYINPUT94), .B(KEYINPUT96), .Z(n348) );
  NAND2_X1 U402 ( .A1(G225GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U404 ( .A(n349), .B(KEYINPUT5), .Z(n353) );
  XNOR2_X1 U405 ( .A(G120GAT), .B(G148GAT), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n350), .B(G57GAT), .ZN(n429) );
  XNOR2_X1 U407 ( .A(n351), .B(n429), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U409 ( .A(n355), .B(n354), .ZN(n395) );
  XOR2_X1 U410 ( .A(KEYINPUT22), .B(KEYINPUT93), .Z(n357) );
  XNOR2_X1 U411 ( .A(G50GAT), .B(KEYINPUT75), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U413 ( .A(G148GAT), .B(KEYINPUT24), .Z(n359) );
  XNOR2_X1 U414 ( .A(KEYINPUT23), .B(KEYINPUT89), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U416 ( .A(n361), .B(n360), .Z(n371) );
  XOR2_X1 U417 ( .A(KEYINPUT90), .B(G218GAT), .Z(n363) );
  XNOR2_X1 U418 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U420 ( .A(G197GAT), .B(n364), .Z(n378) );
  XOR2_X1 U421 ( .A(G78GAT), .B(G204GAT), .Z(n366) );
  XNOR2_X1 U422 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n424) );
  XOR2_X1 U424 ( .A(G22GAT), .B(n424), .Z(n368) );
  NAND2_X1 U425 ( .A1(G228GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n378), .B(n369), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n373), .B(n372), .ZN(n547) );
  XOR2_X1 U430 ( .A(G169GAT), .B(G8GAT), .Z(n444) );
  XOR2_X1 U431 ( .A(n374), .B(n444), .Z(n376) );
  NAND2_X1 U432 ( .A1(G226GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U434 ( .A(n377), .B(G204GAT), .Z(n380) );
  XNOR2_X1 U435 ( .A(G36GAT), .B(n378), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U437 ( .A(n381), .B(KEYINPUT98), .Z(n384) );
  XNOR2_X1 U438 ( .A(G176GAT), .B(G92GAT), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n382), .B(G64GAT), .ZN(n428) );
  XNOR2_X1 U440 ( .A(KEYINPUT80), .B(n428), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n541) );
  NAND2_X1 U443 ( .A1(n550), .A2(n494), .ZN(n387) );
  NAND2_X1 U444 ( .A1(n547), .A2(n387), .ZN(n388) );
  XOR2_X1 U445 ( .A(KEYINPUT25), .B(n388), .Z(n392) );
  NOR2_X1 U446 ( .A1(n550), .A2(n547), .ZN(n389) );
  XOR2_X1 U447 ( .A(KEYINPUT99), .B(n389), .Z(n390) );
  XNOR2_X1 U448 ( .A(n390), .B(KEYINPUT26), .ZN(n567) );
  XOR2_X1 U449 ( .A(n541), .B(KEYINPUT27), .Z(n396) );
  NAND2_X1 U450 ( .A1(n567), .A2(n396), .ZN(n391) );
  NAND2_X1 U451 ( .A1(n392), .A2(n391), .ZN(n393) );
  NAND2_X1 U452 ( .A1(n395), .A2(n393), .ZN(n394) );
  XOR2_X1 U453 ( .A(KEYINPUT100), .B(n394), .Z(n400) );
  NAND2_X1 U454 ( .A1(n396), .A2(n545), .ZN(n516) );
  XOR2_X1 U455 ( .A(KEYINPUT28), .B(KEYINPUT65), .Z(n397) );
  XOR2_X1 U456 ( .A(n547), .B(n397), .Z(n519) );
  OR2_X1 U457 ( .A1(n519), .A2(n550), .ZN(n398) );
  NOR2_X1 U458 ( .A1(n516), .A2(n398), .ZN(n399) );
  NOR2_X2 U459 ( .A1(n400), .A2(n399), .ZN(n461) );
  XOR2_X1 U460 ( .A(KEYINPUT80), .B(G78GAT), .Z(n402) );
  XNOR2_X1 U461 ( .A(G155GAT), .B(G211GAT), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U463 ( .A(G71GAT), .B(KEYINPUT13), .Z(n433) );
  XOR2_X1 U464 ( .A(n403), .B(n433), .Z(n405) );
  XNOR2_X1 U465 ( .A(G183GAT), .B(G127GAT), .ZN(n404) );
  XNOR2_X1 U466 ( .A(n405), .B(n404), .ZN(n410) );
  XNOR2_X1 U467 ( .A(G15GAT), .B(G22GAT), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n406), .B(KEYINPUT66), .ZN(n441) );
  XOR2_X1 U469 ( .A(G57GAT), .B(n441), .Z(n408) );
  NAND2_X1 U470 ( .A1(G231GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U472 ( .A(n410), .B(n409), .Z(n418) );
  XOR2_X1 U473 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n412) );
  XNOR2_X1 U474 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U476 ( .A(KEYINPUT12), .B(G64GAT), .Z(n414) );
  XNOR2_X1 U477 ( .A(G8GAT), .B(G1GAT), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n507) );
  INV_X1 U481 ( .A(n507), .ZN(n576) );
  NOR2_X1 U482 ( .A1(n461), .A2(n576), .ZN(n419) );
  XOR2_X1 U483 ( .A(KEYINPUT102), .B(n419), .Z(n420) );
  NOR2_X1 U484 ( .A1(n579), .A2(n420), .ZN(n422) );
  XOR2_X1 U485 ( .A(KEYINPUT103), .B(KEYINPUT37), .Z(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n491) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n437) );
  XOR2_X1 U488 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n426) );
  NAND2_X1 U489 ( .A1(G230GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U491 ( .A(n427), .B(KEYINPUT32), .Z(n431) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U494 ( .A(n432), .B(KEYINPUT33), .Z(n435) );
  XNOR2_X1 U495 ( .A(n433), .B(KEYINPUT31), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n573) );
  XOR2_X1 U498 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n439) );
  XNOR2_X1 U499 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n448) );
  XOR2_X1 U501 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U502 ( .A1(G229GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n292), .B(n444), .ZN(n446) );
  XNOR2_X1 U504 ( .A(G141GAT), .B(G197GAT), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n450) );
  INV_X1 U507 ( .A(n569), .ZN(n478) );
  XNOR2_X1 U508 ( .A(KEYINPUT69), .B(n478), .ZN(n552) );
  NAND2_X1 U509 ( .A1(n573), .A2(n552), .ZN(n451) );
  XNOR2_X1 U510 ( .A(n451), .B(KEYINPUT74), .ZN(n462) );
  XNOR2_X2 U511 ( .A(n452), .B(KEYINPUT38), .ZN(n474) );
  NAND2_X1 U512 ( .A1(n550), .A2(n474), .ZN(n456) );
  XOR2_X1 U513 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n454) );
  XNOR2_X1 U514 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n453) );
  XNOR2_X1 U515 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n464) );
  XOR2_X1 U516 ( .A(KEYINPUT83), .B(KEYINPUT16), .Z(n459) );
  NAND2_X1 U517 ( .A1(n457), .A2(n576), .ZN(n458) );
  XNOR2_X1 U518 ( .A(n459), .B(n458), .ZN(n460) );
  OR2_X1 U519 ( .A1(n461), .A2(n460), .ZN(n479) );
  NOR2_X1 U520 ( .A1(n462), .A2(n479), .ZN(n469) );
  NAND2_X1 U521 ( .A1(n469), .A2(n545), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n464), .B(n463), .ZN(G1324GAT) );
  NAND2_X1 U523 ( .A1(n494), .A2(n469), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n465), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U525 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n467) );
  NAND2_X1 U526 ( .A1(n469), .A2(n550), .ZN(n466) );
  XNOR2_X1 U527 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U528 ( .A(G15GAT), .B(n468), .Z(G1326GAT) );
  NAND2_X1 U529 ( .A1(n519), .A2(n469), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n470), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U531 ( .A(G29GAT), .B(KEYINPUT39), .Z(n472) );
  NAND2_X1 U532 ( .A1(n474), .A2(n545), .ZN(n471) );
  XNOR2_X1 U533 ( .A(n472), .B(n471), .ZN(G1328GAT) );
  NAND2_X1 U534 ( .A1(n474), .A2(n494), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n473), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n476) );
  NAND2_X1 U537 ( .A1(n474), .A2(n519), .ZN(n475) );
  XNOR2_X1 U538 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U539 ( .A(G50GAT), .B(n477), .ZN(G1331GAT) );
  XNOR2_X1 U540 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n573), .B(KEYINPUT41), .ZN(n533) );
  XNOR2_X1 U542 ( .A(KEYINPUT108), .B(n533), .ZN(n557) );
  NAND2_X1 U543 ( .A1(n557), .A2(n478), .ZN(n490) );
  NOR2_X1 U544 ( .A1(n490), .A2(n479), .ZN(n486) );
  NAND2_X1 U545 ( .A1(n486), .A2(n545), .ZN(n480) );
  XNOR2_X1 U546 ( .A(n481), .B(n480), .ZN(G1332GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n483) );
  NAND2_X1 U548 ( .A1(n486), .A2(n494), .ZN(n482) );
  XNOR2_X1 U549 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U550 ( .A(G64GAT), .B(n484), .ZN(G1333GAT) );
  NAND2_X1 U551 ( .A1(n486), .A2(n550), .ZN(n485) );
  XNOR2_X1 U552 ( .A(n485), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n488) );
  NAND2_X1 U554 ( .A1(n486), .A2(n519), .ZN(n487) );
  XNOR2_X1 U555 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U556 ( .A(G78GAT), .B(n489), .Z(G1335GAT) );
  XNOR2_X1 U557 ( .A(G85GAT), .B(KEYINPUT112), .ZN(n493) );
  NOR2_X1 U558 ( .A1(n491), .A2(n490), .ZN(n497) );
  NAND2_X1 U559 ( .A1(n497), .A2(n545), .ZN(n492) );
  XNOR2_X1 U560 ( .A(n493), .B(n492), .ZN(G1336GAT) );
  NAND2_X1 U561 ( .A1(n494), .A2(n497), .ZN(n495) );
  XNOR2_X1 U562 ( .A(n495), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U563 ( .A1(n497), .A2(n550), .ZN(n496) );
  XNOR2_X1 U564 ( .A(n496), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n499) );
  NAND2_X1 U566 ( .A1(n497), .A2(n519), .ZN(n498) );
  XNOR2_X1 U567 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U568 ( .A(G106GAT), .B(n500), .ZN(G1339GAT) );
  NAND2_X1 U569 ( .A1(n569), .A2(n533), .ZN(n501) );
  XNOR2_X1 U570 ( .A(KEYINPUT46), .B(n501), .ZN(n502) );
  NAND2_X1 U571 ( .A1(n502), .A2(n507), .ZN(n503) );
  NOR2_X1 U572 ( .A1(n563), .A2(n503), .ZN(n506) );
  XNOR2_X1 U573 ( .A(KEYINPUT45), .B(KEYINPUT115), .ZN(n509) );
  NOR2_X1 U574 ( .A1(n579), .A2(n507), .ZN(n508) );
  XOR2_X1 U575 ( .A(n509), .B(n508), .Z(n510) );
  NAND2_X1 U576 ( .A1(n573), .A2(n510), .ZN(n511) );
  NOR2_X1 U577 ( .A1(n552), .A2(n511), .ZN(n512) );
  XNOR2_X1 U578 ( .A(KEYINPUT116), .B(n512), .ZN(n513) );
  NOR2_X1 U579 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(KEYINPUT48), .ZN(n542) );
  NOR2_X1 U581 ( .A1(n542), .A2(n516), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n550), .A2(n530), .ZN(n517) );
  XOR2_X1 U583 ( .A(KEYINPUT117), .B(n517), .Z(n518) );
  NOR2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n552), .A2(n527), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G113GAT), .B(n520), .ZN(G1340GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n522) );
  NAND2_X1 U588 ( .A1(n527), .A2(n557), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G120GAT), .B(n523), .ZN(G1341GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n525) );
  NAND2_X1 U592 ( .A1(n527), .A2(n576), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U594 ( .A(G127GAT), .B(n526), .ZN(G1342GAT) );
  XOR2_X1 U595 ( .A(G134GAT), .B(KEYINPUT51), .Z(n529) );
  NAND2_X1 U596 ( .A1(n527), .A2(n563), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(G1343GAT) );
  NAND2_X1 U598 ( .A1(n567), .A2(n530), .ZN(n531) );
  XOR2_X1 U599 ( .A(KEYINPUT120), .B(n531), .Z(n539) );
  NAND2_X1 U600 ( .A1(n569), .A2(n539), .ZN(n532) );
  XNOR2_X1 U601 ( .A(G141GAT), .B(n532), .ZN(G1344GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT52), .B(KEYINPUT121), .Z(n535) );
  NAND2_X1 U603 ( .A1(n539), .A2(n533), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n535), .B(n534), .ZN(n537) );
  XOR2_X1 U605 ( .A(G148GAT), .B(KEYINPUT53), .Z(n536) );
  XNOR2_X1 U606 ( .A(n537), .B(n536), .ZN(G1345GAT) );
  NAND2_X1 U607 ( .A1(n539), .A2(n576), .ZN(n538) );
  XNOR2_X1 U608 ( .A(n538), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U609 ( .A1(n539), .A2(n563), .ZN(n540) );
  XNOR2_X1 U610 ( .A(n540), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT122), .B(KEYINPUT55), .Z(n549) );
  NOR2_X1 U612 ( .A1(n542), .A2(n541), .ZN(n544) );
  INV_X1 U613 ( .A(KEYINPUT54), .ZN(n543) );
  XNOR2_X1 U614 ( .A(n544), .B(n543), .ZN(n546) );
  NOR2_X1 U615 ( .A1(n546), .A2(n545), .ZN(n566) );
  NAND2_X1 U616 ( .A1(n566), .A2(n547), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(n551) );
  NAND2_X1 U618 ( .A1(n562), .A2(n552), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n555) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U623 ( .A(KEYINPUT123), .B(n556), .Z(n559) );
  NAND2_X1 U624 ( .A1(n557), .A2(n562), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  XOR2_X1 U626 ( .A(G183GAT), .B(KEYINPUT125), .Z(n561) );
  NAND2_X1 U627 ( .A1(n562), .A2(n576), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1350GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT58), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT126), .B(n568), .Z(n577) );
  NAND2_X1 U635 ( .A1(n569), .A2(n577), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .Z(n575) );
  INV_X1 U639 ( .A(n577), .ZN(n580) );
  OR2_X1 U640 ( .A1(n580), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

