//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G116), .A2(G270), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n202), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n211), .B(new_n216), .C1(G97), .C2(G257), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G1), .B2(G20), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT1), .Z(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR3_X1   g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G20), .ZN(new_n224));
  OR3_X1    g0024(.A1(new_n224), .A2(KEYINPUT64), .A3(G13), .ZN(new_n225));
  OAI21_X1  g0025(.A(KEYINPUT64), .B1(new_n224), .B2(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NOR3_X1   g0029(.A1(new_n219), .A2(new_n223), .A3(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G1), .ZN(new_n246));
  OAI211_X1 g0046(.A(new_n246), .B(G274), .C1(G41), .C2(G45), .ZN(new_n247));
  AOI21_X1  g0047(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n246), .B1(G41), .B2(G45), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n247), .B1(new_n251), .B2(new_n213), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n252), .B(KEYINPUT65), .Z(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT66), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT66), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G1698), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n258), .B1(G222), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(new_n259), .ZN(new_n266));
  INV_X1    g0066(.A(new_n258), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n266), .B(new_n248), .C1(G77), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n253), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G200), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n203), .A2(G20), .ZN(new_n271));
  INV_X1    g0071(.A(G150), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n221), .A2(new_n256), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT8), .B(G58), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n221), .A2(G33), .ZN(new_n275));
  OAI221_X1 g0075(.A(new_n271), .B1(new_n272), .B2(new_n273), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n222), .ZN(new_n278));
  INV_X1    g0078(.A(G13), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G1), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n276), .A2(new_n278), .B1(new_n202), .B2(new_n282), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n277), .B(new_n222), .C1(G1), .C2(new_n221), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n283), .B1(new_n202), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT9), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n253), .A2(G190), .A3(new_n268), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n285), .A2(new_n286), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n270), .A2(new_n287), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT10), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n285), .B1(new_n269), .B2(G179), .ZN(new_n292));
  AOI21_X1  g0092(.A(G169), .B1(new_n253), .B2(new_n268), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n263), .A2(G232), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(new_n267), .C1(new_n215), .C2(new_n259), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n298), .B(new_n248), .C1(G107), .C2(new_n267), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n299), .B(new_n247), .C1(new_n208), .C2(new_n251), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n300), .A2(G179), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n281), .A2(G77), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n273), .A2(KEYINPUT67), .ZN(new_n303));
  INV_X1    g0103(.A(new_n274), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n273), .A2(KEYINPUT67), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  XOR2_X1   g0106(.A(KEYINPUT15), .B(G87), .Z(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n306), .B1(new_n221), .B2(new_n207), .C1(new_n275), .C2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n302), .B1(new_n309), .B2(new_n278), .ZN(new_n310));
  INV_X1    g0110(.A(new_n284), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G77), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n300), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n301), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n296), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT14), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G97), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n263), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n258), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n248), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n249), .A2(G238), .A3(new_n250), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(new_n247), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT13), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT13), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n323), .A2(new_n327), .A3(new_n247), .A4(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n319), .B1(new_n329), .B2(G169), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  AOI211_X1 g0131(.A(KEYINPUT14), .B(new_n314), .C1(new_n326), .C2(new_n328), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n331), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n273), .A2(new_n202), .B1(new_n275), .B2(new_n207), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n221), .A2(G68), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n278), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT11), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n340), .A2(new_n341), .B1(new_n214), .B2(new_n284), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n340), .A2(new_n341), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n280), .A2(new_n339), .ZN(new_n344));
  XOR2_X1   g0144(.A(new_n344), .B(KEYINPUT12), .Z(new_n345));
  NOR3_X1   g0145(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n337), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G190), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n346), .B1(new_n329), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G200), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(new_n326), .B2(new_n328), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n318), .A2(new_n348), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n278), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n221), .A2(KEYINPUT7), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n256), .A2(KEYINPUT68), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT68), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G33), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n360), .A3(new_n254), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n357), .B1(new_n361), .B2(new_n257), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT7), .B1(new_n258), .B2(new_n221), .ZN(new_n363));
  OAI21_X1  g0163(.A(G68), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AND2_X1   g0164(.A1(G58), .A2(G68), .ZN(new_n365));
  OAI21_X1  g0165(.A(G20), .B1(new_n365), .B2(new_n201), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT69), .ZN(new_n367));
  INV_X1    g0167(.A(new_n273), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G159), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT69), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(G20), .C1(new_n365), .C2(new_n201), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n367), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n364), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT70), .B(KEYINPUT16), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n356), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n254), .B1(new_n358), .B2(new_n360), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n376), .B(new_n221), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G68), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT68), .B(G33), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n255), .B1(new_n381), .B2(new_n254), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n376), .B1(new_n382), .B2(new_n221), .ZN(new_n383));
  OAI211_X1 g0183(.A(KEYINPUT16), .B(new_n372), .C1(new_n380), .C2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT71), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n304), .A2(new_n284), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n281), .A2(new_n274), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(new_n385), .A3(new_n387), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(KEYINPUT72), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT72), .ZN(new_n392));
  INV_X1    g0192(.A(new_n390), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(new_n388), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n375), .A2(new_n384), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n249), .A2(G232), .A3(new_n250), .ZN(new_n396));
  XNOR2_X1  g0196(.A(KEYINPUT66), .B(G1698), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n397), .A2(new_n265), .B1(new_n213), .B2(new_n259), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n358), .A2(new_n360), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n378), .B1(new_n399), .B2(KEYINPUT3), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n398), .A2(new_n400), .B1(G33), .B2(G87), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n396), .B(new_n247), .C1(new_n401), .C2(new_n249), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n351), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G190), .B2(new_n402), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n395), .A2(new_n404), .A3(KEYINPUT17), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT17), .B1(new_n395), .B2(new_n404), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n373), .A2(new_n374), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(new_n278), .A3(new_n384), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n394), .A2(new_n391), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n402), .A2(G169), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n334), .B2(new_n402), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT18), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n411), .A2(new_n413), .A3(KEYINPUT18), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n310), .A2(new_n312), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n300), .A2(G200), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n419), .B(new_n420), .C1(new_n349), .C2(new_n300), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n407), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n355), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT5), .B(G41), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n246), .A2(G45), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G274), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n249), .A3(G270), .ZN(new_n431));
  INV_X1    g0231(.A(G303), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n255), .B2(new_n257), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G264), .A2(G1698), .ZN(new_n434));
  INV_X1    g0234(.A(G257), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n434), .B1(new_n397), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n433), .B1(new_n400), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n430), .B(new_n431), .C1(new_n437), .C2(new_n249), .ZN(new_n438));
  INV_X1    g0238(.A(G116), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n277), .A2(new_n222), .B1(G20), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G283), .ZN(new_n441));
  INV_X1    g0241(.A(G97), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n441), .B(new_n221), .C1(G33), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT20), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n445), .A2(KEYINPUT77), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(KEYINPUT77), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n280), .A2(G20), .A3(new_n439), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n246), .A2(G33), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n356), .A2(new_n281), .A3(G116), .A4(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n440), .A2(KEYINPUT77), .A3(new_n443), .A4(new_n445), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n448), .A2(new_n449), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n438), .A2(new_n454), .A3(new_n334), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n438), .A2(G169), .A3(new_n453), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT21), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT21), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n438), .A2(new_n458), .A3(G169), .A4(new_n453), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n455), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n438), .A2(G200), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n461), .B(new_n454), .C1(new_n349), .C2(new_n438), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n282), .A2(new_n442), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n356), .A2(new_n281), .A3(new_n450), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G97), .ZN(new_n467));
  OAI21_X1  g0267(.A(G107), .B1(new_n362), .B2(new_n363), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n368), .A2(G77), .ZN(new_n469));
  INV_X1    g0269(.A(G107), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(KEYINPUT6), .A3(G97), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n442), .A2(new_n470), .ZN(new_n472));
  NOR2_X1   g0272(.A1(G97), .A2(G107), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n471), .B1(new_n474), .B2(KEYINPUT6), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G20), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n468), .A2(new_n469), .A3(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n464), .B(new_n467), .C1(new_n477), .C2(new_n356), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n428), .A2(new_n249), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n430), .B1(new_n435), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n359), .A2(G33), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n256), .A2(KEYINPUT68), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT3), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n483), .A2(G244), .A3(new_n255), .A4(new_n263), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n397), .A2(new_n485), .A3(new_n208), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n210), .A2(new_n259), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n267), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n486), .A2(new_n489), .A3(new_n441), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n480), .B1(new_n490), .B2(new_n248), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n478), .B1(G190), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n248), .ZN(new_n493));
  INV_X1    g0293(.A(new_n480), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G200), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n491), .A2(new_n334), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT73), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n484), .A2(new_n485), .B1(G33), .B2(G283), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n249), .B1(new_n500), .B2(new_n489), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n314), .B1(new_n501), .B2(new_n480), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT73), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n491), .A2(new_n503), .A3(new_n334), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n499), .A2(new_n502), .A3(new_n478), .A4(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n428), .A2(new_n249), .A3(G264), .ZN(new_n506));
  INV_X1    g0306(.A(G294), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n399), .A2(new_n507), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n397), .A2(new_n210), .B1(new_n435), .B2(new_n259), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(new_n400), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n430), .B(new_n506), .C1(new_n510), .C2(new_n249), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G169), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT78), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n511), .A2(new_n334), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n511), .A2(KEYINPUT78), .A3(G169), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n470), .A2(G20), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n280), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT25), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n465), .A2(new_n470), .B1(KEYINPUT25), .B2(new_n521), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n358), .A2(new_n360), .A3(G116), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n209), .A2(G20), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(new_n255), .A3(new_n257), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT22), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n528), .A2(new_n221), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n483), .A2(KEYINPUT22), .A3(new_n255), .A4(new_n529), .ZN(new_n533));
  XOR2_X1   g0333(.A(new_n519), .B(KEYINPUT23), .Z(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT24), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT24), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n532), .A2(new_n533), .A3(new_n537), .A4(new_n534), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n525), .B(new_n527), .C1(new_n539), .C2(new_n356), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n518), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n356), .B1(new_n536), .B2(new_n538), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n542), .A2(new_n524), .A3(new_n526), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n511), .A2(new_n351), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(G190), .B2(new_n511), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n497), .A2(new_n505), .A3(new_n541), .A4(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT75), .ZN(new_n548));
  OAI211_X1 g0348(.A(G244), .B(new_n255), .C1(new_n381), .C2(new_n254), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(new_n259), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n397), .A2(new_n215), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n528), .B1(new_n400), .B2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n400), .A2(KEYINPUT75), .A3(G244), .A4(G1698), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n248), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT74), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n426), .A2(new_n556), .A3(G250), .ZN(new_n557));
  AOI21_X1  g0357(.A(G274), .B1(KEYINPUT74), .B2(G250), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n557), .B1(new_n426), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n249), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n314), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT76), .ZN(new_n563));
  NOR4_X1   g0363(.A1(new_n377), .A2(G20), .A3(new_n214), .A4(new_n378), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n320), .A2(KEYINPUT19), .A3(G20), .ZN(new_n565));
  NOR2_X1   g0365(.A1(G87), .A2(G97), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n470), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n320), .A2(new_n221), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n565), .B1(new_n569), .B2(KEYINPUT19), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n278), .B1(new_n564), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n307), .A2(new_n281), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n563), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n483), .A2(new_n221), .A3(G68), .A4(new_n255), .ZN(new_n575));
  INV_X1    g0375(.A(new_n565), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n566), .A2(new_n470), .B1(new_n320), .B2(new_n221), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n356), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n580), .A2(KEYINPUT76), .A3(new_n572), .ZN(new_n581));
  OAI22_X1  g0381(.A1(new_n574), .A2(new_n581), .B1(new_n308), .B2(new_n465), .ZN(new_n582));
  INV_X1    g0382(.A(new_n560), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n583), .B1(new_n554), .B2(new_n248), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n334), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n562), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n465), .A2(new_n209), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n571), .A2(new_n563), .A3(new_n573), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT76), .B1(new_n580), .B2(new_n572), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n555), .A2(G190), .A3(new_n560), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n590), .B(new_n591), .C1(new_n351), .C2(new_n584), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n586), .A2(new_n592), .ZN(new_n593));
  NOR4_X1   g0393(.A1(new_n424), .A2(new_n463), .A3(new_n547), .A4(new_n593), .ZN(G372));
  AND2_X1   g0394(.A1(new_n582), .A2(new_n585), .ZN(new_n595));
  XOR2_X1   g0395(.A(new_n560), .B(KEYINPUT79), .Z(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n555), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n314), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n511), .A2(KEYINPUT78), .A3(G169), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT78), .B1(new_n511), .B2(G169), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n601), .A2(new_n602), .A3(new_n515), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n460), .B1(new_n603), .B2(new_n543), .ZN(new_n604));
  INV_X1    g0404(.A(new_n597), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n591), .B(new_n590), .C1(new_n605), .C2(new_n351), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n604), .A2(new_n497), .A3(new_n546), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n502), .A2(new_n478), .ZN(new_n608));
  NOR4_X1   g0408(.A1(new_n501), .A2(KEYINPUT73), .A3(G179), .A4(new_n480), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n503), .B1(new_n491), .B2(new_n334), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT26), .B1(new_n611), .B2(new_n606), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n593), .A2(new_n505), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT26), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n600), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n424), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g0417(.A(new_n617), .B(KEYINPUT80), .Z(new_n618));
  OAI21_X1  g0418(.A(new_n348), .B1(new_n353), .B2(new_n316), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT81), .ZN(new_n620));
  OR2_X1    g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n407), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n418), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n294), .B1(new_n624), .B2(new_n291), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n618), .A2(new_n625), .ZN(G369));
  INV_X1    g0426(.A(G330), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n279), .A2(G20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n246), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(G213), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(G343), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n454), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n463), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n460), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n636), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT82), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT82), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n637), .A2(new_n642), .A3(new_n639), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n627), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n541), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n645), .A2(KEYINPUT83), .A3(new_n634), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT83), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n541), .B2(new_n635), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n541), .B(new_n546), .C1(new_n543), .C2(new_n635), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n460), .A2(new_n634), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n651), .A2(new_n653), .B1(new_n645), .B2(new_n635), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(G399));
  OAI21_X1  g0455(.A(KEYINPUT86), .B1(new_n616), .B2(new_n634), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT29), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT86), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n607), .A2(new_n612), .B1(new_n614), .B2(KEYINPUT26), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n658), .B(new_n635), .C1(new_n659), .C2(new_n600), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n656), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT87), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n611), .A2(new_n606), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT26), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n600), .B1(new_n614), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n497), .A2(new_n505), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(KEYINPUT88), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT88), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n497), .B2(new_n505), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n604), .A2(new_n546), .A3(new_n606), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n665), .B(new_n667), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(KEYINPUT29), .A3(new_n635), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n656), .A2(KEYINPUT87), .A3(new_n657), .A4(new_n660), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n663), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n605), .A2(G179), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT84), .ZN(new_n679));
  INV_X1    g0479(.A(new_n511), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n491), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n491), .A2(new_n680), .A3(new_n679), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n678), .B(new_n438), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT85), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n683), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n681), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n688), .A2(KEYINPUT85), .A3(new_n438), .A4(new_n678), .ZN(new_n689));
  INV_X1    g0489(.A(new_n437), .ZN(new_n690));
  INV_X1    g0490(.A(new_n479), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n690), .A2(new_n248), .B1(G270), .B2(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n515), .A2(new_n491), .A3(new_n584), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT30), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n686), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n634), .ZN(new_n696));
  NOR4_X1   g0496(.A1(new_n547), .A2(new_n463), .A3(new_n593), .A4(new_n634), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n694), .A2(new_n684), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(KEYINPUT31), .A3(new_n634), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n677), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n246), .ZN(new_n705));
  INV_X1    g0505(.A(new_n227), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n566), .A2(new_n470), .A3(new_n439), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n707), .A2(new_n246), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n220), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(new_n707), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT28), .Z(new_n712));
  NAND2_X1  g0512(.A1(new_n705), .A2(new_n712), .ZN(G364));
  NAND2_X1  g0513(.A1(new_n641), .A2(new_n643), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n628), .A2(G45), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n716), .A2(KEYINPUT89), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(KEYINPUT89), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n707), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n715), .A2(new_n644), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g0521(.A(new_n721), .B(KEYINPUT90), .Z(new_n722));
  NOR2_X1   g0522(.A1(new_n334), .A2(new_n351), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n221), .A2(G190), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G317), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT33), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n727), .A2(KEYINPUT33), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G179), .A2(G200), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n724), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G329), .ZN(new_n734));
  INV_X1    g0534(.A(G283), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n351), .A2(G179), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n724), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n730), .B(new_n734), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n221), .A2(new_n349), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n334), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n267), .B(new_n738), .C1(G322), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n740), .A2(new_n724), .ZN(new_n744));
  INV_X1    g0544(.A(G311), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n221), .B1(new_n731), .B2(G190), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n744), .A2(new_n745), .B1(new_n746), .B2(new_n507), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n739), .A2(new_n723), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n747), .B1(G326), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT92), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n739), .A2(new_n736), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n743), .B(new_n751), .C1(new_n432), .C2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G58), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n754), .A2(new_n741), .B1(new_n752), .B2(new_n209), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n267), .B1(new_n737), .B2(new_n470), .C1(new_n214), .C2(new_n725), .ZN(new_n756));
  INV_X1    g0556(.A(new_n744), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n755), .B(new_n756), .C1(G77), .C2(new_n757), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n746), .A2(KEYINPUT91), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n746), .A2(KEYINPUT91), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G97), .ZN(new_n763));
  INV_X1    g0563(.A(G159), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n732), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT32), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n758), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n748), .A2(new_n202), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n753), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n222), .B1(G20), .B2(new_n314), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n770), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n706), .A2(new_n258), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G355), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n706), .A2(new_n400), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G45), .B2(new_n220), .ZN(new_n778));
  INV_X1    g0578(.A(G45), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n241), .A2(new_n779), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n776), .B1(G116), .B2(new_n227), .C1(new_n778), .C2(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n769), .A2(new_n770), .B1(new_n774), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n773), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n720), .B(new_n782), .C1(new_n714), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n722), .A2(new_n784), .ZN(G396));
  NAND2_X1  g0585(.A1(new_n313), .A2(new_n634), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n421), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n317), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n316), .A2(new_n634), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n656), .A2(new_n660), .A3(new_n791), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n635), .B(new_n790), .C1(new_n659), .C2(new_n600), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n703), .ZN(new_n795));
  INV_X1    g0595(.A(new_n720), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n794), .A2(new_n703), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G143), .A2(new_n742), .B1(new_n726), .B2(G150), .ZN(new_n799));
  INV_X1    g0599(.A(G137), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n799), .B1(new_n800), .B2(new_n748), .C1(new_n764), .C2(new_n744), .ZN(new_n801));
  XOR2_X1   g0601(.A(KEYINPUT94), .B(KEYINPUT34), .Z(new_n802));
  XNOR2_X1  g0602(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G132), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n737), .A2(new_n214), .B1(new_n732), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n746), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n382), .B(new_n805), .C1(G58), .C2(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n803), .B(new_n807), .C1(new_n202), .C2(new_n752), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n741), .A2(new_n507), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n748), .A2(new_n432), .B1(new_n725), .B2(new_n735), .ZN(new_n810));
  INV_X1    g0610(.A(new_n752), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n809), .B(new_n810), .C1(G107), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n737), .A2(new_n209), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n258), .B1(new_n744), .B2(new_n439), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G311), .B2(new_n733), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n812), .A2(new_n763), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n808), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n770), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n770), .A2(new_n771), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n720), .B1(G77), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT93), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n819), .B(new_n823), .C1(new_n790), .C2(new_n772), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n798), .A2(new_n824), .ZN(G384));
  INV_X1    g0625(.A(new_n789), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n793), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n347), .B(new_n634), .C1(new_n337), .C2(new_n353), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n347), .A2(new_n634), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n330), .A2(new_n332), .A3(new_n335), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n354), .B(new_n829), .C1(new_n830), .C2(new_n346), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n827), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT96), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n827), .A2(KEYINPUT96), .A3(new_n833), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n632), .B(KEYINPUT97), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n411), .B1(new_n413), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT37), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n395), .A2(new_n404), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT98), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n839), .A2(KEYINPUT98), .A3(new_n840), .A4(new_n841), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n372), .B1(new_n380), .B2(new_n383), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n847), .A2(new_n374), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n384), .A2(new_n278), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n389), .A2(new_n390), .ZN(new_n851));
  INV_X1    g0651(.A(new_n632), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n850), .A2(new_n851), .B1(new_n413), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n840), .B1(new_n853), .B2(new_n841), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n846), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n852), .B1(new_n850), .B2(new_n851), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n407), .B2(new_n418), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n856), .A2(new_n859), .A3(KEYINPUT38), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n854), .B1(new_n844), .B2(new_n845), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n861), .B1(new_n862), .B2(new_n858), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n860), .A2(new_n863), .A3(KEYINPUT99), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT99), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n865), .B(new_n861), .C1(new_n862), .C2(new_n858), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(KEYINPUT100), .A3(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT100), .B1(new_n864), .B2(new_n866), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n836), .B(new_n837), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n418), .A2(new_n838), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n870), .A2(KEYINPUT101), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT101), .B1(new_n870), .B2(new_n872), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n846), .A2(KEYINPUT103), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n839), .A2(new_n841), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT102), .B1(new_n876), .B2(new_n840), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT103), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n844), .A2(new_n878), .A3(new_n845), .ZN(new_n879));
  OR3_X1    g0679(.A1(new_n876), .A2(KEYINPUT102), .A3(new_n840), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n875), .A2(new_n877), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n407), .A2(new_n418), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(new_n411), .A3(new_n838), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT38), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n860), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT39), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n864), .A2(KEYINPUT39), .A3(new_n866), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n348), .A2(new_n634), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n873), .A2(new_n874), .A3(new_n891), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n663), .A2(new_n675), .A3(new_n423), .A4(new_n676), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n625), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n892), .B(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n695), .A2(KEYINPUT31), .A3(new_n634), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n791), .B(new_n832), .C1(new_n699), .C2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n868), .B2(new_n869), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n884), .A2(new_n885), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(KEYINPUT40), .A3(new_n897), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n699), .A2(new_n896), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n423), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n903), .B(new_n905), .Z(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(G330), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n895), .B(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n246), .B2(new_n628), .ZN(new_n909));
  OAI21_X1  g0709(.A(G77), .B1(new_n754), .B2(new_n214), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n910), .A2(new_n220), .B1(G50), .B2(new_n214), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(G1), .A3(new_n279), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n439), .B1(new_n475), .B2(KEYINPUT35), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n222), .A2(new_n221), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n913), .B(new_n914), .C1(KEYINPUT35), .C2(new_n475), .ZN(new_n915));
  XOR2_X1   g0715(.A(KEYINPUT95), .B(KEYINPUT36), .Z(new_n916));
  XNOR2_X1  g0716(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n909), .A2(new_n912), .A3(new_n917), .ZN(G367));
  INV_X1    g0718(.A(new_n737), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(G97), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n920), .B1(new_n735), .B2(new_n744), .C1(new_n727), .C2(new_n732), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(G303), .B2(new_n742), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n752), .A2(new_n439), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT46), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(G107), .B2(new_n806), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n726), .A2(G294), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n400), .B1(G311), .B2(new_n749), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n922), .A2(new_n925), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n737), .A2(new_n207), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(G150), .B2(new_n742), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n764), .B2(new_n725), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(G50), .B2(new_n757), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n762), .A2(G68), .ZN(new_n933));
  INV_X1    g0733(.A(G143), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n267), .B1(new_n748), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(G137), .B2(new_n733), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n932), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n752), .A2(new_n754), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n928), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n796), .B1(new_n941), .B2(new_n770), .ZN(new_n942));
  INV_X1    g0742(.A(new_n777), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n774), .B1(new_n227), .B2(new_n308), .C1(new_n943), .C2(new_n237), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n590), .A2(new_n635), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n599), .A2(new_n606), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n599), .B2(new_n945), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n942), .B(new_n944), .C1(new_n947), .C2(new_n783), .ZN(new_n948));
  INV_X1    g0748(.A(new_n652), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n668), .B(KEYINPUT88), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n478), .A2(new_n634), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n505), .A2(new_n635), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(new_n654), .A3(KEYINPUT45), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT45), .B1(new_n955), .B2(new_n654), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n654), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n953), .B1(new_n950), .B2(new_n951), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT44), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT44), .B1(new_n955), .B2(new_n654), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n949), .B1(new_n959), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT45), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n960), .B2(new_n961), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n956), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n969), .A2(new_n652), .A3(new_n964), .A4(new_n963), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n651), .A2(new_n653), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT106), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n974), .A2(new_n644), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n644), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n975), .A2(new_n976), .B1(new_n651), .B2(new_n653), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n974), .A2(new_n644), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n651), .A2(new_n653), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n974), .A2(new_n644), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n703), .B(new_n677), .C1(new_n971), .C2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n707), .B(KEYINPUT41), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n719), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n950), .A2(new_n645), .A3(new_n951), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n505), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n635), .ZN(new_n988));
  OAI21_X1  g0788(.A(KEYINPUT42), .B1(new_n961), .B2(new_n972), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT105), .ZN(new_n991));
  OR3_X1    g0791(.A1(new_n961), .A2(new_n972), .A3(KEYINPUT42), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT105), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n988), .A2(new_n993), .A3(new_n989), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n947), .B(KEYINPUT104), .Z(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n995), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n991), .A2(new_n992), .A3(new_n994), .A4(new_n998), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n652), .A2(new_n961), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1000), .A2(new_n1003), .A3(new_n1001), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n948), .B1(new_n985), .B2(new_n1007), .ZN(G387));
  NAND2_X1  g0808(.A1(new_n977), .A2(new_n981), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n719), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G311), .A2(new_n726), .B1(new_n742), .B2(G317), .ZN(new_n1011));
  INV_X1    g0811(.A(G322), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1011), .B1(new_n432), .B2(new_n744), .C1(new_n1012), .C2(new_n748), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT48), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n735), .B2(new_n746), .C1(new_n507), .C2(new_n752), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT109), .Z(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT49), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(KEYINPUT49), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n733), .A2(G326), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n400), .B1(G116), .B2(new_n919), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n744), .A2(new_n214), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n811), .A2(G77), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n274), .B2(new_n725), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G50), .B2(new_n742), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n920), .B1(new_n764), .B2(new_n748), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G150), .B2(new_n733), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n762), .A2(new_n307), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1025), .A2(new_n1027), .A3(new_n400), .A4(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1021), .B1(new_n1022), .B2(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n775), .A2(new_n708), .B1(new_n470), .B2(new_n706), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n304), .A2(new_n202), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n708), .B1(new_n1032), .B2(KEYINPUT50), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n779), .C1(KEYINPUT50), .C2(new_n1032), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n214), .A2(new_n207), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n777), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT108), .Z(new_n1037));
  NOR2_X1   g0837(.A1(new_n234), .A2(new_n779), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1031), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1030), .A2(new_n770), .B1(new_n774), .B2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1040), .B(new_n720), .C1(new_n651), .C2(new_n783), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n982), .A2(new_n704), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(KEYINPUT110), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1009), .A2(new_n703), .A3(new_n677), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n707), .B1(new_n1042), .B2(KEYINPUT110), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1010), .B(new_n1041), .C1(new_n1045), .C2(new_n1046), .ZN(G393));
  OR2_X1    g0847(.A1(new_n971), .A2(new_n1044), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n707), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n971), .B2(new_n1044), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n966), .A2(new_n970), .A3(new_n719), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n774), .B1(new_n442), .B2(new_n227), .C1(new_n943), .C2(new_n244), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n258), .B1(new_n744), .B2(new_n507), .C1(new_n470), .C2(new_n737), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G116), .B2(new_n806), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n748), .A2(new_n727), .B1(new_n741), .B2(new_n745), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT52), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n726), .A2(G303), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n752), .A2(new_n735), .B1(new_n732), .B2(new_n1012), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT112), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n744), .A2(new_n274), .B1(new_n732), .B2(new_n934), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n761), .A2(new_n207), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(G68), .C2(new_n811), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n748), .A2(new_n272), .B1(new_n741), .B2(new_n764), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT111), .Z(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT51), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n382), .B(new_n813), .C1(G50), .C2(new_n726), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1066), .B2(KEYINPUT51), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1061), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n796), .B1(new_n1071), .B2(new_n770), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1053), .B(new_n1072), .C1(new_n955), .C2(new_n783), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1051), .A2(new_n1052), .A3(new_n1073), .ZN(G390));
  NAND3_X1  g0874(.A1(new_n423), .A2(G330), .A3(new_n904), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n893), .A2(new_n625), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n790), .A2(G330), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n833), .B1(new_n904), .B2(new_n1078), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1077), .B(new_n832), .C1(new_n699), .C2(new_n701), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n674), .B(new_n635), .C1(new_n317), .C2(new_n787), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1082), .A2(new_n826), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n547), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n463), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n593), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .A4(new_n635), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1087), .A2(KEYINPUT31), .B1(new_n634), .B2(new_n695), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n896), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n833), .B(new_n1078), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1077), .B1(new_n699), .B2(new_n701), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1090), .B1(new_n833), .B2(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1081), .A2(new_n1083), .B1(new_n1092), .B2(new_n827), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1076), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1090), .A2(KEYINPUT113), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n889), .B1(new_n827), .B2(new_n833), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n886), .A2(new_n887), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n832), .B1(new_n1082), .B2(new_n826), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n884), .A2(new_n885), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n1098), .A2(new_n1099), .A3(new_n889), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1095), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1097), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n901), .B(new_n890), .C1(new_n1083), .C2(new_n832), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n904), .A2(KEYINPUT113), .A3(new_n1078), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n1080), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1102), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1094), .A2(new_n1101), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT114), .B1(new_n1107), .B2(new_n707), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1106), .A2(new_n1101), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(KEYINPUT115), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1076), .A2(new_n1093), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT115), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1106), .A2(new_n1101), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1111), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1107), .A2(KEYINPUT114), .A3(new_n707), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1109), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n888), .A2(new_n771), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n748), .A2(new_n735), .B1(new_n744), .B2(new_n442), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G107), .B2(new_n726), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT117), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(G68), .A2(new_n919), .B1(new_n733), .B2(G294), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1063), .B1(G116), .B2(new_n742), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n258), .B1(new_n752), .B2(new_n209), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT118), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(G128), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n748), .A2(new_n1127), .B1(new_n744), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n811), .A2(G150), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT53), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1129), .B(new_n1131), .C1(G132), .C2(new_n742), .ZN(new_n1132));
  INV_X1    g0932(.A(G125), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n267), .B1(new_n732), .B2(new_n1133), .C1(new_n202), .C2(new_n737), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(KEYINPUT116), .A2(new_n1135), .B1(new_n762), .B2(G159), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1132), .B(new_n1136), .C1(KEYINPUT116), .C2(new_n1135), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n725), .A2(new_n800), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1126), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1139), .A2(new_n770), .B1(new_n274), .B2(new_n820), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1118), .A2(new_n720), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n719), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(new_n1110), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1117), .A2(new_n1144), .ZN(G378));
  NAND3_X1  g0945(.A1(new_n904), .A2(new_n790), .A3(new_n833), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n864), .A2(new_n866), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT100), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1146), .B1(new_n1149), .B2(new_n867), .ZN(new_n1150));
  OAI211_X1 g0950(.A(G330), .B(new_n902), .C1(new_n1150), .C2(KEYINPUT40), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n296), .B(KEYINPUT55), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n285), .A2(new_n852), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT56), .Z(new_n1154));
  XNOR2_X1  g0954(.A(new_n1152), .B(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1155), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n900), .A2(G330), .A3(new_n902), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT120), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1159), .B1(new_n892), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n870), .A2(new_n872), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT101), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n891), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n870), .A2(KEYINPUT101), .A3(new_n872), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1167), .A2(KEYINPUT120), .A3(new_n1158), .A4(new_n1156), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1076), .B(KEYINPUT121), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1107), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1161), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n873), .A2(new_n874), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1174), .A2(new_n1165), .A3(new_n1158), .A4(new_n1156), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1159), .A2(new_n1167), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1172), .B1(new_n1107), .B2(new_n1169), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1049), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1173), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1161), .A2(new_n719), .A3(new_n1168), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1155), .A2(new_n771), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n820), .A2(new_n202), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G58), .A2(new_n919), .B1(new_n733), .B2(G283), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n308), .B2(new_n744), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1023), .B1(new_n442), .B2(new_n725), .C1(new_n439), .C2(new_n748), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(G107), .C2(new_n742), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n400), .A2(G41), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n933), .A3(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT58), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n748), .A2(new_n1133), .B1(new_n744), .B2(new_n800), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n1127), .A2(new_n741), .B1(new_n725), .B2(new_n804), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(new_n762), .C2(G150), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n752), .B2(new_n1128), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n733), .A2(G124), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(G33), .A2(G41), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT119), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G159), .B2(new_n919), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n202), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1190), .B(new_n1201), .C1(new_n1188), .C2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n796), .B1(new_n1203), .B2(new_n770), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1182), .A2(new_n1183), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1181), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1180), .A2(new_n1207), .ZN(G375));
  NAND2_X1  g1008(.A1(new_n1076), .A2(new_n1093), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1112), .A2(new_n984), .A3(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1093), .A2(new_n1142), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n744), .A2(new_n470), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n748), .A2(new_n507), .B1(new_n741), .B2(new_n735), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(G97), .C2(new_n811), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n726), .A2(G116), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n267), .B(new_n929), .C1(G303), .C2(new_n733), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1214), .A2(new_n1028), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n382), .B1(G58), .B2(new_n919), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT122), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n725), .A2(new_n1128), .B1(new_n732), .B2(new_n1127), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n748), .A2(new_n804), .B1(new_n744), .B2(new_n272), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(G159), .C2(new_n811), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1219), .B(new_n1222), .C1(new_n202), .C2(new_n761), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n741), .A2(new_n800), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1217), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n770), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(G68), .B2(new_n821), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n832), .B2(new_n771), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1211), .B1(new_n720), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1210), .A2(new_n1229), .ZN(G381));
  AOI21_X1  g1030(.A(new_n1206), .B1(new_n1173), .B2(new_n1179), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1107), .A2(KEYINPUT114), .A3(new_n707), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(new_n1108), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1143), .B1(new_n1233), .B2(new_n1115), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n983), .A2(new_n984), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1142), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1051), .A2(new_n1052), .A3(new_n1073), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n1241), .A3(new_n948), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1243));
  INV_X1    g1043(.A(G396), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1243), .A2(new_n1244), .A3(new_n1010), .A4(new_n1041), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(new_n1242), .A2(new_n1245), .A3(G384), .A4(G381), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1236), .A2(new_n1246), .ZN(G407));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n633), .ZN(new_n1248));
  OAI21_X1  g1048(.A(G213), .B1(new_n1248), .B2(new_n1235), .ZN(G409));
  NAND2_X1  g1049(.A1(G387), .A2(G390), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1242), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1245), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1245), .A2(new_n1252), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(new_n1242), .A3(new_n1250), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT125), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1257), .B(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G375), .A2(G378), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT62), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT60), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1209), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1076), .A2(new_n1093), .A3(KEYINPUT60), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1263), .A2(new_n1112), .A3(new_n707), .A4(new_n1264), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1265), .A2(G384), .A3(new_n1229), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G384), .B1(new_n1265), .B2(new_n1229), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(G213), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(G343), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1161), .A2(new_n1168), .A3(new_n984), .A4(new_n1170), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1159), .A2(new_n1167), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1174), .A2(new_n1165), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n719), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1271), .A2(new_n1274), .A3(new_n1205), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1270), .B1(new_n1275), .B2(new_n1234), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1260), .A2(new_n1261), .A3(new_n1268), .A4(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1270), .A2(G2897), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1265), .A2(new_n1229), .ZN(new_n1281));
  INV_X1    g1081(.A(G384), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1265), .A2(G384), .A3(new_n1229), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1279), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1280), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1234), .B1(new_n1180), .B2(new_n1207), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1270), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1271), .A2(new_n1274), .A3(new_n1205), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1289), .B1(G378), .B2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1287), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1277), .A2(new_n1278), .A3(new_n1292), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n1295), .B2(new_n1268), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1259), .B1(new_n1293), .B2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(KEYINPUT63), .A3(new_n1268), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1257), .A2(KEYINPUT61), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT63), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1275), .A2(new_n1234), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1301), .B(new_n1289), .C1(new_n1231), .C2(new_n1234), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT123), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1280), .A2(new_n1286), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1280), .B2(new_n1286), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1300), .B1(new_n1302), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1268), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1302), .A2(new_n1308), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1298), .B(new_n1299), .C1(new_n1307), .C2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1297), .A2(new_n1310), .ZN(G405));
  NAND3_X1  g1111(.A1(new_n1257), .A2(KEYINPUT126), .A3(new_n1268), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT126), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1254), .B(new_n1256), .C1(new_n1313), .C2(new_n1308), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1268), .A2(KEYINPUT126), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(new_n1236), .A2(new_n1288), .A3(new_n1316), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1315), .B(new_n1317), .ZN(G402));
endmodule


