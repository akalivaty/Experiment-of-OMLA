//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n187));
  NOR2_X1   g001(.A1(G475), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G113), .B(G122), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G237), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G214), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT85), .ZN(new_n196));
  AOI21_X1  g010(.A(G143), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G214), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n198), .A2(G237), .A3(G953), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT85), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT88), .ZN(new_n202));
  AOI21_X1  g016(.A(G131), .B1(new_n199), .B2(G143), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n197), .A2(new_n200), .B1(G143), .B2(new_n199), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n202), .B1(new_n201), .B2(new_n203), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT89), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n208), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n199), .A2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n201), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G131), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT89), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n213), .A3(new_n214), .A4(new_n204), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT64), .A2(G146), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT64), .A2(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G125), .B(G140), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT19), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT73), .B(G125), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G140), .ZN(new_n223));
  NOR2_X1   g037(.A1(G125), .A2(G140), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n218), .B(new_n221), .C1(new_n226), .C2(new_n220), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT16), .ZN(new_n228));
  INV_X1    g042(.A(G140), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n222), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n224), .B1(new_n222), .B2(G140), .ZN(new_n231));
  OAI211_X1 g045(.A(G146), .B(new_n230), .C1(new_n231), .C2(new_n228), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n209), .A2(new_n215), .A3(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(KEYINPUT18), .A2(G131), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n212), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT86), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n212), .A2(KEYINPUT86), .A3(new_n235), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n212), .A2(new_n235), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n231), .A2(KEYINPUT87), .A3(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n218), .A2(new_n219), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT87), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n245), .B1(new_n226), .B2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n241), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n240), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n192), .B1(new_n234), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n226), .A2(KEYINPUT16), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n251), .A2(KEYINPUT74), .A3(G146), .A4(new_n230), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT74), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n232), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n230), .B1(new_n231), .B2(new_n228), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n246), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n212), .A2(KEYINPUT17), .A3(G131), .ZN(new_n257));
  AND4_X1   g071(.A1(new_n252), .A2(new_n254), .A3(new_n256), .A4(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT17), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n210), .A2(new_n213), .A3(new_n259), .A4(new_n204), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n258), .A2(new_n260), .B1(new_n240), .B2(new_n248), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n250), .A2(KEYINPUT90), .B1(new_n261), .B2(new_n192), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n234), .A2(new_n249), .ZN(new_n263));
  INV_X1    g077(.A(new_n192), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT90), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n189), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT20), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n187), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n263), .A2(KEYINPUT90), .A3(new_n264), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n261), .A2(new_n192), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n250), .A2(KEYINPUT90), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n188), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT92), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT20), .B1(new_n189), .B2(new_n277), .ZN(new_n278));
  OAI221_X1 g092(.A(new_n278), .B1(new_n277), .B2(new_n189), .C1(new_n273), .C2(new_n274), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n270), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  XOR2_X1   g094(.A(KEYINPUT93), .B(G475), .Z(new_n281));
  XNOR2_X1  g095(.A(new_n261), .B(new_n264), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(G902), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT99), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT97), .ZN(new_n285));
  INV_X1    g099(.A(G134), .ZN(new_n286));
  INV_X1    g100(.A(G143), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G128), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT13), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n289), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT95), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G128), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G143), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n288), .A2(KEYINPUT95), .A3(new_n289), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n290), .B1(new_n297), .B2(KEYINPUT96), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT96), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n293), .A2(new_n299), .A3(new_n295), .A4(new_n296), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n286), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(KEYINPUT65), .A2(G134), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(KEYINPUT65), .A2(G134), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n288), .A3(new_n295), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G122), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT94), .B1(new_n308), .B2(G116), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT94), .ZN(new_n310));
  INV_X1    g124(.A(G116), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n311), .A3(G122), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n308), .A2(G116), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G107), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G107), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n313), .A2(new_n318), .A3(new_n315), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n307), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n285), .B1(new_n301), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n296), .A2(new_n295), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT95), .B1(new_n288), .B2(new_n289), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT96), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n290), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n300), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G134), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(KEYINPUT97), .A3(new_n320), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n305), .B1(new_n288), .B2(new_n295), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n319), .B1(new_n307), .B2(new_n330), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n313), .A2(KEYINPUT14), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n316), .B1(new_n313), .B2(KEYINPUT14), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n318), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n322), .A2(new_n329), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT9), .B(G234), .ZN(new_n338));
  INV_X1    g152(.A(G217), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n338), .A2(new_n339), .A3(G953), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n328), .A2(new_n320), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n335), .B1(new_n343), .B2(new_n285), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n329), .A3(new_n340), .ZN(new_n345));
  AOI21_X1  g159(.A(G902), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G478), .ZN(new_n347));
  NOR2_X1   g161(.A1(KEYINPUT98), .A2(KEYINPUT15), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(KEYINPUT98), .A2(KEYINPUT15), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n347), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  AOI211_X1 g167(.A(G902), .B(new_n351), .C1(new_n342), .C2(new_n345), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n284), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G902), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n337), .A2(new_n341), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n340), .B1(new_n344), .B2(new_n329), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n351), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n346), .A2(new_n352), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(KEYINPUT99), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n194), .A2(G952), .ZN(new_n364));
  NAND2_X1  g178(.A1(G234), .A2(G237), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT21), .B(G898), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n365), .A2(G902), .A3(G953), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT100), .ZN(new_n371));
  AND4_X1   g185(.A1(new_n280), .A2(new_n283), .A3(new_n363), .A4(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT6), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n374), .B1(new_n191), .B2(G107), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n318), .A2(KEYINPUT3), .A3(G104), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT77), .B1(new_n318), .B2(G104), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT77), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n191), .A3(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G101), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT2), .B(G113), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(G116), .B(G119), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n311), .A2(G119), .ZN(new_n388));
  INV_X1    g202(.A(G119), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(G116), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n384), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G101), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n377), .A2(new_n393), .A3(new_n378), .A4(new_n380), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n378), .A2(new_n380), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n393), .B1(new_n396), .B2(new_n377), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n383), .B(new_n392), .C1(new_n395), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n386), .A2(KEYINPUT5), .ZN(new_n399));
  INV_X1    g213(.A(G113), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT5), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n400), .B1(new_n388), .B2(new_n401), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n399), .A2(new_n402), .B1(new_n385), .B2(new_n386), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT78), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n191), .A2(G107), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n318), .A2(G104), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n404), .B(G101), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(G104), .B(G107), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT78), .B1(new_n408), .B2(new_n393), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n403), .A2(new_n394), .A3(new_n407), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n398), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G110), .B(G122), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n373), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n397), .A2(new_n382), .B1(new_n387), .B2(new_n391), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n381), .A2(G101), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT4), .A3(new_n394), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n394), .A2(new_n407), .A3(new_n409), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n415), .A2(new_n417), .B1(new_n418), .B2(new_n403), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT80), .B1(new_n419), .B2(new_n412), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n398), .A2(KEYINPUT80), .A3(new_n410), .A4(new_n412), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n414), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n419), .A2(KEYINPUT6), .A3(new_n412), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT64), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n246), .ZN(new_n427));
  NAND2_X1  g241(.A1(KEYINPUT64), .A2(G146), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(G143), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT1), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n287), .A2(G146), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n429), .A2(new_n430), .A3(G128), .A4(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n222), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n216), .A2(new_n217), .A3(new_n287), .ZN(new_n436));
  OAI21_X1  g250(.A(G128), .B1(new_n436), .B2(new_n430), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n287), .B1(new_n216), .B2(new_n217), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n287), .A2(G146), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT69), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n294), .B1(new_n429), .B2(KEYINPUT1), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT64), .B(G146), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n439), .B1(new_n444), .B2(new_n287), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT69), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n435), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(KEYINPUT0), .A2(G128), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n429), .A2(new_n431), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT0), .B(G128), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n438), .B2(new_n440), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n222), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT81), .B(G224), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n194), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n446), .B1(new_n443), .B2(new_n445), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n430), .B1(new_n218), .B2(G143), .ZN(new_n458));
  OAI211_X1 g272(.A(KEYINPUT69), .B(new_n441), .C1(new_n458), .C2(new_n294), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n429), .A2(new_n431), .A3(new_n449), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n461), .B1(new_n445), .B2(new_n451), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n460), .A2(new_n435), .B1(new_n222), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(KEYINPUT81), .A2(G224), .ZN(new_n464));
  NOR2_X1   g278(.A1(KEYINPUT81), .A2(G224), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n194), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n456), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n423), .A2(new_n425), .A3(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n412), .B(KEYINPUT8), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n394), .A2(new_n407), .A3(new_n409), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n399), .A2(new_n402), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n387), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n471), .B1(new_n410), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n466), .A2(KEYINPUT7), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n454), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT82), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n466), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n455), .A2(KEYINPUT82), .A3(new_n194), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT7), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n462), .B2(new_n222), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n448), .A2(KEYINPUT83), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT83), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n434), .B1(new_n457), .B2(new_n459), .ZN(new_n486));
  INV_X1    g300(.A(new_n482), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n453), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n485), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n478), .A2(new_n490), .A3(KEYINPUT84), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n398), .A2(new_n410), .A3(new_n412), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT80), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n421), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT84), .B1(new_n478), .B2(new_n490), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n356), .B(new_n469), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G210), .B1(G237), .B2(G902), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n424), .B1(new_n495), .B2(new_n414), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n502), .B2(new_n468), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT84), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n484), .A2(new_n489), .ZN(new_n505));
  INV_X1    g319(.A(new_n477), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n410), .A2(new_n475), .ZN(new_n507));
  OAI22_X1  g321(.A1(new_n463), .A2(new_n506), .B1(new_n507), .B2(new_n471), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n504), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n495), .A3(new_n491), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n503), .A2(new_n510), .A3(new_n499), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n501), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(G214), .B1(G237), .B2(G902), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n372), .A2(new_n515), .ZN(new_n516));
  XOR2_X1   g330(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n517));
  NAND3_X1  g331(.A1(new_n193), .A2(new_n194), .A3(G210), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(G101), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT28), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n460), .A2(new_n432), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT11), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n524), .B1(new_n305), .B2(G137), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT66), .ZN(new_n526));
  NAND2_X1  g340(.A1(KEYINPUT11), .A2(G134), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n526), .B1(new_n527), .B2(G137), .ZN(new_n528));
  INV_X1    g342(.A(G137), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n529), .A2(KEYINPUT66), .A3(KEYINPUT11), .A4(G134), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OR2_X1    g345(.A1(KEYINPUT65), .A2(G134), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(G137), .A3(new_n302), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n525), .A2(new_n205), .A3(new_n531), .A4(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(G137), .B1(new_n532), .B2(new_n302), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT68), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT68), .B1(new_n529), .B2(G134), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n537), .B(G131), .C1(new_n535), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n523), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT67), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n531), .B(new_n533), .C1(new_n535), .C2(KEYINPUT11), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G131), .ZN(new_n545));
  AOI211_X1 g359(.A(new_n543), .B(new_n462), .C1(new_n545), .C2(new_n534), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n534), .ZN(new_n547));
  INV_X1    g361(.A(new_n462), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT67), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n542), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n392), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n548), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n392), .B(KEYINPUT70), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n542), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n522), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n522), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n521), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n542), .A2(KEYINPUT30), .A3(new_n552), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n540), .B1(new_n460), .B2(new_n432), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n552), .A2(new_n543), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n547), .A2(KEYINPUT67), .A3(new_n548), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n392), .B(new_n560), .C1(new_n564), .C2(KEYINPUT30), .ZN(new_n565));
  INV_X1    g379(.A(new_n521), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n555), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT29), .B1(new_n559), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n552), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n553), .B1(new_n569), .B2(new_n561), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT72), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n555), .A3(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(KEYINPUT72), .B(new_n553), .C1(new_n569), .C2(new_n561), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n557), .B1(new_n574), .B2(new_n522), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n521), .A2(KEYINPUT29), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n356), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G472), .B1(new_n568), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n566), .B1(new_n556), .B2(new_n558), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n555), .A2(new_n521), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n565), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT31), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT31), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n565), .A2(new_n583), .A3(new_n580), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n579), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT32), .ZN(new_n586));
  NOR2_X1   g400(.A1(G472), .A2(G902), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n586), .B1(new_n585), .B2(new_n587), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n578), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n523), .A2(KEYINPUT10), .A3(new_n418), .ZN(new_n591));
  INV_X1    g405(.A(new_n547), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n429), .A2(new_n431), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n294), .B1(new_n440), .B2(KEYINPUT1), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n432), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n418), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n417), .A2(new_n548), .A3(new_n383), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n591), .A2(new_n592), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n596), .B1(new_n523), .B2(new_n418), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(KEYINPUT12), .A3(new_n547), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT12), .B1(new_n601), .B2(new_n547), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n194), .A2(G227), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT76), .ZN(new_n607));
  XNOR2_X1  g421(.A(G110), .B(G140), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n609), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n600), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT79), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n591), .A2(new_n598), .A3(new_n599), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n547), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n600), .A2(KEYINPUT79), .A3(new_n611), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n610), .A2(new_n618), .A3(G469), .ZN(new_n619));
  INV_X1    g433(.A(G469), .ZN(new_n620));
  INV_X1    g434(.A(new_n604), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n612), .B1(new_n602), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n611), .B1(new_n616), .B2(new_n600), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n620), .B(new_n356), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(G469), .A2(G902), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n619), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(G221), .B1(new_n338), .B2(G902), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n339), .B1(G234), .B2(new_n356), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n252), .A2(new_n256), .A3(new_n254), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT23), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n389), .B2(G128), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n294), .A2(KEYINPUT23), .A3(G119), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n632), .B(new_n633), .C1(G119), .C2(new_n294), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT24), .B(G110), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(G119), .B(G128), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n634), .A2(G110), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n630), .A2(new_n639), .ZN(new_n640));
  OAI22_X1  g454(.A1(new_n634), .A2(G110), .B1(new_n636), .B2(new_n637), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n232), .A2(new_n243), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT22), .B(G137), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n640), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n645), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n630), .A2(new_n639), .ZN(new_n648));
  INV_X1    g462(.A(new_n642), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT75), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT25), .ZN(new_n652));
  AOI21_X1  g466(.A(G902), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n646), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n629), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n655), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n646), .A2(new_n650), .A3(new_n657), .A4(new_n653), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n646), .A2(new_n650), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n628), .A2(G902), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n656), .A2(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n626), .A2(new_n627), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n590), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n516), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n393), .ZN(G3));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n503), .A2(new_n510), .A3(new_n666), .A4(new_n499), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n667), .A2(new_n513), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n501), .A2(KEYINPUT101), .A3(new_n511), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n668), .A2(new_n669), .A3(KEYINPUT102), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT102), .B1(new_n668), .B2(new_n669), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n359), .A2(KEYINPUT103), .A3(new_n347), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(new_n346), .B2(G478), .ZN(new_n675));
  OAI21_X1  g489(.A(KEYINPUT33), .B1(new_n357), .B2(new_n358), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT33), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n342), .A2(new_n677), .A3(new_n345), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n347), .A2(G902), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n673), .A2(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n280), .B2(new_n283), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n672), .A2(new_n371), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(G472), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n585), .B2(new_n356), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n587), .B2(new_n585), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n687), .A2(new_n662), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT34), .B(G104), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G6));
  AND2_X1   g505(.A1(new_n355), .A2(new_n362), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n268), .A2(new_n269), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n270), .A2(new_n276), .A3(new_n693), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n692), .A2(new_n694), .A3(new_n283), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n672), .A2(new_n371), .A3(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n688), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT35), .B(G107), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G9));
  NAND2_X1  g514(.A1(new_n656), .A2(new_n658), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n640), .A2(new_n642), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n647), .A2(KEYINPUT36), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n660), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n626), .A2(new_n706), .A3(new_n627), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n687), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n516), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT37), .B(G110), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G12));
  XNOR2_X1  g525(.A(KEYINPUT104), .B(G900), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n712), .A2(new_n369), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n366), .ZN(new_n714));
  AND4_X1   g528(.A1(new_n283), .A2(new_n692), .A3(new_n694), .A4(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n672), .A2(new_n715), .A3(new_n590), .A4(new_n707), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G128), .ZN(G30));
  XOR2_X1   g531(.A(new_n512), .B(KEYINPUT38), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n714), .B(KEYINPUT39), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n626), .A2(new_n627), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n718), .B1(new_n720), .B2(KEYINPUT40), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(KEYINPUT40), .B2(new_n720), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n363), .B1(new_n280), .B2(new_n283), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n701), .A2(new_n705), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n513), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n574), .A2(new_n566), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n356), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n566), .B1(new_n565), .B2(new_n555), .ZN(new_n731));
  OAI21_X1  g545(.A(G472), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n588), .B2(new_n589), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT105), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n722), .A2(new_n727), .A3(new_n728), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G143), .ZN(G45));
  NAND2_X1  g551(.A1(new_n668), .A2(new_n669), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT102), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n668), .A2(new_n669), .A3(KEYINPUT102), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n590), .A2(new_n740), .A3(new_n741), .A4(new_n707), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n682), .A2(new_n714), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT107), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n626), .A2(new_n706), .A3(new_n627), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n585), .A2(new_n587), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT32), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n745), .B1(new_n749), .B2(new_n578), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n751));
  INV_X1    g565(.A(new_n714), .ZN(new_n752));
  AOI211_X1 g566(.A(new_n681), .B(new_n752), .C1(new_n280), .C2(new_n283), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n750), .A2(new_n751), .A3(new_n672), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n744), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G146), .ZN(G48));
  NOR2_X1   g570(.A1(new_n622), .A2(new_n623), .ZN(new_n757));
  OAI21_X1  g571(.A(G469), .B1(new_n757), .B2(G902), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n758), .A2(new_n627), .A3(new_n624), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n590), .A2(new_n661), .A3(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n683), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g575(.A(KEYINPUT41), .B(G113), .Z(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G15));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n764));
  INV_X1    g578(.A(new_n760), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n697), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT108), .B1(new_n696), .B2(new_n760), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g582(.A(KEYINPUT109), .B(G116), .Z(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(G18));
  NAND2_X1  g584(.A1(new_n672), .A2(new_n759), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n372), .A2(new_n590), .A3(new_n706), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(new_n389), .ZN(G21));
  NAND2_X1  g588(.A1(new_n672), .A2(new_n723), .ZN(new_n775));
  INV_X1    g589(.A(new_n587), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n582), .A2(new_n584), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n575), .A2(new_n566), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n686), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(new_n371), .A3(new_n661), .A4(new_n759), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n775), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n308), .ZN(G24));
  NOR3_X1   g597(.A1(new_n779), .A2(new_n686), .A3(new_n724), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n672), .A2(new_n753), .A3(new_n759), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G125), .ZN(G27));
  NAND2_X1  g600(.A1(new_n512), .A2(new_n513), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n626), .A2(new_n627), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n590), .A3(new_n661), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT111), .B1(KEYINPUT110), .B2(KEYINPUT42), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(KEYINPUT111), .B2(KEYINPUT42), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n753), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n792), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n790), .B2(new_n743), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n205), .ZN(G33));
  NAND2_X1  g613(.A1(new_n791), .A2(new_n715), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G134), .ZN(G36));
  NAND2_X1  g615(.A1(new_n280), .A2(new_n283), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT112), .B1(new_n802), .B2(new_n681), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT43), .Z(new_n804));
  OR2_X1    g618(.A1(new_n687), .A2(new_n724), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT44), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n787), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n806), .A2(new_n807), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n610), .A2(new_n618), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT45), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n620), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n812), .B2(new_n811), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n625), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT46), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n814), .A2(KEYINPUT46), .A3(new_n625), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n624), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n627), .ZN(new_n820));
  INV_X1    g634(.A(new_n719), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(KEYINPUT113), .B(G137), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n823), .B(new_n824), .ZN(G39));
  INV_X1    g639(.A(KEYINPUT47), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n820), .B(new_n826), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n743), .A2(new_n590), .A3(new_n661), .A4(new_n787), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n828), .A2(KEYINPUT114), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(KEYINPUT114), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G140), .ZN(G42));
  NAND2_X1  g646(.A1(new_n780), .A2(new_n661), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n804), .A2(new_n366), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n759), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n718), .A2(new_n513), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT50), .Z(new_n838));
  AND2_X1   g652(.A1(new_n758), .A2(new_n624), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n627), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n834), .B(new_n809), .C1(new_n827), .C2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n366), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n835), .A2(new_n787), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n734), .A2(new_n843), .A3(new_n661), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n681), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n845), .A2(new_n802), .A3(new_n846), .ZN(new_n847));
  NOR4_X1   g661(.A1(new_n804), .A2(new_n366), .A3(new_n835), .A4(new_n787), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n847), .B1(new_n848), .B2(new_n784), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n838), .A2(new_n842), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n848), .A2(new_n661), .A3(new_n590), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT48), .ZN(new_n854));
  INV_X1    g668(.A(new_n682), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n364), .B1(new_n845), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n771), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n856), .B1(new_n857), .B2(new_n834), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n852), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n850), .A2(new_n851), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n788), .A2(new_n706), .A3(new_n752), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n672), .A2(new_n723), .A3(new_n733), .A4(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n716), .A2(new_n785), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n865), .A2(KEYINPUT117), .A3(new_n755), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT117), .B1(new_n865), .B2(new_n755), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n744), .A2(new_n754), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n716), .A2(new_n785), .A3(new_n864), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n865), .A2(new_n755), .A3(KEYINPUT117), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT52), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n862), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n868), .B1(new_n866), .B2(new_n867), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n873), .A2(KEYINPUT52), .A3(new_n874), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n878), .A3(KEYINPUT118), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n802), .B1(new_n360), .B2(new_n361), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(new_n682), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n687), .A2(new_n515), .A3(new_n371), .A4(new_n662), .ZN(new_n883));
  OAI22_X1  g697(.A1(new_n882), .A2(new_n883), .B1(new_n775), .B2(new_n781), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n683), .A2(new_n760), .B1(new_n771), .B2(new_n772), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n516), .B1(new_n663), .B2(new_n708), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n768), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n753), .A2(new_n784), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n590), .A2(new_n706), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n353), .A2(new_n354), .A3(new_n752), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n694), .A2(new_n283), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n890), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n789), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(new_n797), .A3(new_n795), .A4(new_n800), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n880), .B1(new_n889), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n896), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n898), .A2(KEYINPUT116), .A3(new_n768), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n876), .A2(new_n879), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT53), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n868), .B1(new_n865), .B2(new_n755), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n875), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT53), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n901), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n903), .A2(KEYINPUT54), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n902), .A2(new_n906), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n910));
  INV_X1    g724(.A(new_n905), .ZN(new_n911));
  INV_X1    g725(.A(new_n889), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(KEYINPUT53), .A3(new_n898), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n909), .A2(new_n910), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n861), .A2(new_n908), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(G952), .B2(G953), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT49), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n839), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n661), .A2(new_n513), .A3(new_n627), .ZN(new_n920));
  NOR4_X1   g734(.A1(new_n919), .A2(new_n802), .A3(new_n681), .A4(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT115), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n718), .B1(new_n918), .B2(new_n839), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n734), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n917), .A2(new_n924), .ZN(G75));
  NOR2_X1   g739(.A1(new_n194), .A2(G952), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n356), .B1(new_n909), .B2(new_n914), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT56), .B1(new_n928), .B2(G210), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n502), .B(new_n468), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT55), .Z(new_n931));
  OAI21_X1  g745(.A(new_n927), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n929), .A2(new_n931), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT119), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n929), .A2(KEYINPUT119), .A3(new_n931), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(G51));
  NAND2_X1  g751(.A1(new_n877), .A2(new_n878), .ZN(new_n938));
  AOI22_X1  g752(.A1(new_n938), .A2(new_n862), .B1(new_n897), .B2(new_n900), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT53), .B1(new_n939), .B2(new_n879), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n911), .A2(new_n913), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT54), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n942), .A2(KEYINPUT120), .A3(new_n915), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n944), .B(KEYINPUT54), .C1(new_n940), .C2(new_n941), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n625), .B(KEYINPUT57), .Z(new_n946));
  NAND3_X1  g760(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n757), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n928), .B(new_n813), .C1(new_n812), .C2(new_n811), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n926), .B1(new_n949), .B2(new_n950), .ZN(G54));
  NAND3_X1  g765(.A1(new_n928), .A2(KEYINPUT58), .A3(G475), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n273), .A2(new_n274), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n927), .B1(new_n952), .B2(new_n954), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n953), .B1(new_n952), .B2(new_n954), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(G60));
  NAND2_X1  g772(.A1(G478), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT59), .Z(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n908), .B2(new_n915), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n927), .B1(new_n961), .B2(new_n679), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n943), .A2(new_n945), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n960), .B1(new_n676), .B2(new_n678), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(G63));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT60), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n940), .B2(new_n941), .ZN(new_n969));
  INV_X1    g783(.A(new_n659), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n926), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT122), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT61), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n704), .B(new_n968), .C1(new_n940), .C2(new_n941), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n971), .B(new_n974), .C1(new_n972), .C2(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(G66));
  INV_X1    g792(.A(new_n455), .ZN(new_n979));
  OAI21_X1  g793(.A(G953), .B1(new_n979), .B2(new_n367), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n912), .B2(G953), .ZN(new_n981));
  INV_X1    g795(.A(new_n502), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(G898), .B2(new_n194), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n981), .B(new_n983), .ZN(G69));
  OAI21_X1  g798(.A(new_n560), .B1(new_n564), .B2(KEYINPUT30), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT123), .Z(new_n986));
  OAI21_X1  g800(.A(new_n221), .B1(new_n226), .B2(new_n220), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n986), .B(new_n987), .Z(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(G900), .B2(G953), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n823), .A2(new_n831), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n755), .A2(new_n716), .A3(new_n785), .ZN(new_n993));
  INV_X1    g807(.A(new_n800), .ZN(new_n994));
  INV_X1    g808(.A(new_n822), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT125), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n672), .A2(new_n661), .A3(new_n590), .A4(new_n723), .ZN(new_n997));
  OR3_X1    g811(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n996), .B1(new_n995), .B2(new_n997), .ZN(new_n999));
  AOI211_X1 g813(.A(new_n798), .B(new_n994), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n992), .A2(new_n993), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n991), .B1(new_n1001), .B2(new_n194), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n993), .A2(new_n736), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n882), .A2(new_n790), .A3(new_n821), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT124), .Z(new_n1006));
  OR2_X1    g820(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n992), .A2(new_n1004), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n988), .B1(new_n1008), .B2(new_n194), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n1010));
  OAI22_X1  g824(.A1(new_n1002), .A2(new_n1009), .B1(KEYINPUT126), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(KEYINPUT126), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1011), .B(new_n1012), .ZN(G72));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n1008), .B2(new_n889), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n731), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1015), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1018), .B1(new_n1001), .B2(new_n912), .ZN(new_n1019));
  OAI211_X1 g833(.A(new_n1017), .B(new_n927), .C1(new_n567), .C2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n567), .A2(new_n1015), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1021), .A2(new_n731), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n903), .A2(new_n907), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT127), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1020), .B1(new_n1025), .B2(new_n1026), .ZN(G57));
endmodule


