//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT64), .Z(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AND2_X1   g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G20), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT65), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n202), .A2(KEYINPUT66), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(KEYINPUT66), .ZN(new_n214));
  AND3_X1   g0014(.A1(new_n213), .A2(G50), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n209), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT67), .B(G244), .Z(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G77), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G116), .A2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT68), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n205), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n216), .B1(KEYINPUT1), .B2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT69), .ZN(new_n237));
  XOR2_X1   g0037(.A(G58), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G351));
  XNOR2_X1  g0044(.A(KEYINPUT3), .B(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G1698), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n245), .A2(G222), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n245), .A2(G223), .A3(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(G77), .ZN(new_n249));
  OAI211_X1 g0049(.A(new_n247), .B(new_n248), .C1(new_n249), .C2(new_n245), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n251), .B1(G33), .B2(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(new_n258), .A3(G274), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n252), .A2(new_n256), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n260), .B1(G226), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n253), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G190), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n265), .B1(G200), .B2(new_n263), .ZN(new_n266));
  INV_X1    g0066(.A(G13), .ZN(new_n267));
  INV_X1    g0067(.A(G20), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n267), .A2(new_n268), .A3(G1), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(KEYINPUT70), .A3(new_n251), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(KEYINPUT70), .B1(new_n271), .B2(new_n251), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OR3_X1    g0075(.A1(new_n268), .A2(KEYINPUT71), .A3(G1), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT71), .B1(new_n268), .B2(G1), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G50), .ZN(new_n279));
  OAI22_X1  g0079(.A1(new_n275), .A2(new_n279), .B1(G50), .B2(new_n270), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT72), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n273), .A2(new_n274), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n268), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(G150), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n284), .A2(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G50), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n268), .B1(new_n201), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n283), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n282), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n266), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT76), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n245), .A2(G232), .A3(G1698), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n245), .A2(G226), .A3(new_n246), .ZN(new_n300));
  INV_X1    g0100(.A(G33), .ZN(new_n301));
  INV_X1    g0101(.A(G97), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n299), .B(new_n300), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n252), .ZN(new_n304));
  INV_X1    g0104(.A(G1), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(G41), .B2(G45), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n258), .A2(G238), .A3(new_n306), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n259), .A2(new_n307), .A3(KEYINPUT74), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT74), .B1(new_n259), .B2(new_n307), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n304), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT13), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT13), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n304), .B(new_n312), .C1(new_n309), .C2(new_n308), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(G190), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n274), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n269), .B1(new_n315), .B2(new_n272), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(G68), .A3(new_n278), .ZN(new_n317));
  INV_X1    g0117(.A(G68), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n269), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n319), .B(KEYINPUT12), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n285), .A2(new_n249), .B1(new_n268), .B2(G68), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n321), .A2(KEYINPUT75), .B1(new_n290), .B2(new_n288), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n321), .A2(KEYINPUT75), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n283), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT11), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n317), .B(new_n320), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n324), .A2(new_n325), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n314), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n311), .B2(new_n313), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n298), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n331), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n333), .A2(KEYINPUT76), .A3(new_n328), .A4(new_n314), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n311), .A2(new_n313), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G169), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT14), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(G179), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT14), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n336), .A2(new_n341), .A3(G169), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n328), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n293), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n263), .A2(new_n338), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(G179), .B2(new_n263), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n245), .A2(G232), .A3(new_n246), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n245), .A2(G238), .A3(G1698), .ZN(new_n351));
  INV_X1    g0151(.A(G107), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n350), .B(new_n351), .C1(new_n352), .C2(new_n245), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n252), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n260), .B1(new_n217), .B2(new_n261), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G179), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G20), .A2(G77), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n359), .B1(new_n284), .B2(new_n288), .C1(new_n285), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n283), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n316), .A2(G77), .A3(new_n278), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n269), .A2(new_n249), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n358), .B(new_n365), .C1(G169), .C2(new_n356), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n349), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT73), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n330), .B1(new_n354), .B2(new_n355), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n365), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n365), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n371), .A2(KEYINPUT73), .B1(G190), .B2(new_n356), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n367), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n297), .A2(new_n335), .A3(new_n345), .A4(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT18), .ZN(new_n375));
  INV_X1    g0175(.A(G58), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(new_n318), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n377), .A2(new_n201), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(G20), .B1(G159), .B2(new_n287), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n301), .A2(KEYINPUT3), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT3), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G33), .ZN(new_n383));
  AOI211_X1 g0183(.A(new_n380), .B(G20), .C1(new_n381), .C2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n382), .A2(G33), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n301), .A2(KEYINPUT3), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT77), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT77), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n381), .A2(new_n383), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n268), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n384), .B1(new_n390), .B2(new_n380), .ZN(new_n391));
  OAI211_X1 g0191(.A(KEYINPUT16), .B(new_n379), .C1(new_n391), .C2(new_n318), .ZN(new_n392));
  XOR2_X1   g0192(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n393));
  INV_X1    g0193(.A(new_n379), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n380), .B1(new_n245), .B2(G20), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n381), .A2(new_n383), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(KEYINPUT7), .A3(new_n268), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n318), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n393), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n392), .A2(new_n283), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n284), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n278), .A2(new_n401), .ZN(new_n402));
  OAI22_X1  g0202(.A1(new_n275), .A2(new_n402), .B1(new_n270), .B2(new_n401), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT79), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT79), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n405), .B1(new_n270), .B2(new_n401), .C1(new_n275), .C2(new_n402), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n381), .A2(new_n383), .A3(G226), .A4(G1698), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n381), .A2(new_n383), .A3(G223), .A4(new_n246), .ZN(new_n410));
  INV_X1    g0210(.A(G87), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n409), .B(new_n410), .C1(new_n301), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n252), .ZN(new_n413));
  INV_X1    g0213(.A(G274), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n210), .B2(new_n257), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n261), .A2(G232), .B1(new_n256), .B2(new_n415), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n413), .A2(new_n416), .A3(G179), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n338), .B1(new_n413), .B2(new_n416), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n375), .B1(new_n408), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n283), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT7), .B1(new_n396), .B2(new_n268), .ZN(new_n423));
  OAI21_X1  g0223(.A(G68), .B1(new_n423), .B2(new_n384), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n379), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n422), .B1(new_n425), .B2(new_n393), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(new_n392), .B1(new_n404), .B2(new_n406), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n427), .A2(KEYINPUT18), .A3(new_n419), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT80), .B1(new_n421), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n413), .A2(new_n416), .A3(new_n264), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n413), .A2(new_n416), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(G200), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n400), .A2(new_n407), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT81), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT81), .B1(new_n427), .B2(new_n432), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT17), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT17), .B1(new_n427), .B2(new_n432), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n408), .A2(new_n375), .A3(new_n420), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT18), .B1(new_n427), .B2(new_n419), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT80), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n429), .A2(new_n437), .A3(new_n439), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n258), .A2(G274), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n255), .A2(G1), .ZN(new_n446));
  AND2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT5), .B(G41), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n252), .B1(new_n446), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n450), .B1(G270), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n245), .A2(G264), .A3(G1698), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n245), .A2(G257), .A3(new_n246), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n396), .A2(G303), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n252), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(KEYINPUT21), .A3(G169), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT87), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n305), .A2(G33), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n270), .B(new_n462), .C1(new_n273), .C2(new_n274), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n316), .A2(KEYINPUT87), .A3(G116), .A4(new_n462), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(new_n268), .C1(G33), .C2(new_n302), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n271), .A2(new_n251), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n464), .A2(G20), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n470), .A2(KEYINPUT88), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT88), .B1(new_n470), .B2(new_n471), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT20), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(KEYINPUT20), .B(new_n469), .C1(new_n472), .C2(new_n473), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n476), .A2(new_n477), .B1(new_n464), .B2(new_n269), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n460), .B1(new_n467), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n467), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n453), .A2(new_n458), .A3(G179), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n479), .A2(KEYINPUT89), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n459), .A2(G169), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT21), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT89), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n478), .A2(new_n467), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(new_n460), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n459), .A2(G200), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n489), .B(new_n491), .C1(new_n264), .C2(new_n459), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n483), .A2(new_n487), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n449), .A2(G257), .A3(new_n258), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n415), .A2(new_n446), .A3(new_n451), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n381), .A2(new_n383), .A3(G244), .A4(new_n246), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n245), .A2(KEYINPUT4), .A3(G244), .A4(new_n246), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n245), .A2(G250), .A3(G1698), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n468), .A4(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n496), .B1(new_n502), .B2(new_n252), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n503), .A2(KEYINPUT82), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(KEYINPUT82), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G190), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n287), .A2(G77), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT6), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n509), .A2(new_n302), .A3(G107), .ZN(new_n510));
  XNOR2_X1  g0310(.A(G97), .B(G107), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(new_n509), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n508), .B1(new_n512), .B2(new_n268), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n352), .B1(new_n395), .B2(new_n397), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n283), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n463), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G97), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n269), .A2(new_n302), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n502), .A2(new_n252), .ZN(new_n520));
  INV_X1    g0320(.A(new_n496), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n519), .B1(G200), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n503), .A2(new_n357), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n338), .B1(new_n504), .B2(new_n505), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n507), .A2(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT22), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n268), .A2(KEYINPUT90), .A3(G87), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n396), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n529), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n245), .A2(new_n531), .A3(KEYINPUT22), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G116), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(G20), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT23), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n268), .B2(G107), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n352), .A2(KEYINPUT23), .A3(G20), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n530), .A2(new_n532), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT24), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n530), .A2(new_n532), .A3(new_n538), .A4(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n422), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n305), .A2(new_n352), .A3(G13), .A4(G20), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT25), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g0346(.A(new_n546), .B(KEYINPUT91), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n544), .A2(new_n545), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT92), .ZN(new_n549));
  XNOR2_X1  g0349(.A(new_n548), .B(new_n549), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n547), .A2(new_n550), .B1(new_n352), .B2(new_n463), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT93), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n452), .A2(new_n553), .A3(G264), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n449), .A2(G264), .A3(new_n258), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT93), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n245), .A2(G257), .A3(G1698), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n245), .A2(G250), .A3(new_n246), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G294), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n554), .A2(new_n556), .B1(new_n560), .B2(new_n252), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n561), .A2(new_n264), .A3(new_n495), .ZN(new_n562));
  AOI21_X1  g0362(.A(G200), .B1(new_n561), .B2(new_n495), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n552), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n381), .A2(new_n383), .A3(G238), .A4(new_n246), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT84), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT84), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n245), .A2(new_n567), .A3(G238), .A4(new_n246), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n245), .A2(G244), .A3(G1698), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n566), .A2(new_n568), .A3(new_n533), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n252), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n305), .A2(G45), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G250), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n252), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT83), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n415), .B2(new_n446), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n415), .A2(new_n575), .A3(new_n446), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n574), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n571), .A2(new_n579), .A3(new_n264), .ZN(new_n580));
  AND4_X1   g0380(.A1(new_n575), .A2(new_n258), .A3(G274), .A4(new_n446), .ZN(new_n581));
  OAI22_X1  g0381(.A1(new_n576), .A2(new_n581), .B1(new_n252), .B2(new_n573), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n252), .B2(new_n570), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n580), .B1(new_n583), .B2(G200), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n411), .A2(new_n302), .A3(new_n352), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT85), .ZN(new_n586));
  NOR2_X1   g0386(.A1(G87), .A2(G97), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT85), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(new_n352), .ZN(new_n589));
  NAND3_X1  g0389(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n586), .A2(new_n589), .B1(new_n268), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n268), .A2(G33), .A3(G97), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT19), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n318), .A2(G20), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n594), .B1(new_n396), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT86), .B1(new_n591), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n590), .A2(new_n268), .ZN(new_n599));
  INV_X1    g0399(.A(new_n589), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n588), .B1(new_n587), .B2(new_n352), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT86), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n245), .A2(new_n595), .B1(new_n593), .B2(new_n592), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n598), .A2(new_n605), .A3(new_n283), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n360), .A2(new_n269), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n516), .A2(G87), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n584), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n571), .A2(new_n579), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n338), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n463), .A2(new_n360), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n606), .A2(new_n613), .A3(new_n607), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n571), .A2(new_n579), .A3(new_n357), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n564), .A2(new_n610), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n561), .A2(new_n495), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(G169), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n618), .A2(G179), .B1(new_n543), .B2(new_n551), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n527), .A2(new_n617), .A3(new_n624), .ZN(new_n625));
  NOR4_X1   g0425(.A1(new_n374), .A2(new_n444), .A3(new_n493), .A4(new_n625), .ZN(G372));
  NOR2_X1   g0426(.A1(new_n374), .A2(new_n444), .ZN(new_n627));
  INV_X1    g0427(.A(new_n616), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n610), .A2(new_n526), .A3(new_n525), .A4(new_n616), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n571), .A2(new_n579), .A3(new_n357), .ZN(new_n632));
  AOI21_X1  g0432(.A(G169), .B1(new_n571), .B2(new_n579), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n634), .A2(new_n614), .B1(new_n584), .B2(new_n609), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n519), .A2(new_n524), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT82), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n522), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n503), .A2(KEYINPUT82), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n636), .B1(new_n640), .B2(new_n338), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n635), .A2(new_n641), .A3(KEYINPUT26), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n628), .B1(new_n631), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n480), .A2(new_n482), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n480), .A2(new_n485), .A3(KEYINPUT89), .A4(KEYINPUT21), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n490), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n484), .B1(new_n467), .B2(new_n478), .ZN(new_n647));
  OAI22_X1  g0447(.A1(new_n620), .A2(new_n622), .B1(new_n647), .B2(KEYINPUT21), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n527), .B(new_n617), .C1(new_n646), .C2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n627), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n349), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n421), .A2(new_n428), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n329), .A2(new_n331), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n366), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n343), .A2(new_n344), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n437), .A2(new_n439), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n652), .B1(new_n659), .B2(new_n297), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n651), .A2(new_n660), .ZN(G369));
  NAND3_X1  g0461(.A1(new_n305), .A2(new_n268), .A3(G13), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n489), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n646), .B2(new_n486), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n493), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT94), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n552), .A2(new_n668), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT95), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n676), .A2(new_n564), .A3(new_n624), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n624), .A2(new_n668), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n490), .A2(new_n644), .A3(new_n645), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n667), .B1(new_n681), .B2(new_n487), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n623), .A2(new_n621), .A3(new_n668), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n680), .A2(new_n685), .ZN(G399));
  NAND3_X1  g0486(.A1(new_n586), .A2(new_n464), .A3(new_n589), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n206), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n691), .A3(G1), .ZN(new_n692));
  INV_X1    g0492(.A(new_n215), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(new_n691), .ZN(new_n694));
  XOR2_X1   g0494(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n695));
  XNOR2_X1  g0495(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n629), .A2(new_n630), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT26), .B1(new_n635), .B2(new_n641), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n616), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT99), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT100), .B1(new_n646), .B2(new_n648), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n486), .B1(new_n621), .B2(new_n623), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT100), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(new_n490), .A4(new_n483), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n526), .A2(new_n525), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n523), .B1(new_n264), .B2(new_n640), .ZN(new_n707));
  AND4_X1   g0507(.A1(new_n706), .A2(new_n707), .A3(new_n564), .A4(new_n635), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n702), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT99), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n643), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n701), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n697), .B1(new_n712), .B2(new_n668), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n667), .B1(new_n643), .B2(new_n649), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(KEYINPUT29), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n481), .A2(KEYINPUT97), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT97), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n453), .A2(new_n458), .A3(new_n720), .A4(G179), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n719), .A2(new_n561), .A3(new_n583), .A4(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n718), .B1(new_n722), .B2(new_n640), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n583), .A2(new_n503), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n357), .A3(new_n459), .A4(new_n618), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n638), .A2(KEYINPUT30), .A3(new_n639), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n722), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n667), .B1(new_n724), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n723), .B(new_n726), .C1(new_n722), .C2(new_n727), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT31), .B1(new_n732), .B2(new_n667), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT98), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n729), .A2(new_n730), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT98), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n493), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n739), .A2(new_n708), .A3(new_n624), .A4(new_n668), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n734), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G330), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n717), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n696), .B1(new_n744), .B2(G1), .ZN(G364));
  NOR2_X1   g0545(.A1(new_n267), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n305), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n690), .A2(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n264), .A2(G179), .A3(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n268), .ZN(new_n751));
  INV_X1    g0551(.A(G294), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n268), .A2(new_n357), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G317), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n758), .A2(KEYINPUT33), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(KEYINPUT33), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n757), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n755), .A2(new_n264), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n753), .B(new_n761), .C1(G326), .C2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n754), .A2(G190), .A3(new_n330), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n268), .A2(G179), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G190), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n765), .A2(G322), .B1(new_n769), .B2(G329), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n754), .A2(new_n767), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n770), .B(new_n396), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G283), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n766), .A2(new_n264), .A3(G200), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n766), .A2(G190), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(G303), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n757), .A2(new_n318), .B1(new_n775), .B2(new_n352), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n245), .B1(new_n772), .B2(new_n249), .C1(new_n376), .C2(new_n764), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n751), .A2(new_n302), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n776), .A2(new_n411), .ZN(new_n783));
  NOR4_X1   g0583(.A1(new_n780), .A2(new_n781), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n762), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT32), .ZN(new_n786));
  XNOR2_X1  g0586(.A(KEYINPUT102), .B(G159), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n768), .A2(new_n787), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n785), .A2(new_n290), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(new_n786), .B2(new_n788), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n763), .A2(new_n779), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n251), .B1(G20), .B2(new_n338), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n749), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n689), .A2(new_n396), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n795), .A2(G355), .B1(new_n464), .B2(new_n689), .ZN(new_n796));
  AND3_X1   g0596(.A1(new_n381), .A2(new_n383), .A3(new_n388), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n388), .B1(new_n381), .B2(new_n383), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n689), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(new_n255), .B2(new_n215), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT101), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n255), .B2(new_n239), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n803), .A2(new_n804), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n796), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n792), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n794), .B1(new_n808), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n811), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n671), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n749), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n671), .B2(G330), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n815), .B1(new_n674), .B2(new_n817), .ZN(G396));
  NAND2_X1  g0618(.A1(new_n656), .A2(new_n668), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n372), .A2(new_n370), .B1(new_n365), .B2(new_n667), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n820), .B2(new_n656), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n714), .B(new_n822), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n742), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n749), .B1(new_n742), .B2(new_n823), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n792), .A2(new_n809), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n749), .B1(G77), .B2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT103), .Z(new_n830));
  NOR2_X1   g0630(.A1(new_n822), .A2(new_n810), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n757), .A2(new_n774), .B1(new_n776), .B2(new_n352), .ZN(new_n832));
  INV_X1    g0632(.A(new_n775), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(G87), .B2(new_n833), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n764), .A2(new_n752), .B1(new_n768), .B2(new_n771), .ZN(new_n835));
  INV_X1    g0635(.A(new_n772), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n245), .B(new_n835), .C1(G116), .C2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n782), .B1(G303), .B2(new_n762), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n834), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  XOR2_X1   g0639(.A(KEYINPUT104), .B(G143), .Z(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n787), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n765), .A2(new_n841), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(G137), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n843), .B1(new_n785), .B2(new_n844), .C1(new_n286), .C2(new_n757), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT105), .Z(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(KEYINPUT34), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n775), .A2(new_n318), .ZN(new_n848));
  INV_X1    g0648(.A(new_n751), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(G58), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n290), .B2(new_n776), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n799), .B(new_n851), .C1(G132), .C2(new_n769), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n846), .A2(KEYINPUT34), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n839), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n830), .B(new_n831), .C1(new_n792), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n826), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  NOR2_X1   g0658(.A1(new_n746), .A2(new_n305), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT40), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n740), .A2(new_n735), .A3(new_n737), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n335), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n344), .A2(new_n667), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OR3_X1    g0666(.A1(new_n328), .A2(KEYINPUT107), .A3(new_n668), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n864), .A2(KEYINPUT107), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n345), .A2(new_n655), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n861), .A2(new_n870), .A3(new_n822), .ZN(new_n871));
  INV_X1    g0671(.A(new_n403), .ZN(new_n872));
  INV_X1    g0672(.A(new_n393), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT7), .B1(new_n799), .B2(new_n268), .ZN(new_n874));
  OAI21_X1  g0674(.A(G68), .B1(new_n874), .B2(new_n384), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n875), .B2(new_n379), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n392), .A2(new_n283), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n665), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n444), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n433), .A2(new_n434), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n427), .A2(KEYINPUT81), .A3(new_n432), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n419), .A2(new_n665), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT37), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n408), .B1(new_n420), .B2(new_n879), .ZN(new_n889));
  XNOR2_X1  g0689(.A(KEYINPUT108), .B(KEYINPUT37), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n889), .A2(new_n883), .A3(new_n884), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n882), .A2(KEYINPUT38), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n408), .A2(new_n879), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n438), .B1(new_n885), .B2(KEYINPUT17), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n653), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n889), .A2(new_n433), .ZN(new_n898));
  INV_X1    g0698(.A(new_n890), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n891), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n894), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n893), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n860), .B1(new_n871), .B2(new_n904), .ZN(new_n905));
  AOI221_X4 g0705(.A(new_n894), .B1(new_n888), .B2(new_n891), .C1(new_n444), .C2(new_n881), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n882), .B2(new_n892), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n861), .A2(new_n870), .A3(new_n860), .A4(new_n822), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT109), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n627), .A2(new_n861), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(G330), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  INV_X1    g0717(.A(new_n895), .ZN(new_n918));
  INV_X1    g0718(.A(new_n653), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n918), .B1(new_n658), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n920), .B2(new_n901), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n917), .B1(new_n906), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n442), .B1(new_n440), .B2(new_n441), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n880), .B1(new_n925), .B2(new_n896), .ZN(new_n926));
  INV_X1    g0726(.A(new_n892), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n894), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(KEYINPUT39), .A3(new_n893), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n343), .A2(new_n344), .A3(new_n668), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n667), .B(new_n821), .C1(new_n643), .C2(new_n649), .ZN(new_n933));
  INV_X1    g0733(.A(new_n819), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n870), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n908), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n653), .A2(new_n879), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n932), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n627), .B1(new_n713), .B2(new_n716), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n660), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n938), .B(new_n940), .Z(new_n941));
  AOI21_X1  g0741(.A(new_n859), .B1(new_n916), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n941), .B2(new_n916), .ZN(new_n943));
  INV_X1    g0743(.A(new_n512), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n944), .A2(KEYINPUT35), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(KEYINPUT35), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n945), .A2(G116), .A3(new_n212), .A4(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT36), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n693), .A2(new_n249), .A3(new_n377), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n318), .A2(G50), .ZN(new_n950));
  OAI211_X1 g0750(.A(G1), .B(new_n267), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT106), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n943), .A2(new_n948), .A3(new_n952), .ZN(G367));
  OAI221_X1 g0753(.A(new_n812), .B1(new_n206), .B2(new_n360), .C1(new_n802), .C2(new_n234), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n954), .A2(new_n749), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n609), .A2(new_n668), .ZN(new_n956));
  MUX2_X1   g0756(.A(new_n635), .B(new_n628), .S(new_n956), .Z(new_n957));
  OAI22_X1  g0757(.A1(new_n757), .A2(new_n752), .B1(new_n775), .B2(new_n302), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(G311), .B2(new_n762), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n764), .A2(new_n777), .B1(new_n772), .B2(new_n774), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G317), .B2(new_n769), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n800), .B1(G107), .B2(new_n849), .ZN(new_n962));
  INV_X1    g0762(.A(new_n776), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(G116), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT46), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n959), .A2(new_n961), .A3(new_n962), .A4(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n762), .A2(new_n841), .B1(new_n765), .B2(G150), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n318), .B2(new_n751), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT111), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n245), .B1(new_n768), .B2(new_n844), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G50), .B2(new_n836), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n776), .A2(new_n376), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n775), .A2(new_n249), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(new_n756), .C2(new_n842), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n969), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n968), .A2(KEYINPUT111), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n966), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT47), .Z(new_n978));
  OAI221_X1 g0778(.A(new_n955), .B1(new_n957), .B2(new_n814), .C1(new_n978), .C2(new_n793), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT44), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n707), .A2(new_n706), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n519), .A2(new_n667), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n981), .A2(new_n982), .B1(new_n706), .B2(new_n668), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n685), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n980), .B1(new_n685), .B2(new_n983), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n685), .A2(new_n983), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n685), .A2(KEYINPUT45), .A3(new_n983), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n680), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n985), .A2(new_n984), .B1(new_n989), .B2(new_n990), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n680), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n683), .B1(new_n679), .B2(new_n682), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n673), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n673), .A2(new_n998), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n744), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n690), .B(KEYINPUT41), .Z(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n748), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n677), .A2(new_n682), .A3(new_n983), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1006), .A2(KEYINPUT42), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n624), .B1(new_n507), .B2(new_n523), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n668), .B1(new_n1008), .B2(new_n641), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1006), .A2(KEYINPUT42), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n957), .B(KEYINPUT43), .ZN(new_n1017));
  AND3_X1   g0817(.A1(new_n1012), .A2(new_n1017), .A3(new_n1013), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n993), .B(new_n983), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1018), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n993), .A2(new_n983), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(new_n1015), .C2(new_n1014), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n979), .B1(new_n1005), .B2(new_n1023), .ZN(G387));
  NOR2_X1   g0824(.A1(new_n1001), .A2(new_n747), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT112), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1001), .A2(new_n743), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1001), .A2(new_n743), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n690), .B(KEYINPUT115), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n801), .B1(new_n231), .B2(new_n255), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n795), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1032), .B1(new_n688), .B2(new_n1033), .ZN(new_n1034));
  OR3_X1    g0834(.A1(new_n284), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1035));
  OAI21_X1  g0835(.A(KEYINPUT50), .B1(new_n284), .B2(G50), .ZN(new_n1036));
  AOI21_X1  g0836(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n688), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1034), .A2(new_n1038), .B1(new_n352), .B2(new_n689), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n812), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n749), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n776), .A2(new_n249), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n800), .B1(new_n286), .B2(new_n768), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(G97), .C2(new_n833), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT113), .Z(new_n1045));
  NOR2_X1   g0845(.A1(new_n751), .A2(new_n360), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n765), .A2(G50), .B1(new_n836), .B2(G68), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n284), .B2(new_n757), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1046), .B(new_n1048), .C1(G159), .C2(new_n762), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n764), .A2(new_n758), .B1(new_n772), .B2(new_n777), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT114), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(KEYINPUT114), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G311), .A2(new_n756), .B1(new_n762), .B2(G322), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT48), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n751), .A2(new_n774), .B1(new_n776), .B2(new_n752), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(KEYINPUT49), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n800), .B1(G326), .B2(new_n769), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n464), .C2(new_n775), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT49), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1050), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1041), .B1(new_n1064), .B2(new_n792), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n679), .B2(new_n814), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1026), .A2(new_n1031), .A3(new_n1066), .ZN(G393));
  NOR2_X1   g0867(.A1(new_n983), .A2(new_n814), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n812), .B1(new_n302), .B2(new_n206), .C1(new_n802), .C2(new_n243), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n751), .A2(new_n249), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n290), .B2(new_n757), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n840), .A2(new_n768), .B1(new_n772), .B2(new_n284), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n318), .A2(new_n776), .B1(new_n775), .B2(new_n411), .ZN(new_n1074));
  NOR4_X1   g0874(.A1(new_n1072), .A2(new_n799), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(G159), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n785), .A2(new_n286), .B1(new_n1076), .B2(new_n764), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT51), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n785), .A2(new_n758), .B1(new_n771), .B2(new_n764), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT52), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n757), .A2(new_n777), .B1(new_n464), .B2(new_n751), .ZN(new_n1081));
  INV_X1    g0881(.A(G322), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n396), .B1(new_n768), .B2(new_n1082), .C1(new_n752), .C2(new_n772), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n352), .A2(new_n775), .B1(new_n776), .B2(new_n774), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n1081), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1075), .A2(new_n1078), .B1(new_n1080), .B2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n749), .B(new_n1069), .C1(new_n1086), .C2(new_n793), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1068), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1030), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n997), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n1027), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n992), .A2(new_n993), .A3(KEYINPUT116), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n994), .A2(KEYINPUT116), .A3(new_n996), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n1028), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1088), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT117), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n994), .A2(KEYINPUT116), .A3(new_n996), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1097), .B1(new_n1098), .B2(new_n1092), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1093), .A2(new_n1094), .A3(KEYINPUT117), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(new_n748), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1096), .A2(new_n1101), .ZN(G390));
  OAI221_X1 g0902(.A(new_n1071), .B1(new_n785), .B2(new_n774), .C1(new_n352), .C2(new_n757), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n765), .A2(G116), .B1(new_n769), .B2(G294), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1104), .B(new_n396), .C1(new_n302), .C2(new_n772), .ZN(new_n1105));
  NOR4_X1   g0905(.A1(new_n1103), .A2(new_n1105), .A3(new_n783), .A4(new_n848), .ZN(new_n1106));
  XOR2_X1   g0906(.A(KEYINPUT54), .B(G143), .Z(new_n1107));
  AOI22_X1  g0907(.A1(new_n849), .A2(G159), .B1(new_n836), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n844), .B2(new_n757), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT119), .Z(new_n1110));
  NOR2_X1   g0910(.A1(new_n776), .A2(new_n286), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT53), .ZN(new_n1112));
  INV_X1    g0912(.A(G132), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n245), .B1(new_n764), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G125), .B2(new_n769), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n762), .A2(G128), .B1(new_n833), .B2(G50), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1112), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1106), .B1(new_n1110), .B2(new_n1117), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n749), .B1(new_n401), .B2(new_n828), .C1(new_n1118), .C2(new_n793), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n930), .B2(new_n809), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT120), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n820), .A2(new_n656), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n712), .A2(new_n668), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n819), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n870), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n931), .B1(new_n906), .B2(new_n921), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n935), .A2(new_n931), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n930), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n741), .A2(G330), .A3(new_n822), .A4(new_n870), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n735), .A2(new_n737), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n625), .A2(new_n493), .A3(new_n667), .ZN(new_n1134));
  OAI21_X1  g0934(.A(G330), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n868), .B(new_n867), .C1(new_n331), .C2(new_n329), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n343), .B2(new_n344), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n864), .B1(new_n862), .B2(new_n335), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n822), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1126), .B1(new_n1124), .B2(new_n870), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n922), .A2(new_n929), .B1(new_n931), .B2(new_n935), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1132), .A2(new_n1143), .A3(new_n748), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1121), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT118), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1132), .A2(new_n1143), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n870), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n1135), .B2(new_n821), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1131), .A2(new_n1149), .A3(new_n819), .A4(new_n1123), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n933), .A2(new_n934), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n738), .A2(new_n740), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n736), .B1(new_n735), .B2(new_n737), .ZN(new_n1153));
  OAI211_X1 g0953(.A(G330), .B(new_n822), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1140), .B1(new_n1154), .B2(new_n1148), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1150), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n627), .A2(G330), .A3(new_n861), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n939), .A2(new_n1157), .A3(new_n660), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1146), .B1(new_n1147), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1154), .A2(new_n1148), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1140), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1151), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1158), .B1(new_n1166), .B2(new_n1150), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1167), .A2(KEYINPUT118), .A3(new_n1132), .A4(new_n1143), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1161), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1089), .B1(new_n1147), .B2(new_n1160), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1145), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(G378));
  AOI22_X1  g0972(.A1(new_n765), .A2(G107), .B1(new_n769), .B2(G283), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n360), .B2(new_n772), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1042), .B(new_n1174), .C1(G68), .C2(new_n849), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n775), .A2(new_n376), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n757), .A2(new_n302), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(G116), .C2(new_n762), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1175), .A2(new_n254), .A3(new_n799), .A4(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT58), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  AOI21_X1  g0982(.A(G50), .B1(new_n301), .B2(new_n254), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n800), .B2(G41), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n963), .A2(new_n1107), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT122), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G128), .B2(new_n765), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n756), .A2(G132), .B1(new_n836), .B2(G137), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT121), .Z(new_n1190));
  AOI22_X1  g0990(.A1(G150), .A2(new_n849), .B1(new_n762), .B2(G125), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT123), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1188), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G33), .B(G41), .C1(new_n769), .C2(G124), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n775), .B2(new_n787), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n1193), .B2(KEYINPUT59), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1181), .B(new_n1185), .C1(new_n1194), .C2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(new_n793), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT124), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n816), .B(new_n1200), .C1(new_n290), .C2(new_n827), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n297), .A2(new_n349), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n346), .A2(new_n665), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1203), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1208), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(new_n1206), .A3(new_n1202), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1211), .A3(new_n809), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1201), .A2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(G330), .B1(new_n905), .B2(new_n910), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(new_n1211), .A3(new_n1209), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1216), .B(G330), .C1(new_n905), .C2(new_n910), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n1215), .A2(new_n938), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n938), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1213), .B1(new_n1220), .B2(new_n747), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1169), .A2(new_n1159), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT57), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1158), .B1(new_n1161), .B2(new_n1168), .ZN(new_n1226));
  OAI21_X1  g1026(.A(KEYINPUT57), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1030), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1222), .B1(new_n1225), .B2(new_n1228), .ZN(G375));
  NOR2_X1   g1029(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1230));
  OR3_X1    g1030(.A1(new_n1230), .A2(new_n1167), .A3(new_n1003), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G50), .A2(new_n849), .B1(new_n756), .B2(new_n1107), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n1113), .B2(new_n785), .C1(new_n1076), .C2(new_n776), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n765), .A2(G137), .B1(new_n769), .B2(G128), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n286), .B2(new_n772), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1233), .A2(new_n799), .A3(new_n1176), .A4(new_n1235), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G116), .A2(new_n756), .B1(new_n762), .B2(G294), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n302), .B2(new_n776), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n245), .B1(new_n769), .B2(G303), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n352), .B2(new_n772), .C1(new_n774), .C2(new_n764), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1238), .A2(new_n1240), .A3(new_n973), .A4(new_n1046), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n792), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(new_n749), .C1(G68), .C2(new_n828), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1148), .B2(new_n809), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1156), .B2(new_n748), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1231), .A2(new_n1245), .ZN(G381));
  INV_X1    g1046(.A(KEYINPUT125), .ZN(new_n1247));
  AOI21_X1  g1047(.A(G378), .B1(G375), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1247), .B2(G375), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(G390), .A2(G387), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1250), .A2(new_n1245), .A3(new_n1231), .A4(new_n1251), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1249), .A2(new_n1252), .ZN(G407));
  OAI211_X1 g1053(.A(G407), .B(G213), .C1(G343), .C2(new_n1249), .ZN(G409));
  OAI211_X1 g1054(.A(G378), .B(new_n1222), .C1(new_n1225), .C2(new_n1228), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1226), .A2(new_n1220), .A3(new_n1003), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1171), .B1(new_n1256), .B2(new_n1221), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n666), .A2(G213), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1259), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT60), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1160), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT126), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(KEYINPUT126), .A3(new_n1160), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1089), .B1(new_n1230), .B2(KEYINPUT60), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1269), .A2(G384), .A3(new_n1245), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G384), .B1(new_n1269), .B2(new_n1245), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G2897), .B(new_n1261), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1271), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1269), .A2(G384), .A3(new_n1245), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1261), .A2(G2897), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1272), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT61), .B1(new_n1260), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1279), .B1(new_n1260), .B2(new_n1281), .ZN(new_n1282));
  XOR2_X1   g1082(.A(G393), .B(G396), .Z(new_n1283));
  AND2_X1   g1083(.A1(G390), .A2(G387), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1283), .B1(new_n1284), .B2(new_n1250), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1005), .A2(new_n1023), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1286), .A2(new_n979), .A3(new_n1101), .A4(new_n1096), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(G393), .B(G396), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G390), .A2(G387), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1285), .A2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1261), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(KEYINPUT63), .A3(new_n1280), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1278), .A2(new_n1282), .A3(new_n1291), .A4(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT62), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1292), .A2(new_n1295), .A3(new_n1280), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1272), .A2(new_n1276), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1297), .B1(new_n1292), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1295), .B1(new_n1292), .B2(new_n1280), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1296), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1294), .B1(new_n1301), .B2(new_n1291), .ZN(G405));
  NAND2_X1  g1102(.A1(new_n1255), .A2(KEYINPUT127), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1285), .A2(new_n1290), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1280), .A2(G375), .A3(new_n1171), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G375), .A2(new_n1171), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1281), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(new_n1305), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1304), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1303), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1307), .A2(new_n1305), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1291), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1313), .A2(KEYINPUT127), .A3(new_n1255), .A4(new_n1308), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1311), .A2(new_n1314), .ZN(G402));
endmodule


