//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT31), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n194), .B(KEYINPUT1), .C1(new_n191), .C2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n194), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n193), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(G134), .B(G137), .ZN(new_n203));
  INV_X1    g017(.A(G131), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT66), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G137), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT11), .A3(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(G137), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n208), .A2(new_n210), .A3(new_n204), .A4(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n207), .A2(G137), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n209), .A2(G134), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n213), .B(G131), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n205), .A2(new_n212), .A3(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT0), .A4(G128), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n199), .A2(new_n220), .A3(KEYINPUT0), .A4(G128), .ZN(new_n221));
  XOR2_X1   g035(.A(KEYINPUT0), .B(G128), .Z(new_n222));
  AOI22_X1  g036(.A1(new_n219), .A2(new_n221), .B1(new_n193), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n204), .A2(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n225), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n227), .A2(new_n208), .A3(new_n210), .A4(new_n211), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n202), .A2(new_n217), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G116), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT68), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G116), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n234), .A3(G119), .ZN(new_n235));
  INV_X1    g049(.A(G119), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G116), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT2), .B(G113), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n235), .A2(KEYINPUT69), .A3(new_n237), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT69), .B1(new_n235), .B2(new_n237), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n240), .B1(new_n243), .B2(new_n239), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n230), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n217), .A2(new_n202), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n219), .A2(new_n221), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n222), .A2(new_n193), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n229), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT30), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT30), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n230), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n238), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n235), .A2(KEYINPUT69), .A3(new_n237), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n239), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n240), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n246), .B1(new_n255), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(G237), .A2(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G210), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G101), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n188), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n247), .A2(new_n253), .A3(new_n250), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n253), .B1(new_n247), .B2(new_n250), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n261), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n271), .A2(new_n188), .A3(new_n245), .A4(new_n267), .ZN(new_n272));
  INV_X1    g086(.A(new_n267), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n244), .A2(KEYINPUT28), .A3(new_n250), .A4(new_n247), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n251), .A2(new_n261), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT28), .B1(new_n230), .B2(new_n244), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n273), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n187), .B1(new_n268), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n271), .A2(new_n245), .A3(new_n267), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT31), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(new_n272), .A3(new_n278), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT70), .A3(new_n187), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n282), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n276), .A2(new_n277), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n290), .B1(new_n292), .B2(new_n273), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n262), .A2(new_n267), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n289), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n275), .A2(new_n245), .A3(KEYINPUT71), .ZN(new_n296));
  OR3_X1    g110(.A1(new_n230), .A2(new_n244), .A3(KEYINPUT71), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT28), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n277), .B(KEYINPUT72), .ZN(new_n300));
  NOR4_X1   g114(.A1(new_n299), .A2(new_n300), .A3(new_n290), .A4(new_n273), .ZN(new_n301));
  OAI21_X1  g115(.A(G472), .B1(new_n295), .B2(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(KEYINPUT32), .B(new_n187), .C1(new_n268), .C2(new_n279), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n288), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G475), .ZN(new_n305));
  INV_X1    g119(.A(G140), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G125), .ZN(new_n307));
  INV_X1    g121(.A(G125), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G140), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n309), .A3(KEYINPUT16), .ZN(new_n310));
  OR3_X1    g124(.A1(new_n308), .A2(KEYINPUT16), .A3(G140), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n310), .A2(G146), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(G146), .B1(new_n310), .B2(new_n311), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT91), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n263), .A2(G143), .A3(G214), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(G143), .B1(new_n263), .B2(G214), .ZN(new_n319));
  OAI21_X1  g133(.A(G131), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n319), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n204), .A3(new_n317), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT17), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n317), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(KEYINPUT17), .A3(G131), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT91), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(new_n312), .B2(new_n314), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n316), .A2(new_n324), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n307), .A2(new_n309), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G125), .B(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT75), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n334), .A3(new_n189), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n189), .B2(new_n333), .ZN(new_n336));
  NAND2_X1  g150(.A1(KEYINPUT18), .A2(G131), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n321), .A2(new_n317), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n325), .A2(KEYINPUT18), .A3(G131), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n329), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(G113), .B(G122), .ZN(new_n342));
  INV_X1    g156(.A(G104), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n329), .A2(new_n344), .A3(new_n340), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n305), .B1(new_n348), .B2(new_n289), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n312), .B1(new_n320), .B2(new_n322), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT19), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n332), .A2(new_n334), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n352), .B1(new_n351), .B2(new_n333), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n350), .B1(new_n353), .B2(G146), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n340), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n345), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n347), .ZN(new_n357));
  NOR2_X1   g171(.A1(G475), .A2(G902), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT20), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT20), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n361), .A3(new_n358), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n349), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G128), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G143), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT13), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n207), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G128), .B(G143), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n367), .B(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT68), .B(G116), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G122), .ZN(new_n371));
  INV_X1    g185(.A(G107), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n231), .A2(G122), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n372), .B1(new_n371), .B2(new_n373), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n369), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n370), .A2(KEYINPUT14), .A3(G122), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n371), .A2(new_n373), .ZN(new_n379));
  OAI211_X1 g193(.A(G107), .B(new_n378), .C1(new_n379), .C2(KEYINPUT14), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n191), .A2(G128), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n365), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT92), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n368), .A2(KEYINPUT92), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G134), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n386), .A3(new_n207), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n374), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n377), .B1(new_n381), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT9), .B(G234), .ZN(new_n392));
  INV_X1    g206(.A(G217), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n392), .A2(new_n393), .A3(G953), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n380), .A2(new_n374), .A3(new_n389), .A4(new_n388), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n377), .A3(new_n394), .ZN(new_n398));
  AOI21_X1  g212(.A(G902), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G478), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n399), .B1(KEYINPUT15), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n398), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n394), .B1(new_n397), .B2(new_n377), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n289), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n400), .A2(KEYINPUT15), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n363), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G952), .ZN(new_n410));
  AOI211_X1 g224(.A(G953), .B(new_n410), .C1(G234), .C2(G237), .ZN(new_n411));
  NAND2_X1  g225(.A1(G234), .A2(G237), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(G902), .A3(G953), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT93), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT21), .B(G898), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT25), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n313), .A2(new_n315), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n364), .A2(KEYINPUT23), .A3(G119), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT73), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT74), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n423), .B1(new_n236), .B2(G128), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT23), .B1(new_n364), .B2(G119), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n364), .A2(KEYINPUT74), .A3(G119), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G110), .ZN(new_n429));
  XOR2_X1   g243(.A(G119), .B(G128), .Z(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT24), .B(G110), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n419), .B(new_n429), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n431), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n428), .B2(G110), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n335), .A3(new_n313), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT22), .B(G137), .ZN(new_n436));
  INV_X1    g250(.A(G953), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(G221), .A3(G234), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n436), .B(new_n438), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n432), .A2(new_n435), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n432), .B2(new_n435), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n440), .A2(new_n441), .A3(G902), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT76), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n418), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n441), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n432), .A2(new_n435), .A3(new_n439), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n289), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(KEYINPUT76), .A3(KEYINPUT25), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n393), .B1(G234), .B2(new_n289), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n440), .A2(new_n441), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n449), .A2(G902), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT77), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT78), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n454), .A2(KEYINPUT78), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n450), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n304), .A2(new_n417), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G214), .B1(G237), .B2(G902), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT67), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(G128), .A3(new_n195), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n193), .A2(new_n364), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n462), .A2(new_n193), .B1(new_n463), .B2(new_n200), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n308), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n308), .B2(new_n223), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT7), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT88), .B(G224), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(G953), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n466), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  OAI221_X1 g284(.A(new_n465), .B1(new_n308), .B2(new_n223), .C1(G953), .C2(new_n468), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(new_n467), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT81), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n372), .A3(G104), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT3), .ZN(new_n475));
  INV_X1    g289(.A(G101), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT3), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n473), .A2(new_n477), .A3(new_n372), .A4(G104), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n343), .A2(G107), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n475), .A2(new_n476), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT82), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n372), .A3(G104), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(KEYINPUT82), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n343), .A2(G107), .ZN(new_n484));
  OAI211_X1 g298(.A(G101), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT84), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT84), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n480), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT5), .B1(new_n241), .B2(new_n242), .ZN(new_n491));
  OAI21_X1  g305(.A(G113), .B1(new_n237), .B2(KEYINPUT5), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n490), .A2(new_n494), .A3(new_n260), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n475), .A2(new_n478), .A3(new_n479), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(G101), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(G101), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(KEYINPUT4), .A3(new_n480), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n261), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(G110), .B(G122), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n472), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n493), .B1(new_n238), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n490), .A2(new_n260), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n240), .B1(new_n491), .B2(new_n493), .ZN(new_n510));
  INV_X1    g324(.A(new_n486), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n503), .B(KEYINPUT8), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n289), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT87), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n502), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT6), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n495), .A2(KEYINPUT87), .A3(new_n501), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .A4(new_n504), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n466), .A2(new_n469), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n471), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n495), .A2(KEYINPUT87), .A3(new_n501), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT87), .B1(new_n495), .B2(new_n501), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n524), .A2(new_n525), .A3(new_n503), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n500), .A2(new_n498), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n527), .A2(new_n261), .B1(new_n510), .B2(new_n490), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n503), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT6), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n521), .B(new_n523), .C1(new_n526), .C2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT89), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n504), .B1(new_n528), .B2(KEYINPUT87), .ZN(new_n534));
  OAI211_X1 g348(.A(KEYINPUT6), .B(new_n529), .C1(new_n534), .C2(new_n524), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n535), .A2(KEYINPUT89), .A3(new_n521), .A4(new_n523), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n516), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(G210), .B1(G237), .B2(G902), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n538), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT90), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n540), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  AOI211_X1 g356(.A(KEYINPUT90), .B(new_n516), .C1(new_n533), .C2(new_n536), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G469), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT10), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n198), .B2(new_n201), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n480), .A2(new_n485), .A3(new_n488), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n488), .B1(new_n480), .B2(new_n485), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n500), .A2(new_n498), .A3(new_n223), .ZN(new_n551));
  INV_X1    g365(.A(new_n229), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n460), .A2(KEYINPUT83), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT83), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n190), .A2(new_n554), .A3(KEYINPUT1), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(G128), .A3(new_n555), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n556), .A2(new_n193), .B1(new_n463), .B2(new_n200), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n546), .B1(new_n557), .B2(new_n486), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n550), .A2(new_n551), .A3(new_n552), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n437), .A2(G227), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT80), .ZN(new_n561));
  XNOR2_X1  g375(.A(G110), .B(G140), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n561), .B(new_n562), .Z(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n487), .A2(new_n489), .A3(new_n464), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n557), .A2(new_n486), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT12), .B1(new_n229), .B2(KEYINPUT85), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n229), .A3(new_n569), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n548), .A2(new_n549), .A3(new_n202), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n557), .A2(new_n486), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n229), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n568), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n564), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n550), .A2(new_n551), .A3(new_n558), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n229), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n563), .B1(new_n577), .B2(new_n559), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n545), .B(new_n289), .C1(new_n575), .C2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT86), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n569), .B1(new_n567), .B2(new_n229), .ZN(new_n582));
  AOI211_X1 g396(.A(new_n552), .B(new_n568), .C1(new_n565), .C2(new_n566), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n559), .B(new_n563), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n577), .A2(new_n559), .ZN(new_n585));
  INV_X1    g399(.A(new_n563), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n588), .A2(KEYINPUT86), .A3(new_n545), .A4(new_n289), .ZN(new_n589));
  INV_X1    g403(.A(new_n564), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n577), .ZN(new_n591));
  INV_X1    g405(.A(new_n559), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(new_n574), .B2(new_n570), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n591), .B1(new_n593), .B2(new_n563), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n289), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n581), .A2(new_n589), .B1(new_n595), .B2(G469), .ZN(new_n596));
  INV_X1    g410(.A(G221), .ZN(new_n597));
  INV_X1    g411(.A(new_n392), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n597), .B1(new_n598), .B2(new_n289), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n599), .B(KEYINPUT79), .Z(new_n600));
  NOR2_X1   g414(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n458), .A2(new_n459), .A3(new_n544), .A4(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  NAND2_X1  g417(.A1(new_n396), .A2(new_n398), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n400), .A2(G902), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n399), .A2(new_n609), .A3(G478), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT94), .B1(new_n404), .B2(new_n400), .ZN(new_n611));
  OAI22_X1  g425(.A1(new_n606), .A2(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n349), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n361), .B1(new_n357), .B2(new_n358), .ZN(new_n614));
  INV_X1    g428(.A(new_n358), .ZN(new_n615));
  AOI211_X1 g429(.A(KEYINPUT20), .B(new_n615), .C1(new_n356), .C2(new_n347), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n613), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n416), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n533), .A2(new_n536), .ZN(new_n620));
  INV_X1    g434(.A(new_n516), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n538), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI211_X1 g436(.A(new_n540), .B(new_n516), .C1(new_n533), .C2(new_n536), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n459), .B(new_n619), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n286), .ZN(new_n626));
  OAI21_X1  g440(.A(G472), .B1(new_n626), .B2(G902), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n457), .A2(new_n282), .A3(new_n287), .A4(new_n627), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n628), .A2(new_n596), .A3(new_n600), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  OAI21_X1  g446(.A(new_n459), .B1(new_n622), .B2(new_n623), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n360), .A2(KEYINPUT95), .A3(new_n362), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT95), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n614), .B2(new_n616), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n349), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n416), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(new_n638), .A3(new_n407), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT96), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT96), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n637), .A2(new_n641), .A3(new_n638), .A4(new_n407), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n633), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n629), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  NAND3_X1  g461(.A1(new_n627), .A2(new_n282), .A3(new_n287), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n432), .A2(new_n435), .ZN(new_n649));
  INV_X1    g463(.A(new_n439), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n649), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n453), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n450), .A2(new_n653), .ZN(new_n654));
  NOR4_X1   g468(.A1(new_n648), .A2(new_n416), .A3(new_n409), .A4(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n544), .A2(new_n655), .A3(new_n459), .A4(new_n601), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT97), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n656), .B(new_n658), .ZN(G12));
  OAI211_X1 g473(.A(new_n601), .B(new_n459), .C1(new_n622), .C2(new_n623), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n411), .B1(new_n414), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n637), .A2(new_n407), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n654), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n304), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  XOR2_X1   g483(.A(new_n544), .B(KEYINPUT38), .Z(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n262), .A2(new_n273), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n296), .A2(new_n297), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n289), .B1(new_n674), .B2(new_n267), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n288), .A2(new_n303), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT98), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n288), .A2(KEYINPUT98), .A3(new_n303), .A4(new_n676), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n663), .B(KEYINPUT39), .Z(new_n683));
  NAND2_X1  g497(.A1(new_n601), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n684), .A2(KEYINPUT40), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(KEYINPUT40), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n363), .A2(new_n408), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n654), .A2(new_n459), .A3(new_n687), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n682), .A2(new_n685), .A3(new_n686), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n671), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G143), .ZN(G45));
  INV_X1    g505(.A(new_n459), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n620), .A2(new_n621), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n540), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n692), .B1(new_n694), .B2(new_n539), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n612), .A2(new_n617), .A3(new_n664), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n654), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n695), .A2(new_n601), .A3(new_n304), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT99), .B(G146), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G48));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n588), .A2(new_n289), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n581), .A2(new_n589), .B1(G469), .B2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n599), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n703), .A2(KEYINPUT100), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(KEYINPUT100), .B1(new_n703), .B2(new_n704), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n701), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT100), .ZN(new_n708));
  AOI21_X1  g522(.A(G902), .B1(new_n584), .B2(new_n587), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT86), .B1(new_n709), .B2(new_n545), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n579), .A2(new_n580), .ZN(new_n711));
  OAI22_X1  g525(.A1(new_n710), .A2(new_n711), .B1(new_n545), .B2(new_n709), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n708), .B1(new_n712), .B2(new_n599), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n703), .A2(KEYINPUT100), .A3(new_n704), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(KEYINPUT101), .A3(new_n714), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n304), .A2(new_n457), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n625), .A2(new_n707), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND4_X1  g533(.A1(new_n644), .A2(new_n716), .A3(new_n707), .A4(new_n715), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  INV_X1    g535(.A(new_n654), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n304), .A2(new_n417), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n705), .A2(new_n706), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n724), .A3(new_n695), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  OAI211_X1 g540(.A(new_n459), .B(new_n687), .C1(new_n622), .C2(new_n623), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT102), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT72), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n277), .B(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n267), .B1(new_n731), .B2(new_n298), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n729), .B1(new_n732), .B2(new_n268), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n272), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n732), .A2(new_n268), .A3(new_n729), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n187), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n638), .A2(new_n736), .A3(new_n457), .A4(new_n627), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n728), .A2(new_n707), .A3(new_n715), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  INV_X1    g553(.A(new_n696), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n736), .A2(new_n740), .A3(new_n627), .A4(new_n722), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n724), .A3(new_n695), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n692), .B1(new_n537), .B2(new_n538), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n746), .B1(new_n542), .B2(new_n543), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT105), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT105), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n749), .B(new_n746), .C1(new_n542), .C2(new_n543), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT104), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n581), .A2(new_n589), .ZN(new_n752));
  NAND2_X1  g566(.A1(G469), .A2(G902), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT103), .ZN(new_n754));
  INV_X1    g568(.A(new_n594), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n754), .B1(new_n755), .B2(G469), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n751), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n752), .A2(new_n756), .A3(new_n751), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n599), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n748), .A2(new_n716), .A3(new_n750), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n745), .B1(new_n761), .B2(new_n696), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  INV_X1    g577(.A(new_n303), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT32), .B1(new_n286), .B2(new_n187), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n280), .A2(new_n283), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(KEYINPUT106), .A3(new_n303), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n302), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n696), .A2(new_n745), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n769), .A2(new_n457), .A3(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n748), .A2(new_n750), .A3(new_n760), .A4(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n762), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G131), .ZN(G33));
  NOR2_X1   g591(.A1(new_n761), .A2(new_n665), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n207), .ZN(G36));
  NAND2_X1  g593(.A1(new_n612), .A2(new_n363), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT109), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT43), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n648), .A3(new_n722), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(KEYINPUT111), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(KEYINPUT111), .ZN(new_n787));
  OR3_X1    g601(.A1(new_n783), .A2(KEYINPUT110), .A3(new_n784), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT110), .B1(new_n783), .B2(new_n784), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n786), .A2(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n748), .A2(new_n750), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n545), .B1(new_n594), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT108), .ZN(new_n795));
  OAI22_X1  g609(.A1(new_n794), .A2(new_n795), .B1(new_n793), .B2(new_n594), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n754), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(KEYINPUT46), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n752), .B1(new_n798), .B2(KEYINPUT46), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n704), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n683), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n790), .A2(new_n792), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  XNOR2_X1  g619(.A(new_n801), .B(KEYINPUT47), .ZN(new_n806));
  INV_X1    g620(.A(new_n457), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n740), .ZN(new_n808));
  OR4_X1    g622(.A1(new_n304), .A2(new_n806), .A3(new_n791), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  NAND2_X1  g624(.A1(new_n782), .A2(new_n411), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n736), .A2(new_n627), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n457), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n692), .A3(new_n724), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n671), .A2(new_n815), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n816), .A2(KEYINPUT50), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(KEYINPUT50), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n713), .A2(new_n714), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n791), .A2(new_n819), .A3(new_n811), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n812), .A2(new_n722), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n817), .A2(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n791), .A2(new_n819), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n682), .A2(new_n411), .A3(new_n457), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n825), .A2(KEYINPUT115), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(KEYINPUT115), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n612), .A2(new_n617), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n822), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n792), .A2(new_n814), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n703), .A2(new_n600), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n831), .B1(new_n806), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n830), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n819), .A2(new_n633), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n814), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(G952), .A3(new_n437), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n769), .A2(new_n457), .ZN(new_n839));
  NOR4_X1   g653(.A1(new_n791), .A2(new_n819), .A3(new_n839), .A4(new_n811), .ZN(new_n840));
  AND2_X1   g654(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n826), .A2(new_n827), .ZN(new_n844));
  OAI221_X1 g658(.A(new_n842), .B1(new_n840), .B2(new_n843), .C1(new_n844), .C2(new_n618), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n835), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n833), .B1(new_n830), .B2(KEYINPUT116), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n822), .A2(new_n848), .A3(new_n829), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n850), .A2(KEYINPUT117), .A3(new_n834), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT117), .B1(new_n850), .B2(new_n834), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n846), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  MUX2_X1   g667(.A(new_n612), .B(new_n407), .S(new_n363), .Z(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(new_n638), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n629), .A2(new_n544), .A3(new_n855), .A4(new_n459), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n602), .A2(new_n856), .A3(new_n656), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n602), .A2(new_n856), .A3(new_n656), .A4(KEYINPUT112), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI211_X1 g675(.A(new_n407), .B(new_n663), .C1(new_n450), .C2(new_n653), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n304), .A2(new_n601), .A3(new_n637), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n759), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n704), .B1(new_n864), .B2(new_n757), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n865), .B2(new_n741), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(new_n750), .A3(new_n748), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n761), .B2(new_n665), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n720), .A2(new_n717), .A3(new_n738), .A4(new_n725), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n776), .A2(new_n861), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n668), .A2(new_n743), .A3(new_n698), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n722), .A2(new_n663), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n681), .A2(new_n728), .A3(new_n760), .A4(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT52), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n836), .A2(new_n742), .B1(new_n661), .B2(new_n667), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n728), .A2(new_n681), .A3(new_n760), .A4(new_n873), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n876), .A2(new_n877), .A3(new_n698), .A4(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n875), .B(new_n879), .C1(new_n877), .C2(new_n876), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n871), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(KEYINPUT53), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n875), .A2(new_n879), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(new_n776), .A3(new_n861), .A4(new_n870), .ZN(new_n884));
  XNOR2_X1  g698(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n882), .B1(KEYINPUT114), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(KEYINPUT114), .B2(new_n886), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT54), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n776), .A2(new_n861), .A3(new_n870), .ZN(new_n890));
  INV_X1    g704(.A(new_n880), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(KEYINPUT53), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n875), .A2(new_n879), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n885), .B1(new_n871), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n889), .B1(KEYINPUT54), .B2(new_n895), .ZN(new_n896));
  OAI22_X1  g710(.A1(new_n853), .A2(new_n896), .B1(G952), .B2(G953), .ZN(new_n897));
  NOR4_X1   g711(.A1(new_n807), .A2(new_n780), .A3(new_n692), .A4(new_n600), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(KEYINPUT49), .B2(new_n712), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(KEYINPUT49), .B2(new_n712), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n670), .A2(new_n682), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n897), .A2(new_n901), .ZN(G75));
  NOR2_X1   g716(.A1(new_n437), .A2(G952), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AOI22_X1  g718(.A1(new_n881), .A2(KEYINPUT53), .B1(new_n884), .B2(new_n885), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n289), .ZN(new_n906));
  AOI211_X1 g720(.A(KEYINPUT119), .B(KEYINPUT56), .C1(new_n906), .C2(G210), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n535), .A2(new_n521), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n523), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT55), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n904), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n910), .B2(new_n907), .ZN(G51));
  XOR2_X1   g726(.A(new_n588), .B(KEYINPUT120), .Z(new_n913));
  XNOR2_X1  g727(.A(new_n905), .B(KEYINPUT54), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n754), .B(KEYINPUT57), .Z(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n906), .A2(new_n797), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n903), .B1(new_n916), .B2(new_n917), .ZN(G54));
  NAND3_X1  g732(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .ZN(new_n919));
  INV_X1    g733(.A(new_n357), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n921), .A2(new_n922), .A3(new_n903), .ZN(G60));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT59), .Z(new_n925));
  NOR3_X1   g739(.A1(new_n914), .A2(new_n606), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n925), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n896), .A2(new_n927), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n903), .B(new_n926), .C1(new_n928), .C2(new_n606), .ZN(G63));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n930));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT122), .ZN(new_n932));
  XOR2_X1   g746(.A(KEYINPUT121), .B(KEYINPUT60), .Z(new_n933));
  XOR2_X1   g747(.A(new_n932), .B(new_n933), .Z(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n930), .B1(new_n905), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n895), .A2(KEYINPUT123), .A3(new_n934), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n903), .B1(new_n938), .B2(new_n652), .ZN(new_n939));
  INV_X1    g753(.A(new_n451), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n936), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT124), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n936), .A2(new_n937), .A3(new_n943), .A4(new_n940), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n939), .A2(new_n942), .A3(KEYINPUT61), .A4(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT123), .B1(new_n895), .B2(new_n934), .ZN(new_n946));
  AOI211_X1 g760(.A(new_n930), .B(new_n935), .C1(new_n892), .C2(new_n894), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n652), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n948), .A2(new_n904), .A3(new_n941), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n945), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT125), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n945), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(G66));
  AOI211_X1 g770(.A(KEYINPUT126), .B(new_n869), .C1(new_n859), .C2(new_n860), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n958));
  INV_X1    g772(.A(new_n869), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n861), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n437), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(G953), .B1(new_n468), .B2(new_n415), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n908), .B1(G898), .B2(new_n437), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(G69));
  NOR2_X1   g779(.A1(new_n727), .A2(new_n839), .ZN(new_n966));
  AOI211_X1 g780(.A(new_n778), .B(new_n872), .C1(new_n803), .C2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n809), .A2(new_n776), .A3(new_n804), .A4(new_n967), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n968), .A2(G953), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n255), .B(new_n353), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(G900), .B2(G953), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n872), .B1(new_n671), .B2(new_n689), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n974));
  INV_X1    g788(.A(new_n684), .ZN(new_n975));
  AND4_X1   g789(.A1(new_n716), .A2(new_n792), .A3(new_n975), .A4(new_n854), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n973), .B2(KEYINPUT62), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n809), .A2(new_n804), .A3(new_n974), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n437), .ZN(new_n979));
  AOI22_X1  g793(.A1(new_n969), .A2(new_n971), .B1(new_n979), .B2(new_n970), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n437), .B1(G227), .B2(G900), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n980), .B(new_n981), .Z(G72));
  NOR3_X1   g796(.A1(new_n968), .A2(new_n957), .A3(new_n960), .ZN(new_n983));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n273), .B(new_n262), .C1(new_n983), .C2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(KEYINPUT127), .B1(new_n262), .B2(new_n267), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(new_n294), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n888), .A2(new_n985), .A3(new_n989), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n978), .A2(new_n957), .A3(new_n960), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n673), .B1(new_n991), .B2(new_n986), .ZN(new_n992));
  AND4_X1   g806(.A1(new_n904), .A2(new_n987), .A3(new_n990), .A4(new_n992), .ZN(G57));
endmodule


