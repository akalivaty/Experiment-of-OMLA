

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589;

  XOR2_X1 U323 ( .A(n366), .B(n365), .Z(n517) );
  XNOR2_X1 U324 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U325 ( .A(n396), .B(n395), .Z(n291) );
  INV_X1 U326 ( .A(KEYINPUT90), .ZN(n354) );
  XNOR2_X1 U327 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n433) );
  XNOR2_X1 U328 ( .A(n355), .B(n354), .ZN(n356) );
  NOR2_X1 U329 ( .A1(n545), .A2(n520), .ZN(n526) );
  XNOR2_X1 U330 ( .A(n357), .B(n356), .ZN(n438) );
  XNOR2_X1 U331 ( .A(n397), .B(n291), .ZN(n398) );
  NOR2_X1 U332 ( .A1(n471), .A2(n470), .ZN(n484) );
  XNOR2_X1 U333 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U334 ( .A(n326), .B(n325), .ZN(n525) );
  XNOR2_X1 U335 ( .A(n454), .B(KEYINPUT120), .ZN(n455) );
  XNOR2_X1 U336 ( .A(n478), .B(G36GAT), .ZN(n479) );
  XNOR2_X1 U337 ( .A(n456), .B(n455), .ZN(G1348GAT) );
  XNOR2_X1 U338 ( .A(n480), .B(n479), .ZN(G1329GAT) );
  XOR2_X1 U339 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n293) );
  XNOR2_X1 U340 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n292) );
  XNOR2_X1 U341 ( .A(n293), .B(n292), .ZN(n301) );
  XNOR2_X1 U342 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n294), .B(KEYINPUT7), .ZN(n406) );
  XNOR2_X1 U344 ( .A(G22GAT), .B(G1GAT), .ZN(n295) );
  XNOR2_X1 U345 ( .A(n295), .B(KEYINPUT69), .ZN(n373) );
  XNOR2_X1 U346 ( .A(n406), .B(n373), .ZN(n299) );
  XOR2_X1 U347 ( .A(KEYINPUT30), .B(G8GAT), .Z(n297) );
  XNOR2_X1 U348 ( .A(G197GAT), .B(G141GAT), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n309) );
  NAND2_X1 U352 ( .A1(G229GAT), .A2(G233GAT), .ZN(n307) );
  XOR2_X1 U353 ( .A(G15GAT), .B(G113GAT), .Z(n303) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(G50GAT), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n305) );
  XOR2_X1 U356 ( .A(G36GAT), .B(G43GAT), .Z(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n575) );
  XOR2_X1 U360 ( .A(KEYINPUT86), .B(KEYINPUT83), .Z(n315) );
  XOR2_X1 U361 ( .A(KEYINPUT85), .B(KEYINPUT82), .Z(n311) );
  XNOR2_X1 U362 ( .A(G190GAT), .B(KEYINPUT20), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n313) );
  XNOR2_X1 U364 ( .A(G99GAT), .B(G71GAT), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n312), .B(G120GAT), .ZN(n394) );
  XNOR2_X1 U366 ( .A(n313), .B(n394), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U368 ( .A(G15GAT), .B(G127GAT), .Z(n374) );
  XOR2_X1 U369 ( .A(G113GAT), .B(KEYINPUT0), .Z(n338) );
  XOR2_X1 U370 ( .A(n374), .B(n338), .Z(n317) );
  NAND2_X1 U371 ( .A1(G227GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U373 ( .A(n319), .B(n318), .Z(n326) );
  XOR2_X1 U374 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n321) );
  XNOR2_X1 U375 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U377 ( .A(n322), .B(G183GAT), .Z(n324) );
  XNOR2_X1 U378 ( .A(G169GAT), .B(G176GAT), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n351) );
  XOR2_X1 U380 ( .A(G43GAT), .B(G134GAT), .Z(n416) );
  XNOR2_X1 U381 ( .A(n351), .B(n416), .ZN(n325) );
  XOR2_X1 U382 ( .A(KEYINPUT4), .B(G148GAT), .Z(n328) );
  XNOR2_X1 U383 ( .A(G120GAT), .B(G127GAT), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U385 ( .A(KEYINPUT6), .B(KEYINPUT94), .Z(n330) );
  XNOR2_X1 U386 ( .A(KEYINPUT5), .B(KEYINPUT95), .ZN(n329) );
  XNOR2_X1 U387 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U388 ( .A(n332), .B(n331), .Z(n337) );
  XOR2_X1 U389 ( .A(KEYINPUT93), .B(KEYINPUT1), .Z(n334) );
  NAND2_X1 U390 ( .A1(G225GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U392 ( .A(G1GAT), .B(n335), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n342) );
  XOR2_X1 U394 ( .A(G85GAT), .B(G57GAT), .Z(n389) );
  XOR2_X1 U395 ( .A(KEYINPUT75), .B(n389), .Z(n340) );
  XNOR2_X1 U396 ( .A(n338), .B(G162GAT), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U398 ( .A(n342), .B(n341), .Z(n344) );
  XNOR2_X1 U399 ( .A(G29GAT), .B(G134GAT), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n344), .B(n343), .ZN(n349) );
  XOR2_X1 U401 ( .A(KEYINPUT2), .B(KEYINPUT92), .Z(n346) );
  XNOR2_X1 U402 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U404 ( .A(G141GAT), .B(n347), .Z(n437) );
  INV_X1 U405 ( .A(n437), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n514) );
  XNOR2_X1 U407 ( .A(G204GAT), .B(G92GAT), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n350), .B(G64GAT), .ZN(n390) );
  XNOR2_X1 U409 ( .A(n351), .B(n390), .ZN(n366) );
  XOR2_X1 U410 ( .A(G36GAT), .B(G190GAT), .Z(n410) );
  XOR2_X1 U411 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n353) );
  XNOR2_X1 U412 ( .A(G218GAT), .B(KEYINPUT89), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n357) );
  XNOR2_X1 U414 ( .A(G197GAT), .B(G211GAT), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n410), .B(n438), .ZN(n361) );
  INV_X1 U416 ( .A(n361), .ZN(n359) );
  NAND2_X1 U417 ( .A1(G226GAT), .A2(G233GAT), .ZN(n360) );
  INV_X1 U418 ( .A(n360), .ZN(n358) );
  NAND2_X1 U419 ( .A1(n359), .A2(n358), .ZN(n363) );
  NAND2_X1 U420 ( .A1(n361), .A2(n360), .ZN(n362) );
  NAND2_X1 U421 ( .A1(n363), .A2(n362), .ZN(n364) );
  XOR2_X1 U422 ( .A(G8GAT), .B(KEYINPUT77), .Z(n369) );
  XNOR2_X1 U423 ( .A(n364), .B(n369), .ZN(n365) );
  XOR2_X1 U424 ( .A(KEYINPUT117), .B(n517), .Z(n432) );
  XOR2_X1 U425 ( .A(G57GAT), .B(G78GAT), .Z(n368) );
  XNOR2_X1 U426 ( .A(G211GAT), .B(G155GAT), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n370) );
  XOR2_X1 U428 ( .A(n370), .B(n369), .Z(n372) );
  XNOR2_X1 U429 ( .A(G183GAT), .B(G71GAT), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n378) );
  XOR2_X1 U431 ( .A(n374), .B(n373), .Z(n376) );
  NAND2_X1 U432 ( .A1(G231GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U434 ( .A(n378), .B(n377), .Z(n386) );
  XOR2_X1 U435 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n380) );
  XNOR2_X1 U436 ( .A(KEYINPUT13), .B(G64GAT), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U438 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n382) );
  XNOR2_X1 U439 ( .A(KEYINPUT15), .B(KEYINPUT78), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n551) );
  INV_X1 U443 ( .A(n551), .ZN(n584) );
  INV_X1 U444 ( .A(n575), .ZN(n546) );
  XOR2_X1 U445 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n388) );
  XNOR2_X1 U446 ( .A(G176GAT), .B(KEYINPUT70), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n388), .B(n387), .ZN(n401) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n392) );
  AND2_X1 U449 ( .A1(G230GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n399) );
  XNOR2_X1 U451 ( .A(G106GAT), .B(G78GAT), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n393), .B(G148GAT), .ZN(n439) );
  XNOR2_X1 U453 ( .A(n394), .B(n439), .ZN(n397) );
  XOR2_X1 U454 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n396) );
  XNOR2_X1 U455 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n395) );
  XOR2_X1 U456 ( .A(n401), .B(n400), .Z(n581) );
  XNOR2_X1 U457 ( .A(n581), .B(KEYINPUT41), .ZN(n558) );
  NAND2_X1 U458 ( .A1(n546), .A2(n558), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n402), .B(KEYINPUT46), .ZN(n423) );
  XOR2_X1 U460 ( .A(KEYINPUT11), .B(KEYINPUT65), .Z(n404) );
  XNOR2_X1 U461 ( .A(G85GAT), .B(G92GAT), .ZN(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U463 ( .A(KEYINPUT10), .B(n405), .Z(n408) );
  XNOR2_X1 U464 ( .A(n406), .B(KEYINPUT75), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n422) );
  XNOR2_X1 U466 ( .A(G50GAT), .B(KEYINPUT73), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n409), .B(G162GAT), .ZN(n440) );
  XOR2_X1 U468 ( .A(n410), .B(n440), .Z(n412) );
  NAND2_X1 U469 ( .A1(G232GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n412), .B(n411), .ZN(n420) );
  XOR2_X1 U471 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n414) );
  XNOR2_X1 U472 ( .A(G218GAT), .B(KEYINPUT74), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U474 ( .A(n415), .B(G106GAT), .Z(n418) );
  XNOR2_X1 U475 ( .A(G99GAT), .B(n416), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U477 ( .A(n420), .B(n419), .Z(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n570) );
  AND2_X1 U479 ( .A1(n423), .A2(n570), .ZN(n424) );
  AND2_X1 U480 ( .A1(n584), .A2(n424), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n425), .B(KEYINPUT47), .ZN(n430) );
  INV_X1 U482 ( .A(n581), .ZN(n476) );
  XNOR2_X1 U483 ( .A(KEYINPUT36), .B(n570), .ZN(n587) );
  NOR2_X1 U484 ( .A1(n587), .A2(n584), .ZN(n426) );
  XOR2_X1 U485 ( .A(KEYINPUT45), .B(n426), .Z(n427) );
  NOR2_X1 U486 ( .A1(n476), .A2(n427), .ZN(n428) );
  NAND2_X1 U487 ( .A1(n428), .A2(n575), .ZN(n429) );
  NAND2_X1 U488 ( .A1(n430), .A2(n429), .ZN(n431) );
  XNOR2_X1 U489 ( .A(KEYINPUT48), .B(n431), .ZN(n543) );
  NAND2_X1 U490 ( .A1(n432), .A2(n543), .ZN(n434) );
  NOR2_X1 U491 ( .A1(n514), .A2(n435), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n436), .B(KEYINPUT64), .ZN(n574) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n450) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n448) );
  NAND2_X1 U495 ( .A1(G228GAT), .A2(G233GAT), .ZN(n446) );
  XOR2_X1 U496 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n442) );
  XNOR2_X1 U497 ( .A(G22GAT), .B(KEYINPUT88), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U499 ( .A(KEYINPUT24), .B(G204GAT), .Z(n443) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U502 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n450), .B(n449), .ZN(n467) );
  NAND2_X1 U504 ( .A1(n574), .A2(n467), .ZN(n452) );
  XOR2_X1 U505 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n451) );
  XNOR2_X1 U506 ( .A(n452), .B(n451), .ZN(n453) );
  NAND2_X1 U507 ( .A1(n525), .A2(n453), .ZN(n569) );
  NOR2_X1 U508 ( .A1(n575), .A2(n569), .ZN(n456) );
  INV_X1 U509 ( .A(G169GAT), .ZN(n454) );
  INV_X1 U510 ( .A(KEYINPUT100), .ZN(n473) );
  NAND2_X1 U511 ( .A1(n517), .A2(n525), .ZN(n458) );
  INV_X1 U512 ( .A(KEYINPUT97), .ZN(n457) );
  XNOR2_X1 U513 ( .A(n458), .B(n457), .ZN(n459) );
  NAND2_X1 U514 ( .A1(n459), .A2(n467), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n460), .B(KEYINPUT25), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n517), .B(KEYINPUT27), .ZN(n466) );
  NOR2_X1 U517 ( .A1(n525), .A2(n467), .ZN(n461) );
  XNOR2_X1 U518 ( .A(KEYINPUT26), .B(n461), .ZN(n573) );
  AND2_X1 U519 ( .A1(n466), .A2(n573), .ZN(n462) );
  NOR2_X1 U520 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n464), .B(KEYINPUT98), .ZN(n465) );
  NOR2_X1 U522 ( .A1(n514), .A2(n465), .ZN(n471) );
  NAND2_X1 U523 ( .A1(n514), .A2(n466), .ZN(n545) );
  XOR2_X1 U524 ( .A(KEYINPUT28), .B(n467), .Z(n520) );
  XOR2_X1 U525 ( .A(n526), .B(KEYINPUT96), .Z(n469) );
  XOR2_X1 U526 ( .A(n525), .B(KEYINPUT87), .Z(n468) );
  NOR2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n551), .A2(n484), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n473), .B(n472), .ZN(n474) );
  NOR2_X1 U530 ( .A1(n587), .A2(n474), .ZN(n475) );
  XOR2_X1 U531 ( .A(KEYINPUT37), .B(n475), .Z(n513) );
  NOR2_X1 U532 ( .A1(n575), .A2(n476), .ZN(n485) );
  NAND2_X1 U533 ( .A1(n513), .A2(n485), .ZN(n477) );
  XOR2_X1 U534 ( .A(KEYINPUT38), .B(n477), .Z(n499) );
  NAND2_X1 U535 ( .A1(n499), .A2(n517), .ZN(n480) );
  XOR2_X1 U536 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n478) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n482) );
  NAND2_X1 U538 ( .A1(n551), .A2(n570), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(n483) );
  NOR2_X1 U540 ( .A1(n484), .A2(n483), .ZN(n503) );
  AND2_X1 U541 ( .A1(n485), .A2(n503), .ZN(n492) );
  NAND2_X1 U542 ( .A1(n492), .A2(n514), .ZN(n486) );
  XNOR2_X1 U543 ( .A(n486), .B(KEYINPUT34), .ZN(n487) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  XOR2_X1 U545 ( .A(G8GAT), .B(KEYINPUT99), .Z(n489) );
  NAND2_X1 U546 ( .A1(n492), .A2(n517), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT35), .Z(n491) );
  NAND2_X1 U549 ( .A1(n492), .A2(n525), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  NAND2_X1 U551 ( .A1(n520), .A2(n492), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n493), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .Z(n495) );
  NAND2_X1 U554 ( .A1(n514), .A2(n499), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NAND2_X1 U556 ( .A1(n525), .A2(n499), .ZN(n497) );
  XOR2_X1 U557 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n499), .A2(n520), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n500), .B(KEYINPUT104), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(n501), .ZN(G1331GAT) );
  NAND2_X1 U563 ( .A1(n558), .A2(n575), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n502), .B(KEYINPUT105), .ZN(n512) );
  AND2_X1 U565 ( .A1(n512), .A2(n503), .ZN(n508) );
  NAND2_X1 U566 ( .A1(n514), .A2(n508), .ZN(n504) );
  XNOR2_X1 U567 ( .A(KEYINPUT42), .B(n504), .ZN(n505) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n517), .A2(n508), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n508), .A2(n525), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U574 ( .A1(n508), .A2(n520), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(n511), .ZN(G1335GAT) );
  XOR2_X1 U577 ( .A(G85GAT), .B(KEYINPUT107), .Z(n516) );
  AND2_X1 U578 ( .A1(n513), .A2(n512), .ZN(n521) );
  NAND2_X1 U579 ( .A1(n521), .A2(n514), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n517), .A2(n521), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n521), .A2(n525), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n523) );
  NAND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U588 ( .A(G106GAT), .B(n524), .Z(G1339GAT) );
  INV_X1 U589 ( .A(n525), .ZN(n528) );
  NAND2_X1 U590 ( .A1(n543), .A2(n526), .ZN(n527) );
  NOR2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U592 ( .A(KEYINPUT109), .B(n529), .Z(n540) );
  NAND2_X1 U593 ( .A1(n540), .A2(n546), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(KEYINPUT110), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U597 ( .A1(n540), .A2(n558), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(KEYINPUT111), .ZN(n537) );
  XOR2_X1 U600 ( .A(KEYINPUT112), .B(KEYINPUT50), .Z(n535) );
  NAND2_X1 U601 ( .A1(n540), .A2(n551), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n539) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT114), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n542) );
  INV_X1 U607 ( .A(n570), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n540), .A2(n555), .ZN(n541) );
  XOR2_X1 U609 ( .A(n542), .B(n541), .Z(G1343GAT) );
  NAND2_X1 U610 ( .A1(n543), .A2(n573), .ZN(n544) );
  NOR2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n556), .A2(n546), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  NAND2_X1 U615 ( .A1(n556), .A2(n558), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n550), .ZN(G1345GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n553) );
  NAND2_X1 U619 ( .A1(n556), .A2(n551), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n554), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 U624 ( .A(n558), .ZN(n559) );
  NOR2_X1 U625 ( .A1(n559), .A2(n569), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n561) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT121), .B(n562), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  NOR2_X1 U631 ( .A1(n584), .A2(n569), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(G1350GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n568) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n568), .B(n567), .ZN(n572) );
  NOR2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U638 ( .A(n572), .B(n571), .Z(G1351GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n586) );
  NOR2_X1 U640 ( .A1(n575), .A2(n586), .ZN(n580) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT59), .B(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n586), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n586), .ZN(n585) );
  XOR2_X1 U650 ( .A(G211GAT), .B(n585), .Z(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

