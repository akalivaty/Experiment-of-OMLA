//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1165, new_n1166, new_n1167;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G219), .A3(G221), .A4(G220), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT68), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n459), .A2(G137), .A3(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT69), .A4(G125), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n465), .B1(new_n474), .B2(G2105), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(new_n460), .B2(G112), .ZN(new_n476));
  INV_X1    g051(.A(G100), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(new_n460), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT70), .Z(new_n479));
  INV_X1    g054(.A(new_n459), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(new_n460), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n479), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND4_X1  g061(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n460), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n459), .A2(KEYINPUT4), .A3(G138), .A4(new_n460), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n466), .A2(new_n468), .A3(G126), .A4(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n491), .A2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G651), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n502), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT72), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  OAI221_X1 g089(.A(new_n514), .B1(new_n510), .B2(new_n511), .C1(new_n509), .C2(new_n508), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(new_n507), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n513), .A2(new_n515), .B1(G651), .B2(new_n519), .ZN(G166));
  AND3_X1   g095(.A1(new_n499), .A2(new_n501), .A3(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT73), .B(G89), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n502), .A2(new_n525), .B1(G63), .B2(G651), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n522), .B(new_n524), .C1(new_n526), .C2(new_n517), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  NAND2_X1  g103(.A1(new_n521), .A2(G52), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n508), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n498), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n531), .A2(new_n533), .ZN(G171));
  NAND3_X1  g109(.A1(new_n502), .A2(G81), .A3(new_n507), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n521), .A2(G43), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n507), .A2(G56), .ZN(new_n537));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n498), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n539), .A2(KEYINPUT74), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(KEYINPUT74), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n535), .B(new_n536), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n548), .ZN(G188));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n508), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g126(.A(KEYINPUT76), .B1(new_n502), .B2(new_n507), .ZN(new_n552));
  OAI21_X1  g127(.A(G91), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n498), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT9), .B1(new_n510), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n521), .A2(new_n559), .A3(G53), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n558), .B1(new_n557), .B2(new_n560), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n553), .B(new_n555), .C1(new_n561), .C2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  NAND2_X1  g139(.A1(new_n513), .A2(new_n515), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n519), .A2(G651), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(G303));
  INV_X1    g142(.A(G49), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n507), .A2(G74), .ZN(new_n569));
  OAI22_X1  g144(.A1(new_n568), .A2(new_n510), .B1(new_n569), .B2(new_n498), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n508), .B(new_n550), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n570), .B1(new_n571), .B2(G87), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(new_n521), .A2(G48), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n498), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n571), .B2(G86), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G305));
  NAND2_X1  g153(.A1(new_n521), .A2(G47), .ZN(new_n579));
  INV_X1    g154(.A(G85), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n508), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n498), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n581), .A2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n571), .A2(G92), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n521), .A2(G54), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(new_n498), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT77), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n571), .A2(new_n592), .A3(G92), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n587), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n585), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n585), .B1(new_n595), .B2(G868), .ZN(G321));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NOR2_X1   g173(.A1(G168), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G299), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(KEYINPUT78), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(KEYINPUT78), .B2(new_n599), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(KEYINPUT78), .B2(new_n599), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n595), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n595), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n483), .A2(G123), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT80), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n481), .A2(G135), .ZN(new_n614));
  NOR2_X1   g189(.A1(G99), .A2(G2105), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(new_n460), .B2(G111), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT81), .B(G2096), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n459), .A2(new_n463), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT13), .B(G2100), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n619), .A2(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT82), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n631), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  OR3_X1    g212(.A1(new_n636), .A2(KEYINPUT83), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  OAI21_X1  g214(.A(KEYINPUT83), .B1(new_n636), .B2(new_n637), .ZN(new_n640));
  NAND4_X1  g215(.A1(new_n638), .A2(G14), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g220(.A1(new_n645), .A2(KEYINPUT17), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  AOI21_X1  g222(.A(KEYINPUT18), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n645), .B2(KEYINPUT18), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n648), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2096), .B(G2100), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(G227));
  XNOR2_X1  g228(.A(G1971), .B(G1976), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n655), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  AOI22_X1  g236(.A1(new_n659), .A2(KEYINPUT20), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n663), .A2(new_n655), .A3(new_n658), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n662), .B(new_n664), .C1(KEYINPUT20), .C2(new_n659), .ZN(new_n665));
  XOR2_X1   g240(.A(G1991), .B(G1996), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n669), .B(new_n670), .Z(G229));
  INV_X1    g246(.A(G16), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G24), .ZN(new_n673));
  INV_X1    g248(.A(G290), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n673), .B1(new_n674), .B2(new_n672), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT85), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1986), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n672), .A2(G23), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(new_n572), .B2(new_n672), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT33), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G1976), .ZN(new_n681));
  INV_X1    g256(.A(G22), .ZN(new_n682));
  OAI21_X1  g257(.A(KEYINPUT86), .B1(new_n682), .B2(G16), .ZN(new_n683));
  OR3_X1    g258(.A1(new_n682), .A2(KEYINPUT86), .A3(G16), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n683), .B(new_n684), .C1(G166), .C2(new_n672), .ZN(new_n685));
  INV_X1    g260(.A(G1971), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n672), .A2(G6), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n577), .B2(new_n672), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT32), .B(G1981), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n681), .A2(new_n687), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n677), .B1(new_n692), .B2(KEYINPUT34), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n481), .A2(G131), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n483), .A2(G119), .ZN(new_n695));
  NOR2_X1   g270(.A1(G95), .A2(G2105), .ZN(new_n696));
  OAI21_X1  g271(.A(G2104), .B1(new_n460), .B2(G107), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n694), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G25), .B(new_n698), .S(G29), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT84), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT35), .B(G1991), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n693), .B(new_n702), .C1(KEYINPUT34), .C2(new_n692), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT36), .Z(new_n704));
  NOR2_X1   g279(.A1(G5), .A2(G16), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G171), .B2(G16), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1961), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n617), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT94), .ZN(new_n710));
  NOR2_X1   g285(.A1(G164), .A2(new_n708), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G27), .B2(new_n708), .ZN(new_n712));
  INV_X1    g287(.A(G2078), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n708), .A2(G26), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n481), .A2(G140), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n483), .A2(G128), .ZN(new_n719));
  OR2_X1    g294(.A1(G104), .A2(G2105), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n720), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n717), .B1(new_n723), .B2(new_n708), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G2067), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n708), .B1(new_n726), .B2(G28), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n726), .B2(G28), .ZN(new_n728));
  NOR4_X1   g303(.A1(new_n710), .A2(new_n714), .A3(new_n725), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n708), .A2(G33), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n463), .A2(G103), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT88), .B(KEYINPUT25), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n481), .A2(G139), .ZN(new_n734));
  NAND2_X1  g309(.A1(G115), .A2(G2104), .ZN(new_n735));
  INV_X1    g310(.A(G127), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n480), .B2(new_n736), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n733), .B(new_n734), .C1(G2105), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT89), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n730), .B1(new_n740), .B2(new_n708), .ZN(new_n741));
  INV_X1    g316(.A(G2090), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n708), .A2(G35), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G162), .B2(new_n708), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT29), .Z(new_n745));
  OAI221_X1 g320(.A(new_n729), .B1(G2072), .B2(new_n741), .C1(new_n742), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n742), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n741), .A2(G2072), .ZN(new_n748));
  OR2_X1    g323(.A1(KEYINPUT24), .A2(G34), .ZN(new_n749));
  NAND2_X1  g324(.A1(KEYINPUT24), .A2(G34), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n749), .A2(new_n708), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G160), .B2(new_n708), .ZN(new_n752));
  INV_X1    g327(.A(G2084), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n747), .A2(new_n748), .A3(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT31), .B(G11), .Z(new_n756));
  NOR3_X1   g331(.A1(new_n746), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n481), .A2(G141), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n483), .A2(G129), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n463), .A2(G105), .ZN(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT26), .Z(new_n762));
  NAND4_X1  g337(.A1(new_n758), .A2(new_n759), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT90), .Z(new_n764));
  AND3_X1   g339(.A1(new_n764), .A2(KEYINPUT91), .A3(G29), .ZN(new_n765));
  AOI21_X1  g340(.A(KEYINPUT91), .B1(new_n764), .B2(G29), .ZN(new_n766));
  OAI22_X1  g341(.A1(new_n765), .A2(new_n766), .B1(G29), .B2(G32), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n672), .A2(G20), .ZN(new_n770));
  OAI211_X1 g345(.A(KEYINPUT23), .B(new_n770), .C1(new_n601), .C2(new_n672), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(KEYINPUT23), .B2(new_n770), .ZN(new_n772));
  INV_X1    g347(.A(G1956), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n672), .A2(G4), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n595), .B2(new_n672), .ZN(new_n777));
  INV_X1    g352(.A(G1348), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n543), .A2(G16), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G16), .B2(G19), .ZN(new_n781));
  INV_X1    g356(.A(G1341), .ZN(new_n782));
  OAI22_X1  g357(.A1(new_n781), .A2(new_n782), .B1(new_n713), .B2(new_n712), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT92), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G16), .B2(G21), .ZN(new_n785));
  NOR2_X1   g360(.A1(G286), .A2(new_n672), .ZN(new_n786));
  MUX2_X1   g361(.A(new_n785), .B(new_n784), .S(new_n786), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT93), .B(G1966), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n783), .B(new_n789), .C1(new_n782), .C2(new_n781), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n757), .A2(new_n775), .A3(new_n779), .A4(new_n790), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n704), .A2(new_n707), .A3(new_n791), .ZN(G311));
  INV_X1    g367(.A(G311), .ZN(G150));
  NAND2_X1  g368(.A1(new_n521), .A2(G55), .ZN(new_n794));
  INV_X1    g369(.A(G93), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n508), .B2(new_n795), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n797), .A2(new_n498), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n543), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n542), .A2(new_n799), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n803), .B(new_n804), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n595), .A2(G559), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT39), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n805), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(G860), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT96), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n800), .A2(G860), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT37), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n812), .ZN(G145));
  OR2_X1    g388(.A1(G106), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n481), .A2(G142), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(KEYINPUT98), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n481), .A2(KEYINPUT98), .A3(G142), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n483), .A2(G130), .ZN(new_n819));
  AND4_X1   g394(.A1(new_n815), .A2(new_n817), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n698), .B(new_n622), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n820), .B(new_n821), .Z(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n740), .A2(new_n764), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n739), .A2(new_n763), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n492), .A2(new_n495), .A3(KEYINPUT97), .ZN(new_n826));
  AOI21_X1  g401(.A(KEYINPUT97), .B1(new_n492), .B2(new_n495), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n489), .B(new_n490), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n722), .B(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n824), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n829), .B1(new_n824), .B2(new_n825), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n823), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n832), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n834), .A2(new_n822), .A3(new_n830), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n833), .A2(new_n835), .A3(KEYINPUT99), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G162), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n833), .A2(new_n835), .A3(KEYINPUT99), .A4(new_n485), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n617), .B(G160), .Z(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G37), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g421(.A(new_n608), .B(new_n803), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n594), .A2(new_n848), .A3(G299), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(G299), .A2(new_n848), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n553), .A2(new_n555), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n852), .B(KEYINPUT100), .C1(new_n562), .C2(new_n561), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n853), .A3(new_n594), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  OR3_X1    g430(.A1(new_n847), .A2(KEYINPUT101), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n854), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT41), .B1(new_n857), .B2(new_n849), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT41), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n850), .A2(new_n859), .A3(new_n854), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n860), .A3(KEYINPUT102), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n857), .A2(new_n849), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n863), .A3(new_n859), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n861), .A2(new_n847), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT101), .B1(new_n847), .B2(new_n855), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n856), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT42), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT42), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n856), .A2(new_n865), .A3(new_n869), .A4(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(G166), .B(new_n572), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(G305), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G290), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n868), .A2(new_n874), .A3(new_n870), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(G868), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n799), .A2(G868), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(G295));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n879), .A2(new_n883), .A3(new_n881), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n598), .B1(new_n876), .B2(new_n877), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT103), .B1(new_n885), .B2(new_n880), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(G331));
  NOR2_X1   g462(.A1(G171), .A2(KEYINPUT104), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n801), .B2(new_n802), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(G286), .B1(G171), .B2(KEYINPUT104), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n801), .A2(new_n802), .A3(new_n889), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n892), .ZN(new_n895));
  INV_X1    g470(.A(new_n893), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n896), .B2(new_n890), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n861), .A2(new_n864), .A3(new_n894), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n894), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n862), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n874), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT105), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n898), .A2(new_n874), .A3(new_n903), .A4(new_n900), .ZN(new_n904));
  AOI21_X1  g479(.A(G37), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n858), .A2(new_n860), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(new_n906), .B2(new_n858), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n900), .B1(new_n908), .B2(new_n899), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n875), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n905), .A2(KEYINPUT43), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n898), .A2(new_n900), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n875), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT43), .B1(new_n905), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT44), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n905), .A2(new_n916), .A3(new_n910), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n905), .B2(new_n913), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n915), .B1(new_n919), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g495(.A(G1966), .ZN(new_n921));
  INV_X1    g496(.A(G1384), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT45), .B1(new_n828), .B2(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(KEYINPUT45), .B(new_n922), .C1(new_n491), .C2(new_n496), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(G40), .A3(G160), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n921), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT50), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n828), .A2(new_n927), .A3(new_n922), .ZN(new_n928));
  INV_X1    g503(.A(G40), .ZN(new_n929));
  AOI211_X1 g504(.A(new_n929), .B(new_n465), .C1(new_n474), .C2(G2105), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n922), .B1(new_n491), .B2(new_n496), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT50), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n928), .A2(new_n753), .A3(new_n930), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n926), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(G8), .ZN(new_n935));
  INV_X1    g510(.A(G8), .ZN(new_n936));
  NOR3_X1   g511(.A1(G168), .A2(KEYINPUT118), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT118), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(G286), .B2(G8), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT120), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT51), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n935), .A2(new_n940), .A3(new_n941), .A4(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n936), .B1(new_n926), .B2(new_n933), .ZN(new_n946));
  INV_X1    g521(.A(new_n940), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n942), .B(new_n943), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n947), .A2(new_n934), .A3(KEYINPUT119), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT119), .B1(new_n947), .B2(new_n934), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT121), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT62), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n947), .A2(new_n934), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT119), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n947), .A2(new_n934), .A3(KEYINPUT119), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT121), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n948), .A4(new_n945), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n953), .A2(new_n954), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G86), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n508), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(G1981), .B1(new_n576), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1981), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n577), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT111), .B1(new_n577), .B2(new_n966), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n965), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT49), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AND4_X1   g548(.A1(G40), .A2(new_n828), .A3(new_n922), .A4(G160), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(new_n936), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT49), .B(new_n965), .C1(new_n969), .C2(new_n970), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT109), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n980));
  NAND4_X1  g555(.A1(G303), .A2(new_n980), .A3(KEYINPUT55), .A4(G8), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(G166), .B2(new_n936), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n979), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n931), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(KEYINPUT107), .B(G1384), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n828), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n930), .B(new_n987), .C1(new_n990), .C2(new_n986), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n686), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n927), .B(new_n922), .C1(new_n491), .C2(new_n496), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT97), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n496), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n492), .A2(new_n495), .A3(KEYINPUT97), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n491), .ZN(new_n998));
  AOI21_X1  g573(.A(G1384), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n930), .B(new_n993), .C1(new_n999), .C2(new_n927), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n992), .B1(G2090), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G8), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n985), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n572), .A2(G1976), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n975), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1976), .ZN(new_n1009));
  NAND3_X1  g584(.A1(G288), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n975), .A2(KEYINPUT110), .A3(KEYINPUT52), .A4(new_n1004), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n928), .A2(new_n930), .A3(new_n932), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n992), .B1(G2090), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n984), .A2(G8), .A3(new_n1014), .ZN(new_n1015));
  AND4_X1   g590(.A1(new_n977), .A2(new_n1003), .A3(new_n1012), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G160), .A2(G40), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n988), .B1(new_n997), .B2(new_n998), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n1018), .B2(KEYINPUT45), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(new_n713), .A3(new_n987), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OR4_X1    g597(.A1(new_n1021), .A2(new_n923), .A3(new_n925), .A4(G2078), .ZN(new_n1023));
  INV_X1    g598(.A(G1961), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1013), .A2(new_n1024), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(G301), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n962), .A2(new_n1016), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT123), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n953), .A2(new_n961), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT62), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n962), .A2(KEYINPUT123), .A3(new_n1016), .A4(new_n1027), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT124), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n977), .A2(new_n1009), .A3(new_n572), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n969), .A2(new_n970), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n975), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1014), .A2(G8), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n977), .B(new_n1012), .C1(new_n1040), .C2(new_n984), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n946), .A2(G168), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT63), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n984), .B1(new_n1001), .B2(G8), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1042), .A2(KEYINPUT63), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1015), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(new_n977), .A3(new_n1012), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1039), .A2(new_n1043), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT60), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1013), .A2(new_n778), .ZN(new_n1052));
  INV_X1    g627(.A(G2067), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n974), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n594), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n595), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1051), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT61), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1000), .A2(new_n773), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1018), .A2(KEYINPUT45), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT56), .B(G2072), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1062), .A2(new_n930), .A3(new_n987), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT57), .B1(new_n557), .B2(new_n560), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n852), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1067), .B1(new_n601), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g645(.A1(G299), .A2(KEYINPUT57), .B1(new_n852), .B2(new_n1066), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1060), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT58), .B(G1341), .ZN(new_n1074));
  OAI22_X1  g649(.A1(new_n991), .A2(G1996), .B1(new_n974), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n543), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1075), .B(new_n543), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1056), .A2(new_n1051), .A3(new_n595), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1073), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1061), .A2(KEYINPUT113), .A3(new_n1064), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT113), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1069), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1070), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n1088), .A3(KEYINPUT61), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT116), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1087), .A2(new_n1088), .A3(new_n1091), .A4(KEYINPUT61), .ZN(new_n1092));
  AOI211_X1 g667(.A(new_n1059), .B(new_n1084), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1086), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1061), .A2(KEYINPUT113), .A3(new_n1064), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1071), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1058), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1088), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1098), .B(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT117), .B1(new_n1093), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n990), .A2(new_n986), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1019), .A2(KEYINPUT53), .A3(new_n713), .A4(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1022), .A2(new_n1025), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1104), .A2(new_n1105), .A3(G171), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1105), .B1(new_n1104), .B2(G171), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1026), .A2(G301), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1104), .A2(G171), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1108), .B1(new_n1027), .B2(new_n1112), .ZN(new_n1113));
  AND4_X1   g688(.A1(new_n1016), .A2(new_n1111), .A3(new_n1031), .A4(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1084), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1059), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1098), .B(KEYINPUT114), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT117), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1101), .A2(new_n1114), .A3(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1030), .A2(KEYINPUT124), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1036), .A2(new_n1050), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n722), .B(new_n1053), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(G1996), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(new_n764), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n763), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n698), .B(new_n701), .ZN(new_n1130));
  XOR2_X1   g705(.A(new_n1130), .B(KEYINPUT108), .Z(new_n1131));
  NOR2_X1   g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(G290), .B(G1986), .Z(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1102), .A2(new_n1017), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1123), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1126), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT46), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1135), .B1(new_n1125), .B2(new_n763), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT47), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1135), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1143), .A2(G1986), .A3(G290), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1144), .B(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1143), .B2(new_n1132), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1129), .A2(new_n701), .A3(new_n698), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n722), .A2(G2067), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1135), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1142), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1151), .B(KEYINPUT126), .Z(new_n1152));
  NAND2_X1  g727(.A1(new_n1137), .A2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g728(.A(new_n457), .ZN(new_n1155));
  OR2_X1    g729(.A1(G227), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n1157));
  AND2_X1   g731(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1159));
  NOR3_X1   g733(.A1(G401), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g734(.A(new_n1160), .B1(new_n917), .B2(new_n918), .ZN(new_n1161));
  INV_X1    g735(.A(G229), .ZN(new_n1162));
  NAND2_X1  g736(.A1(new_n845), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g737(.A1(new_n1161), .A2(new_n1163), .ZN(G308));
  INV_X1    g738(.A(new_n918), .ZN(new_n1165));
  NAND3_X1  g739(.A1(new_n905), .A2(new_n916), .A3(new_n910), .ZN(new_n1166));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g741(.A1(new_n1167), .A2(new_n1162), .A3(new_n845), .A4(new_n1160), .ZN(G225));
endmodule


