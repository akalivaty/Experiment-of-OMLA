//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n449, new_n450, new_n453, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n589, new_n590, new_n591, new_n592, new_n594, new_n595, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n636, new_n637,
    new_n638, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G101), .A3(G2104), .ZN(new_n473));
  XOR2_X1   g048(.A(new_n473), .B(KEYINPUT70), .Z(new_n474));
  NAND3_X1  g049(.A1(new_n464), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n475), .A2(new_n467), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n477), .B1(new_n466), .B2(G2104), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n476), .A2(G137), .A3(new_n472), .A4(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n471), .A2(new_n474), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND4_X1  g056(.A1(new_n478), .A2(new_n475), .A3(G2105), .A4(new_n467), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT71), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n476), .A2(new_n472), .A3(new_n478), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G136), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  AND4_X1   g069(.A1(G2105), .A2(new_n478), .A3(new_n475), .A4(new_n467), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G126), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n478), .A2(new_n475), .A3(new_n498), .A4(new_n467), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n465), .A2(new_n467), .ZN(new_n501));
  NOR3_X1   g076(.A1(new_n497), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n496), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n499), .A2(KEYINPUT4), .B1(new_n501), .B2(new_n502), .ZN(new_n507));
  INV_X1    g082(.A(new_n492), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n508), .B1(G114), .B2(new_n472), .ZN(new_n509));
  INV_X1    g084(.A(G126), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n482), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT72), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(KEYINPUT74), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(KEYINPUT5), .A3(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT6), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT73), .B1(new_n524), .B2(G651), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n526), .A2(new_n522), .A3(KEYINPUT6), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(new_n520), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n528), .A2(new_n520), .A3(KEYINPUT75), .A4(new_n529), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n532), .A2(G88), .A3(new_n533), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n528), .A2(G543), .A3(new_n529), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G50), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT76), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n534), .A2(new_n539), .A3(new_n536), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n523), .B1(new_n538), .B2(new_n540), .ZN(G166));
  AND2_X1   g116(.A1(new_n532), .A2(new_n533), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n528), .A2(G51), .A3(G543), .A4(new_n529), .ZN(new_n543));
  AND2_X1   g118(.A1(G63), .A2(G651), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n520), .A2(KEYINPUT77), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(KEYINPUT77), .B1(new_n520), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n542), .A2(G89), .B1(KEYINPUT78), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT78), .ZN(new_n549));
  OAI211_X1 g124(.A(new_n549), .B(new_n543), .C1(new_n545), .C2(new_n546), .ZN(new_n550));
  NAND3_X1  g125(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT7), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(G168));
  NAND2_X1  g130(.A1(new_n542), .A2(G90), .ZN(new_n556));
  NAND2_X1  g131(.A1(G77), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(new_n520), .ZN(new_n558));
  INV_X1    g133(.A(G64), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G651), .B1(new_n535), .B2(G52), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n561), .ZN(G301));
  INV_X1    g137(.A(G301), .ZN(G171));
  NAND2_X1  g138(.A1(new_n542), .A2(G81), .ZN(new_n564));
  NAND2_X1  g139(.A1(G68), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G56), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n558), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n567), .A2(G651), .B1(new_n535), .B2(G43), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(new_n571));
  XOR2_X1   g146(.A(new_n571), .B(KEYINPUT79), .Z(G153));
  NAND4_X1  g147(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND4_X1  g150(.A1(G319), .A2(G483), .A3(G661), .A4(new_n575), .ZN(G188));
  NAND2_X1  g151(.A1(new_n542), .A2(G91), .ZN(new_n577));
  NAND2_X1  g152(.A1(G78), .A2(G543), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT81), .Z(new_n579));
  NAND2_X1  g154(.A1(new_n520), .A2(G65), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n522), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(KEYINPUT80), .A2(KEYINPUT9), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n535), .A2(G53), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n528), .A2(G543), .A3(new_n529), .ZN(new_n584));
  INV_X1    g159(.A(G53), .ZN(new_n585));
  OAI211_X1 g160(.A(KEYINPUT80), .B(KEYINPUT9), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n581), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n577), .A2(new_n587), .ZN(G299));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n548), .A2(new_n553), .A3(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n589), .B1(new_n548), .B2(new_n553), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(G286));
  AND3_X1   g168(.A1(new_n534), .A2(new_n539), .A3(new_n536), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n539), .B1(new_n534), .B2(new_n536), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n594), .A2(new_n595), .B1(new_n522), .B2(new_n521), .ZN(G303));
  OR2_X1    g171(.A1(new_n520), .A2(G74), .ZN(new_n597));
  AOI22_X1  g172(.A1(G49), .A2(new_n535), .B1(new_n597), .B2(G651), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n532), .A2(G87), .A3(new_n533), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(G288));
  NAND2_X1  g175(.A1(G73), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G61), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n558), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(new_n535), .B2(G48), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n532), .A2(G86), .A3(new_n533), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n604), .A2(KEYINPUT83), .A3(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT83), .B1(new_n604), .B2(new_n605), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n607), .A2(new_n608), .ZN(G305));
  NAND2_X1  g184(.A1(G72), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G60), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n558), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT84), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n522), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n613), .B2(new_n612), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n542), .A2(G85), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT85), .B(G47), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n535), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(G290));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NOR2_X1   g195(.A1(G301), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(G79), .A2(G543), .ZN(new_n622));
  INV_X1    g197(.A(G66), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n558), .B2(new_n623), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n624), .A2(G651), .B1(new_n535), .B2(G54), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n542), .A2(KEYINPUT10), .A3(G92), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n532), .A2(new_n533), .ZN(new_n629));
  INV_X1    g204(.A(G92), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n626), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT86), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n621), .B1(new_n633), .B2(new_n620), .ZN(G284));
  AOI21_X1  g209(.A(new_n621), .B1(new_n633), .B2(new_n620), .ZN(G321));
  NOR2_X1   g210(.A1(G299), .A2(G868), .ZN(new_n636));
  INV_X1    g211(.A(new_n592), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(new_n590), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n636), .B1(new_n638), .B2(G868), .ZN(G297));
  AOI21_X1  g214(.A(new_n636), .B1(new_n638), .B2(G868), .ZN(G280));
  INV_X1    g215(.A(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n633), .B1(new_n641), .B2(G860), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT87), .Z(G148));
  INV_X1    g218(.A(KEYINPUT88), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n633), .A2(new_n644), .A3(new_n641), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n627), .A2(new_n631), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(new_n625), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT86), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT86), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n632), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n648), .A2(new_n641), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT88), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n620), .B1(new_n645), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n620), .B2(new_n569), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT89), .Z(G323));
  XNOR2_X1  g230(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g231(.A1(new_n483), .A2(G123), .ZN(new_n657));
  OAI21_X1  g232(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n658));
  INV_X1    g233(.A(G111), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n658), .B1(new_n659), .B2(G2105), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n488), .B2(G135), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT90), .B(G2096), .Z(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT12), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT13), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2100), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n665), .A3(new_n669), .ZN(G156));
  XNOR2_X1  g245(.A(KEYINPUT15), .B(G2435), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2438), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2427), .B(G2430), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(KEYINPUT14), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT91), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(new_n672), .B2(new_n673), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2443), .B(G2446), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1341), .B(G1348), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2451), .B(G2454), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT16), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(G14), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n685), .B2(new_n682), .ZN(G401));
  XNOR2_X1  g262(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n688));
  XNOR2_X1  g263(.A(G2084), .B(G2090), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT92), .ZN(new_n690));
  XNOR2_X1  g265(.A(G2067), .B(G2678), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n688), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT94), .B(KEYINPUT17), .ZN(new_n694));
  INV_X1    g269(.A(new_n690), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(new_n691), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n690), .A2(new_n692), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n688), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G2072), .B(G2078), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n693), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n699), .B2(new_n698), .ZN(new_n701));
  XOR2_X1   g276(.A(G2096), .B(G2100), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT95), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n701), .B(new_n703), .ZN(G227));
  XOR2_X1   g279(.A(G1971), .B(G1976), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT19), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1956), .B(G2474), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1961), .B(G1966), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT96), .Z(new_n712));
  OR2_X1    g287(.A1(new_n708), .A2(new_n709), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT20), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n710), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT97), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(new_n707), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n712), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(G1991), .B(G1996), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(G1981), .B(G1986), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(G229));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NOR2_X1   g302(.A1(G171), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G5), .B2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G1961), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n483), .A2(G129), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n488), .A2(G141), .ZN(new_n733));
  NAND3_X1  g308(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT26), .Z(new_n735));
  NAND3_X1  g310(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n732), .A2(new_n733), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  MUX2_X1   g312(.A(G32), .B(new_n737), .S(G29), .Z(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT27), .B(G1996), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G34), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n742), .B2(KEYINPUT24), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(KEYINPUT24), .B2(new_n742), .ZN(new_n744));
  INV_X1    g319(.A(G29), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n480), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G2084), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n731), .A2(new_n741), .A3(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT102), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n727), .A2(G4), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n633), .B2(new_n727), .ZN(new_n752));
  INV_X1    g327(.A(G1348), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n727), .A2(G20), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT23), .Z(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  INV_X1    g333(.A(G1956), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n745), .A2(G35), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G162), .B2(new_n745), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT29), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n760), .B1(new_n763), .B2(G2090), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n727), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n727), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT101), .B(G1966), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n764), .B(new_n768), .C1(G2090), .C2(new_n763), .ZN(new_n769));
  OAI22_X1  g344(.A1(new_n729), .A2(new_n730), .B1(new_n738), .B2(new_n740), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n745), .A2(G33), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n501), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(new_n472), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT99), .Z(new_n774));
  NAND3_X1  g349(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT25), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n488), .B2(G139), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n771), .B1(new_n778), .B2(G29), .ZN(new_n779));
  INV_X1    g354(.A(G2072), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n746), .A2(new_n747), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n657), .A2(G29), .A3(new_n661), .ZN(new_n783));
  INV_X1    g358(.A(G28), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(KEYINPUT30), .ZN(new_n785));
  AOI21_X1  g360(.A(G29), .B1(new_n784), .B2(KEYINPUT30), .ZN(new_n786));
  OR2_X1    g361(.A1(KEYINPUT31), .A2(G11), .ZN(new_n787));
  NAND2_X1  g362(.A1(KEYINPUT31), .A2(G11), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n785), .A2(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n781), .A2(new_n782), .A3(new_n783), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n745), .A2(G27), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G164), .B2(new_n745), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2078), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n770), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n727), .A2(G19), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n570), .B2(new_n727), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(G1341), .Z(new_n797));
  NOR2_X1   g372(.A1(new_n779), .A2(new_n780), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT100), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n745), .A2(G26), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT28), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n483), .A2(G128), .ZN(new_n802));
  OAI21_X1  g377(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n803));
  INV_X1    g378(.A(G116), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G2105), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n488), .B2(G140), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n801), .B1(new_n807), .B2(G29), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2067), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n794), .A2(new_n797), .A3(new_n799), .A4(new_n809), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n755), .A2(new_n769), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n727), .A2(G22), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G166), .B2(new_n727), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT98), .Z(new_n815));
  INV_X1    g390(.A(G1971), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n727), .A2(G23), .ZN(new_n819));
  INV_X1    g394(.A(G288), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(new_n727), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT33), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1976), .ZN(new_n823));
  MUX2_X1   g398(.A(G6), .B(G305), .S(G16), .Z(new_n824));
  XOR2_X1   g399(.A(KEYINPUT32), .B(G1981), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n817), .A2(new_n818), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(KEYINPUT34), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(KEYINPUT34), .ZN(new_n829));
  INV_X1    g404(.A(G290), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n727), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n727), .B2(G24), .ZN(new_n832));
  INV_X1    g407(.A(G1986), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n745), .A2(G25), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n483), .A2(G119), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n838));
  INV_X1    g413(.A(G107), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(G2105), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n488), .B2(G131), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n836), .B1(new_n843), .B2(new_n745), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT35), .B(G1991), .Z(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n844), .B(new_n846), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n834), .A2(new_n835), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n828), .A2(new_n829), .A3(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n849), .A2(KEYINPUT36), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(KEYINPUT36), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n812), .B1(new_n850), .B2(new_n851), .ZN(G311));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n811), .ZN(G150));
  XOR2_X1   g429(.A(KEYINPUT104), .B(G860), .Z(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT103), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n542), .A2(G93), .ZN(new_n858));
  NAND2_X1  g433(.A1(G80), .A2(G543), .ZN(new_n859));
  INV_X1    g434(.A(G67), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n558), .B2(new_n860), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n861), .A2(G651), .B1(new_n535), .B2(G55), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n857), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G93), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n862), .B1(new_n864), .B2(new_n629), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(KEYINPUT103), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n569), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n569), .B2(new_n865), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n633), .A2(G559), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n856), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n872), .B2(new_n871), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n863), .A2(new_n866), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n856), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT37), .Z(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(G145));
  XNOR2_X1  g453(.A(new_n737), .B(new_n807), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n778), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n507), .A2(new_n511), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT105), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n880), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n488), .A2(G142), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n472), .A2(G118), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(G130), .B2(new_n483), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(new_n667), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n842), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT106), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n883), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n883), .A2(new_n891), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n662), .B(new_n490), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(G160), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n895), .B1(new_n883), .B2(new_n890), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n883), .B2(new_n890), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g476(.A(G303), .B(new_n820), .ZN(new_n902));
  OR3_X1    g477(.A1(new_n607), .A2(KEYINPUT108), .A3(new_n608), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT108), .B1(new_n607), .B2(new_n608), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(G290), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G290), .B1(new_n903), .B2(new_n904), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n903), .A2(new_n904), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n830), .ZN(new_n910));
  XNOR2_X1  g485(.A(G303), .B(G288), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n911), .A3(new_n905), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n914));
  OR2_X1    g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n913), .B1(KEYINPUT109), .B2(KEYINPUT42), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n644), .B1(new_n633), .B2(new_n641), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n651), .A2(KEYINPUT88), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n868), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G299), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n632), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n922), .A2(new_n632), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT41), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n647), .A2(G299), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n929), .A3(new_n923), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n926), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n924), .A2(new_n925), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(KEYINPUT107), .A3(new_n929), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n569), .A2(new_n865), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n875), .B2(new_n569), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n645), .A2(new_n652), .A3(new_n936), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n921), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n932), .B1(new_n921), .B2(new_n937), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n918), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n921), .A2(new_n937), .ZN(new_n941));
  INV_X1    g516(.A(new_n932), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n921), .A2(new_n934), .A3(new_n937), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT110), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n917), .A2(new_n940), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n915), .A2(new_n916), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n947), .A2(KEYINPUT110), .A3(new_n944), .A4(new_n943), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n620), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n875), .A2(G868), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(G295));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n946), .A2(new_n948), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(G868), .ZN(new_n954));
  INV_X1    g529(.A(new_n950), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n949), .A2(KEYINPUT111), .A3(new_n950), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(G331));
  AOI21_X1  g533(.A(G301), .B1(new_n637), .B2(new_n590), .ZN(new_n959));
  NOR2_X1   g534(.A1(G168), .A2(G171), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n936), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n638), .A2(G171), .ZN(new_n962));
  INV_X1    g537(.A(new_n960), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n868), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n932), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n936), .B1(new_n959), .B2(new_n960), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n868), .A3(new_n963), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n931), .A2(new_n966), .A3(new_n967), .A4(new_n933), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n968), .A3(new_n913), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n969), .A2(new_n899), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n965), .A2(new_n968), .ZN(new_n971));
  INV_X1    g546(.A(new_n913), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n966), .A2(new_n967), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n930), .B2(new_n926), .ZN(new_n977));
  INV_X1    g552(.A(new_n965), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n970), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n975), .B1(new_n980), .B2(KEYINPUT43), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n973), .A2(new_n984), .A3(new_n899), .A4(new_n969), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT112), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n970), .A2(new_n987), .A3(new_n984), .A4(new_n973), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n982), .B1(new_n980), .B2(KEYINPUT43), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n989), .A2(new_n990), .A3(KEYINPUT113), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT113), .B1(new_n989), .B2(new_n990), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n983), .B1(new_n991), .B2(new_n992), .ZN(G397));
  NAND2_X1  g568(.A1(new_n807), .A2(G2067), .ZN(new_n994));
  INV_X1    g569(.A(G2067), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n802), .A2(new_n995), .A3(new_n806), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1996), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n737), .B(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n843), .A2(new_n845), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n842), .A2(new_n846), .ZN(new_n1001));
  AND4_X1   g576(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(new_n507), .B2(new_n511), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n471), .A2(new_n474), .A3(new_n479), .A4(G40), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1009), .A2(G290), .A3(G1986), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT127), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1010), .B1(KEYINPUT48), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(KEYINPUT48), .B2(new_n1012), .ZN(new_n1014));
  INV_X1    g589(.A(new_n997), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1008), .B1(new_n1015), .B2(new_n737), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1008), .A2(new_n998), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT46), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1019), .B(KEYINPUT47), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT126), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n999), .A2(new_n997), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n996), .B1(new_n1022), .B2(new_n1000), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n1008), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1014), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1020), .A2(KEYINPUT126), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1004), .A2(KEYINPUT114), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1030), .B(new_n1003), .C1(new_n507), .C2(new_n511), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1007), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1384), .B1(new_n506), .B2(new_n512), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1032), .B(new_n1033), .C1(new_n1029), .C2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1028), .A2(new_n1033), .A3(new_n1031), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1035), .A2(new_n753), .B1(new_n995), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT60), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n632), .B2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1038), .B(new_n1041), .C1(new_n1040), .C2(new_n632), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n632), .A2(new_n1040), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1034), .A2(new_n1029), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n753), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1037), .A2(new_n995), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1043), .B1(new_n1048), .B2(new_n1039), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1046), .A2(new_n1047), .A3(new_n1041), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1042), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT121), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n577), .A2(new_n1053), .A3(new_n587), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n577), .B2(new_n587), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1007), .B1(new_n1034), .B2(new_n1029), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT50), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1956), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT56), .B(G2072), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(KEYINPUT45), .B(new_n1003), .C1(new_n507), .C2(new_n511), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1033), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n513), .A2(new_n1003), .ZN(new_n1065));
  AOI211_X1 g640(.A(new_n1062), .B(new_n1064), .C1(new_n1065), .C2(new_n1005), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1056), .B1(new_n1060), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n505), .B1(new_n496), .B2(new_n504), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n507), .A2(new_n511), .A3(KEYINPUT72), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1029), .B(new_n1003), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1033), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1029), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n759), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1065), .A2(new_n1005), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1384), .B1(new_n496), .B2(new_n504), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1007), .B1(new_n1076), .B2(KEYINPUT45), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(new_n1077), .A3(new_n1061), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1073), .A2(new_n1074), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1067), .A2(KEYINPUT61), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT119), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1067), .A2(new_n1079), .A3(new_n1082), .A4(KEYINPUT61), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1067), .A2(new_n1079), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT61), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT118), .B(G1996), .Z(new_n1087));
  OAI211_X1 g662(.A(new_n1077), .B(new_n1087), .C1(new_n1034), .C2(KEYINPUT45), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT58), .B(G1341), .Z(new_n1089));
  NAND2_X1  g664(.A1(new_n1036), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n569), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1085), .A2(new_n1086), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1096), .B(new_n1042), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1052), .A2(new_n1084), .A3(new_n1095), .A4(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1067), .B1(new_n647), .B2(new_n1038), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n1079), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1071), .A2(G2090), .A3(new_n1072), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1971), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1103));
  OAI21_X1  g678(.A(G8), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT55), .ZN(new_n1105));
  INV_X1    g680(.A(G8), .ZN(new_n1106));
  NOR3_X1   g681(.A1(G166), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1105), .B1(G166), .B2(new_n1106), .ZN(new_n1111));
  NAND3_X1  g686(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1034), .A2(KEYINPUT45), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n816), .B1(new_n1114), .B2(new_n1064), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(G2090), .B2(new_n1035), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1116), .A3(G8), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1036), .A2(G8), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT52), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1119), .B(new_n1120), .C1(new_n820), .C2(G1976), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n820), .A2(G1976), .ZN(new_n1122));
  AOI21_X1  g697(.A(G1976), .B1(new_n598), .B2(new_n599), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT115), .B1(new_n1123), .B2(KEYINPUT52), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1118), .A2(new_n1121), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT49), .ZN(new_n1126));
  INV_X1    g701(.A(G1981), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n604), .A2(new_n1127), .A3(new_n605), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1127), .B1(new_n604), .B2(new_n605), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1126), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1130), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(KEYINPUT49), .A3(new_n1128), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1118), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1122), .A2(G8), .A3(new_n1036), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT52), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1125), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1110), .A2(new_n1117), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT51), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1007), .B1(new_n1058), .B2(new_n1005), .ZN(new_n1140));
  OAI211_X1 g715(.A(KEYINPUT45), .B(new_n1003), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT116), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT116), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1034), .A2(new_n1143), .A3(KEYINPUT45), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n767), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n747), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n554), .A2(G8), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1139), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1150), .B(KEYINPUT122), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1145), .A2(new_n767), .B1(new_n1147), .B2(new_n747), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1154), .B1(new_n1155), .B2(new_n1106), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1154), .B(new_n1139), .C1(new_n1155), .C2(new_n1106), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n730), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1160));
  INV_X1    g735(.A(G2078), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1077), .B(new_n1161), .C1(new_n1034), .C2(KEYINPUT45), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT53), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1163), .A2(G2078), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1077), .A2(new_n1006), .A3(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1160), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1167), .A2(G171), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1035), .A2(new_n730), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1140), .A2(new_n1142), .A3(new_n1144), .A4(new_n1165), .ZN(new_n1170));
  AOI21_X1  g745(.A(G301), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1159), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1138), .A2(new_n1157), .A3(new_n1158), .A4(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1167), .A2(new_n1174), .A3(G171), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1174), .B1(new_n1167), .B2(G171), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT54), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1170), .A2(new_n1160), .A3(new_n1164), .A4(G301), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT123), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1173), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1101), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1137), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1118), .ZN(new_n1184));
  NOR2_X1   g759(.A1(G288), .A2(G1976), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1129), .B1(new_n1134), .B2(new_n1185), .ZN(new_n1186));
  OAI22_X1  g761(.A1(new_n1183), .A2(new_n1117), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT117), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1106), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1189), .B1(new_n1190), .B2(new_n638), .ZN(new_n1191));
  NOR4_X1   g766(.A1(new_n1155), .A2(KEYINPUT117), .A3(new_n1106), .A4(G286), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1117), .A2(new_n1137), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1110), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1188), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1116), .A2(G8), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1188), .B1(new_n1197), .B2(new_n1109), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1194), .B(new_n1198), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1187), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1182), .A2(KEYINPUT125), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(KEYINPUT125), .B1(new_n1182), .B2(new_n1200), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n1204));
  OAI211_X1 g779(.A(new_n1138), .B(new_n1171), .C1(new_n1203), .C2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1205), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1206));
  NOR3_X1   g781(.A1(new_n1201), .A2(new_n1202), .A3(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g782(.A(G290), .B(new_n833), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1009), .B1(new_n1002), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1027), .B1(new_n1207), .B2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g785(.A(new_n461), .ZN(new_n1212));
  NOR4_X1   g786(.A1(G229), .A2(G401), .A3(new_n1212), .A4(G227), .ZN(new_n1213));
  NAND3_X1  g787(.A1(new_n1213), .A2(new_n900), .A3(new_n981), .ZN(G225));
  INV_X1    g788(.A(G225), .ZN(G308));
endmodule


