//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT77), .A2(KEYINPUT12), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT76), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT76), .A2(G104), .ZN(new_n193));
  AOI21_X1  g007(.A(G107), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G104), .ZN(new_n196));
  OAI21_X1  g010(.A(G101), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  NOR3_X1   g011(.A1(new_n191), .A2(KEYINPUT3), .A3(G107), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n194), .B2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n192), .A2(G107), .A3(new_n193), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n197), .B1(new_n201), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT1), .B1(new_n206), .B2(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  OAI211_X1 g024(.A(G128), .B(new_n207), .C1(new_n208), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n206), .A2(G146), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n212), .B(new_n213), .C1(KEYINPUT1), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n205), .A2(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT76), .A2(G104), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT76), .A2(G104), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(G101), .B1(new_n220), .B2(G107), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n195), .B1(new_n218), .B2(new_n219), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT3), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(new_n223), .A3(new_n199), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n211), .A2(new_n215), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(new_n197), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n217), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT11), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(G137), .ZN(new_n230));
  INV_X1    g044(.A(G137), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT11), .A3(G134), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(G137), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G131), .ZN(new_n235));
  INV_X1    g049(.A(G131), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n230), .A2(new_n232), .A3(new_n236), .A4(new_n233), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT77), .A2(KEYINPUT12), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n189), .B1(new_n227), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n189), .ZN(new_n244));
  AOI211_X1 g058(.A(new_n241), .B(new_n244), .C1(new_n217), .C2(new_n226), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G143), .B(G146), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT0), .A3(G128), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT0), .B(G128), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n202), .B(new_n199), .C1(new_n194), .C2(new_n200), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G101), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n252), .B1(new_n254), .B2(new_n224), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n198), .B1(new_n222), .B2(KEYINPUT3), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n203), .B1(new_n256), .B2(new_n202), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT4), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n251), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n238), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT10), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n226), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n222), .B1(G104), .B2(new_n195), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n256), .A2(new_n221), .B1(new_n263), .B2(G101), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT10), .A3(new_n225), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n259), .A2(new_n260), .A3(new_n262), .A4(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G110), .B(G140), .ZN(new_n267));
  INV_X1    g081(.A(G953), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n268), .A2(G227), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n267), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n246), .A2(new_n266), .A3(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n201), .A2(new_n204), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT4), .B1(new_n257), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n254), .A2(new_n252), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n250), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n262), .A2(new_n265), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n238), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n271), .B1(new_n278), .B2(new_n266), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n272), .B1(new_n279), .B2(KEYINPUT79), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n272), .A2(KEYINPUT79), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n187), .B(new_n188), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n187), .A2(new_n188), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT78), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n278), .A2(new_n266), .A3(new_n271), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n271), .B1(new_n246), .B2(new_n266), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n286), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n276), .A2(new_n277), .A3(new_n238), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n224), .A2(new_n225), .A3(new_n197), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n224), .A2(new_n197), .B1(new_n215), .B2(new_n211), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n242), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n244), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n227), .A2(new_n242), .A3(new_n189), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n270), .B1(new_n291), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(KEYINPUT78), .A3(new_n287), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n290), .A2(G469), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n283), .A2(new_n285), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT9), .B(G234), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(KEYINPUT75), .ZN(new_n303));
  OAI21_X1  g117(.A(G221), .B1(new_n303), .B2(G902), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G210), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(G125), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n216), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n308), .B1(new_n251), .B2(new_n307), .ZN(new_n309));
  INV_X1    g123(.A(G224), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(G953), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n309), .B(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(G116), .B(G119), .Z(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT2), .B(G113), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G113), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT81), .B(KEYINPUT5), .Z(new_n317));
  INV_X1    g131(.A(G116), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(G119), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n316), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(new_n313), .B2(new_n317), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n264), .A2(new_n315), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G110), .B(G122), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n255), .A2(new_n258), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n313), .B(new_n314), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n322), .B(new_n323), .C1(new_n324), .C2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n322), .B1(new_n324), .B2(new_n326), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n323), .B(KEYINPUT82), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n327), .A2(KEYINPUT6), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n328), .A2(KEYINPUT6), .A3(new_n329), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n312), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT7), .B1(new_n310), .B2(G953), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n309), .B(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n205), .A2(new_n315), .A3(new_n321), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n323), .B(KEYINPUT8), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT83), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT5), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n320), .B1(new_n339), .B2(new_n313), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n205), .B1(new_n315), .B2(new_n340), .ZN(new_n341));
  OR3_X1    g155(.A1(new_n337), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n338), .B1(new_n337), .B2(new_n341), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n334), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(G902), .B1(new_n344), .B2(new_n327), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n306), .B1(new_n332), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n332), .A2(new_n345), .A3(new_n306), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(G214), .B1(G237), .B2(G902), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n350), .B(KEYINPUT80), .Z(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT66), .B(G237), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(G214), .A3(new_n268), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n206), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n355), .A2(G143), .A3(G214), .A4(new_n268), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT18), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(new_n236), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT84), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n359), .A2(KEYINPUT84), .A3(new_n361), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G140), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G125), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n307), .A2(G140), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n368), .A2(new_n369), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT85), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(G146), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n370), .A2(new_n209), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(KEYINPUT86), .A3(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n357), .B(new_n358), .C1(new_n360), .C2(new_n236), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT86), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n372), .A2(new_n379), .A3(G146), .A4(new_n374), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n366), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G113), .B(G122), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(new_n191), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n370), .A2(KEYINPUT16), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n368), .A2(KEYINPUT16), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n386), .A2(G146), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(G146), .B1(new_n386), .B2(new_n387), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n359), .A2(KEYINPUT17), .A3(G131), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT88), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n236), .B1(new_n357), .B2(new_n358), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT17), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n357), .A2(new_n236), .A3(new_n358), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT88), .B1(new_n390), .B2(new_n391), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n383), .B(new_n385), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n385), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n381), .B1(new_n364), .B2(new_n365), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n386), .A2(G146), .A3(new_n387), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n372), .A2(KEYINPUT19), .A3(new_n374), .ZN(new_n404));
  OR2_X1    g218(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n370), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n403), .B1(new_n408), .B2(G146), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n394), .B2(new_n396), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n401), .B1(new_n402), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n400), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(G475), .A2(G902), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n354), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n413), .ZN(new_n415));
  AOI211_X1 g229(.A(KEYINPUT20), .B(new_n415), .C1(new_n400), .C2(new_n411), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n383), .B1(new_n398), .B2(new_n399), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n401), .ZN(new_n418));
  AOI21_X1  g232(.A(G902), .B1(new_n418), .B2(new_n400), .ZN(new_n419));
  XOR2_X1   g233(.A(KEYINPUT89), .B(G475), .Z(new_n420));
  OAI22_X1  g234(.A1(new_n414), .A2(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G478), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(KEYINPUT15), .ZN(new_n424));
  INV_X1    g238(.A(G217), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n303), .A2(new_n425), .A3(G953), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n214), .A2(G143), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT13), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n229), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G128), .B(G143), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G122), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n433), .A2(KEYINPUT90), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(KEYINPUT90), .ZN(new_n435));
  OAI21_X1  g249(.A(G116), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n318), .A2(G122), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n195), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n195), .B1(new_n436), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n432), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT90), .B(G122), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(new_n318), .ZN(new_n443));
  OR3_X1    g257(.A1(new_n433), .A2(KEYINPUT14), .A3(G116), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n437), .A2(KEYINPUT14), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G107), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n431), .B(new_n229), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n438), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT91), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n441), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n450), .B1(new_n441), .B2(new_n449), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n427), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n453), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n426), .A3(new_n451), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n456), .A3(new_n188), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT92), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n424), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n458), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n454), .A2(new_n456), .A3(KEYINPUT92), .A4(new_n188), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n459), .B1(new_n462), .B2(new_n424), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n268), .A2(G952), .ZN(new_n464));
  NAND2_X1  g278(.A1(G234), .A2(G237), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(G898), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(G902), .A3(G953), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n422), .A2(new_n463), .A3(new_n470), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n305), .A2(new_n353), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n355), .A2(G210), .A3(new_n268), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT27), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT26), .B(G101), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT69), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n229), .A2(G137), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n231), .A2(G134), .ZN(new_n480));
  OAI21_X1  g294(.A(G131), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n211), .A2(new_n237), .A3(new_n481), .A4(new_n215), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT64), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n251), .A2(new_n238), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n483), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n325), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n482), .B(KEYINPUT65), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n325), .B1(new_n251), .B2(new_n238), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT28), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n490), .A2(new_n482), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n494), .A2(KEYINPUT28), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n478), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT69), .B1(new_n492), .B2(KEYINPUT28), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n477), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT67), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n487), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n489), .A2(KEYINPUT30), .A3(new_n485), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n325), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n491), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n499), .B1(new_n504), .B2(new_n477), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n503), .A2(KEYINPUT67), .A3(new_n476), .A4(new_n491), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(KEYINPUT31), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n504), .A2(new_n477), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT31), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT68), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT68), .ZN(new_n511));
  NOR4_X1   g325(.A1(new_n504), .A2(new_n511), .A3(KEYINPUT31), .A4(new_n477), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n498), .B(new_n507), .C1(new_n510), .C2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(G472), .A2(G902), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(KEYINPUT32), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT70), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n514), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT32), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n494), .A2(KEYINPUT28), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n489), .A2(new_n485), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n491), .B1(new_n522), .B2(new_n326), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n523), .B2(KEYINPUT28), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT29), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n477), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(G902), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n496), .A2(new_n477), .A3(new_n497), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n504), .A2(new_n477), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n525), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n527), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G472), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n513), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n514), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n517), .A2(new_n520), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G119), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G128), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT71), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(KEYINPUT71), .A3(G128), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n538), .B(new_n539), .C1(new_n535), .C2(G128), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT24), .B(G110), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n214), .A2(KEYINPUT23), .A3(G119), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n535), .A2(G128), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n543), .B(new_n536), .C1(new_n544), .C2(KEYINPUT23), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n542), .B1(G110), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n403), .A3(new_n376), .ZN(new_n547));
  OAI22_X1  g361(.A1(new_n388), .A2(new_n389), .B1(new_n541), .B2(new_n540), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n545), .A2(G110), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT72), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n547), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT22), .B(G137), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n268), .A2(G221), .A3(G234), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT73), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n547), .B(new_n554), .C1(new_n548), .C2(new_n550), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n188), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT25), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n556), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n557), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n425), .B1(G234), .B2(new_n188), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(G902), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT74), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n556), .A2(new_n557), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n472), .A2(new_n534), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(G101), .ZN(G3));
  NAND2_X1  g385(.A1(new_n513), .A2(new_n188), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n572), .A2(G472), .B1(new_n513), .B2(new_n514), .ZN(new_n573));
  INV_X1    g387(.A(new_n304), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n272), .A2(KEYINPUT79), .ZN(new_n575));
  AOI21_X1  g389(.A(G902), .B1(new_n575), .B2(new_n280), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n284), .B1(new_n576), .B2(new_n187), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n574), .B1(new_n577), .B2(new_n300), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n573), .A2(new_n569), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n412), .A2(new_n413), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT20), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n412), .A2(new_n354), .A3(new_n413), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n418), .A2(new_n400), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n188), .ZN(new_n585));
  INV_X1    g399(.A(new_n420), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n457), .A2(new_n423), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n454), .A2(new_n456), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n441), .A2(new_n449), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT93), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT33), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n454), .A2(KEYINPUT33), .A3(new_n456), .A4(new_n591), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n423), .A2(G902), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n583), .A2(new_n587), .B1(new_n588), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n598), .A2(new_n470), .ZN(new_n599));
  INV_X1    g413(.A(new_n350), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n347), .B2(new_n348), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n579), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT34), .B(G104), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G6));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n585), .A2(new_n605), .A3(new_n586), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT94), .B1(new_n419), .B2(new_n420), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n463), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n609), .A3(new_n583), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n470), .B(KEYINPUT95), .Z(new_n611));
  INV_X1    g425(.A(new_n348), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n350), .B(new_n611), .C1(new_n612), .C2(new_n346), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n579), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT35), .B(G107), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G9));
  NAND2_X1  g431(.A1(new_n572), .A2(G472), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n555), .A2(KEYINPUT36), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(new_n551), .Z(new_n620));
  INV_X1    g434(.A(new_n566), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n564), .A2(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n618), .A2(new_n518), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n472), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT37), .B(G110), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G12));
  NAND2_X1  g441(.A1(new_n349), .A2(new_n350), .ZN(new_n628));
  INV_X1    g442(.A(new_n623), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n534), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n606), .A2(new_n607), .B1(new_n581), .B2(new_n582), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n466), .B1(G900), .B2(new_n469), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n609), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n305), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G128), .ZN(G30));
  NAND3_X1  g451(.A1(new_n609), .A2(new_n421), .A3(new_n350), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n612), .A2(new_n346), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT38), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n633), .B(KEYINPUT39), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n578), .A2(new_n641), .ZN(new_n642));
  AOI211_X1 g456(.A(new_n638), .B(new_n640), .C1(KEYINPUT40), .C2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n505), .A2(new_n506), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n477), .B2(new_n523), .ZN(new_n645));
  OAI21_X1  g459(.A(G472), .B1(new_n645), .B2(G902), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n517), .A2(new_n520), .A3(new_n533), .A4(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n623), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n643), .B(new_n649), .C1(KEYINPUT40), .C2(new_n642), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G143), .ZN(G45));
  NAND2_X1  g465(.A1(new_n597), .A2(new_n588), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n421), .A2(new_n652), .A3(new_n633), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n305), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n631), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G146), .ZN(G48));
  NOR2_X1   g471(.A1(new_n281), .A2(new_n282), .ZN(new_n658));
  OAI21_X1  g472(.A(G469), .B1(new_n658), .B2(G902), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n304), .A3(new_n283), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n628), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n534), .A2(new_n661), .A3(new_n569), .A4(new_n599), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT41), .B(G113), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT96), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n662), .B(new_n664), .ZN(G15));
  NOR3_X1   g479(.A1(new_n660), .A2(new_n613), .A3(new_n610), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n534), .A3(new_n569), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT97), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n666), .A2(new_n534), .A3(KEYINPUT97), .A4(new_n569), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G116), .ZN(G18));
  NOR2_X1   g486(.A1(new_n660), .A2(new_n471), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n534), .A2(new_n630), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G119), .ZN(G21));
  OAI221_X1 g489(.A(new_n507), .B1(new_n476), .B2(new_n524), .C1(new_n510), .C2(new_n512), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n514), .B(KEYINPUT98), .Z(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n618), .A2(new_n569), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n611), .ZN(new_n680));
  OAI21_X1  g494(.A(KEYINPUT99), .B1(new_n422), .B2(new_n463), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT99), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n609), .A2(new_n682), .A3(new_n421), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n680), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n679), .A2(new_n661), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G122), .ZN(G24));
  AND4_X1   g500(.A1(new_n618), .A2(new_n623), .A3(new_n653), .A4(new_n678), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT100), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n688), .A3(new_n661), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n618), .A2(new_n623), .A3(new_n653), .A4(new_n678), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n601), .A2(new_n304), .A3(new_n283), .A4(new_n659), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT100), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  AND2_X1   g508(.A1(new_n534), .A2(new_n569), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n298), .A2(new_n287), .ZN(new_n696));
  OR3_X1    g510(.A1(new_n696), .A2(KEYINPUT101), .A3(new_n187), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT101), .B1(new_n696), .B2(new_n187), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n574), .B1(new_n699), .B2(new_n577), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT102), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n639), .A2(new_n350), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n283), .A2(new_n698), .A3(new_n285), .A4(new_n697), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n304), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n695), .A2(new_n701), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n701), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n518), .A2(new_n519), .B1(G472), .B2(new_n531), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n515), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n569), .A3(new_n653), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT42), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n236), .ZN(G33));
  NAND4_X1  g529(.A1(new_n706), .A2(new_n534), .A3(new_n701), .A4(new_n569), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n634), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT103), .B(G134), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G36));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n696), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n290), .A2(new_n299), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n187), .B1(new_n723), .B2(new_n721), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n722), .B1(new_n724), .B2(KEYINPUT104), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT45), .B1(new_n290), .B2(new_n299), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n726), .B1(new_n727), .B2(new_n187), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT105), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n298), .A2(KEYINPUT78), .A3(new_n287), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT78), .B1(new_n298), .B2(new_n287), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n721), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(KEYINPUT104), .A3(G469), .ZN(new_n733));
  INV_X1    g547(.A(new_n722), .ZN(new_n734));
  AND4_X1   g548(.A1(KEYINPUT105), .A2(new_n728), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  OAI211_X1 g549(.A(KEYINPUT46), .B(new_n285), .C1(new_n729), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n283), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT106), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n728), .A2(new_n733), .A3(new_n734), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n725), .A2(KEYINPUT105), .A3(new_n728), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n284), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n738), .B1(new_n743), .B2(KEYINPUT46), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n285), .B1(new_n729), .B2(new_n735), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(KEYINPUT106), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n737), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n641), .A2(new_n304), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n720), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n736), .A2(new_n283), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n743), .A2(new_n738), .A3(KEYINPUT46), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT106), .B1(new_n745), .B2(new_n746), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n749), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(KEYINPUT107), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n702), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n421), .A2(KEYINPUT108), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n421), .A2(KEYINPUT108), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n758), .A2(KEYINPUT43), .A3(new_n652), .A4(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n421), .B1(new_n588), .B2(new_n597), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n760), .B1(KEYINPUT43), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n573), .A2(new_n629), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n757), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n764), .B2(new_n765), .ZN(new_n768));
  AOI211_X1 g582(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n762), .C2(new_n763), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n750), .A2(new_n756), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  OAI21_X1  g586(.A(KEYINPUT47), .B1(new_n748), .B2(new_n574), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n754), .A2(new_n774), .A3(new_n304), .ZN(new_n775));
  NOR4_X1   g589(.A1(new_n534), .A2(new_n569), .A3(new_n654), .A4(new_n702), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT110), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n773), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(KEYINPUT111), .B(G140), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G42));
  INV_X1    g594(.A(new_n660), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n640), .A2(new_n781), .A3(new_n600), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT117), .ZN(new_n783));
  AND4_X1   g597(.A1(new_n465), .A2(new_n762), .A3(new_n464), .A4(new_n679), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT50), .Z(new_n786));
  NOR3_X1   g600(.A1(new_n660), .A2(new_n702), .A3(new_n466), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n787), .A2(new_n569), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n648), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n789), .A2(new_n421), .A3(new_n652), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT118), .Z(new_n791));
  AND3_X1   g605(.A1(new_n618), .A2(new_n623), .A3(new_n678), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n762), .A2(new_n787), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n786), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n659), .A2(new_n283), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT112), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n773), .A2(new_n775), .B1(new_n574), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n784), .A2(new_n757), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n794), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n800), .B1(new_n794), .B2(new_n799), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n568), .B1(new_n710), .B2(new_n515), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n762), .A2(new_n787), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n804), .A2(new_n805), .A3(KEYINPUT48), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n784), .A2(new_n661), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n788), .A2(new_n598), .A3(new_n648), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n808), .A3(new_n464), .ZN(new_n809));
  XNOR2_X1  g623(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n810));
  AOI211_X1 g624(.A(new_n806), .B(new_n809), .C1(new_n804), .C2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n801), .A2(new_n802), .A3(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n662), .A2(new_n685), .A3(new_n674), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n671), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n708), .A2(new_n713), .A3(KEYINPUT53), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n421), .A2(new_n463), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n598), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n349), .A2(new_n352), .A3(new_n611), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n579), .A2(new_n820), .B1(new_n472), .B2(new_n624), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n463), .A2(new_n623), .A3(new_n633), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(new_n632), .A3(new_n639), .A4(new_n350), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n305), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n825), .A3(new_n534), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n825), .B1(new_n824), .B2(new_n534), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n821), .B(new_n570), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  OAI22_X1  g643(.A1(new_n716), .A2(new_n634), .B1(new_n709), .B2(new_n690), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT116), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n816), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n700), .A2(new_n633), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n628), .B1(new_n681), .B2(new_n683), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n647), .A3(new_n629), .A4(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n534), .B(new_n630), .C1(new_n655), .C2(new_n635), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n688), .B1(new_n687), .B2(new_n661), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n690), .A2(new_n691), .A3(KEYINPUT100), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n693), .A2(KEYINPUT52), .A3(new_n836), .A4(new_n835), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT115), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT115), .B1(new_n841), .B2(new_n842), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n687), .A2(new_n706), .A3(new_n701), .ZN(new_n847));
  INV_X1    g661(.A(new_n716), .ZN(new_n848));
  INV_X1    g662(.A(new_n634), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n305), .A2(new_n568), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n820), .A2(new_n852), .A3(new_n573), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n570), .A2(new_n853), .A3(new_n625), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n828), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n826), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n850), .A2(new_n851), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n832), .A2(new_n844), .A3(new_n846), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT113), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n671), .A2(new_n813), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n860), .B1(new_n671), .B2(new_n813), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n803), .A2(new_n706), .A3(new_n653), .A4(new_n701), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n848), .A2(new_n707), .B1(new_n864), .B2(KEYINPUT42), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(new_n850), .A3(new_n855), .A4(new_n857), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n841), .A2(new_n842), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n863), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n859), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n869), .A2(KEYINPUT53), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n866), .A2(new_n861), .A3(new_n862), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n870), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n844), .A2(new_n846), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n873), .B1(new_n878), .B2(new_n872), .ZN(new_n879));
  OAI22_X1  g693(.A1(new_n812), .A2(new_n879), .B1(G952), .B2(G953), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n796), .B(KEYINPUT49), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n569), .A2(new_n304), .A3(new_n652), .A4(new_n352), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n640), .A2(new_n759), .A3(new_n758), .A4(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n648), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n880), .A2(new_n884), .ZN(G75));
  NOR2_X1   g699(.A1(new_n268), .A2(G952), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n188), .B1(new_n859), .B2(new_n871), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT56), .B1(new_n888), .B2(G210), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n330), .A2(new_n331), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(new_n312), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT55), .Z(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n887), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n889), .B2(new_n893), .ZN(G51));
  NOR2_X1   g709(.A1(new_n729), .A2(new_n735), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT53), .B1(new_n875), .B2(new_n868), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n816), .A2(new_n858), .A3(new_n831), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n898), .A2(new_n845), .A3(new_n843), .ZN(new_n899));
  OAI211_X1 g713(.A(G902), .B(new_n896), .C1(new_n897), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT121), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n859), .A2(new_n871), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n902), .A2(new_n903), .A3(G902), .A4(new_n896), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT54), .B1(new_n897), .B2(new_n899), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n873), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n284), .B(KEYINPUT57), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n658), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n905), .B1(new_n909), .B2(KEYINPUT120), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n911));
  INV_X1    g725(.A(new_n908), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n906), .B2(new_n873), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n911), .B1(new_n913), .B2(new_n658), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n886), .B1(new_n910), .B2(new_n914), .ZN(G54));
  NAND3_X1  g729(.A1(new_n888), .A2(KEYINPUT58), .A3(G475), .ZN(new_n916));
  INV_X1    g730(.A(new_n412), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n886), .ZN(G60));
  NAND2_X1  g734(.A1(G478), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT59), .Z(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n907), .A2(new_n595), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n595), .B1(new_n879), .B2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n886), .ZN(G63));
  XNOR2_X1  g740(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n425), .A2(new_n188), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n902), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n567), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n902), .A2(new_n620), .A3(new_n929), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n887), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G66));
  AOI21_X1  g749(.A(new_n268), .B1(new_n468), .B2(G224), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n863), .A2(new_n855), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT123), .Z(new_n938));
  AOI21_X1  g752(.A(new_n936), .B1(new_n938), .B2(new_n268), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n890), .B1(G898), .B2(new_n268), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n939), .B(new_n940), .Z(G69));
  AOI21_X1  g755(.A(new_n268), .B1(G227), .B2(G900), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n408), .B(KEYINPUT124), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT125), .Z(new_n944));
  NAND2_X1  g758(.A1(new_n501), .A2(new_n502), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n944), .B(new_n945), .Z(new_n946));
  AND2_X1   g760(.A1(new_n803), .A2(new_n834), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n750), .A2(new_n756), .A3(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n778), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n693), .A2(new_n836), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n714), .A2(new_n950), .A3(new_n717), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n771), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(G953), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n268), .A2(G900), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT126), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n771), .A2(new_n778), .A3(new_n948), .A4(new_n951), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n268), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n958));
  INV_X1    g772(.A(new_n954), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n946), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n650), .A2(new_n693), .A3(new_n836), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT62), .Z(new_n963));
  NOR3_X1   g777(.A1(new_n642), .A2(new_n702), .A3(new_n818), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n695), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n963), .A2(new_n771), .A3(new_n778), .A4(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n966), .A2(new_n268), .ZN(new_n967));
  INV_X1    g781(.A(new_n946), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n942), .B1(new_n961), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n958), .B1(new_n957), .B2(new_n959), .ZN(new_n971));
  AOI211_X1 g785(.A(KEYINPUT126), .B(new_n954), .C1(new_n956), .C2(new_n268), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n942), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n973), .B(new_n974), .C1(new_n967), .C2(new_n968), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n970), .A2(new_n975), .ZN(G72));
  XNOR2_X1  g790(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n977));
  NAND2_X1  g791(.A1(G472), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n938), .B2(new_n956), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n981), .A2(new_n477), .A3(new_n491), .A4(new_n503), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n980), .B1(new_n938), .B2(new_n966), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n983), .A2(new_n476), .A3(new_n504), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n644), .B1(new_n477), .B2(new_n504), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n878), .A2(new_n979), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n986), .A2(new_n886), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n982), .A2(new_n984), .A3(new_n987), .ZN(G57));
endmodule


