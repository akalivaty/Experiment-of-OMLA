//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906;
  INV_X1    g000(.A(G120gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT1), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI211_X1 g007(.A(KEYINPUT1), .B(G134gat), .C1(new_n203), .C2(new_n205), .ZN(new_n209));
  OAI21_X1  g008(.A(G127gat), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G134gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G127gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n212), .B(new_n213), .C1(new_n206), .C2(new_n207), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT27), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT27), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G183gat), .ZN(new_n220));
  INV_X1    g019(.A(G190gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n222), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT66), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n225), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n218), .A2(new_n220), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT28), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n236), .A3(new_n221), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n223), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n231), .A2(KEYINPUT23), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n239), .A2(new_n224), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(G183gat), .A2(G190gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n245), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT25), .B1(new_n242), .B2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n239), .A2(KEYINPUT25), .A3(new_n241), .A4(new_n224), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n217), .A2(new_n221), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n253), .A2(new_n247), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT24), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n255), .A2(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(KEYINPUT65), .B2(new_n255), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n252), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n238), .B(KEYINPUT68), .C1(new_n251), .C2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n244), .B1(new_n261), .B2(KEYINPUT24), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n255), .A2(KEYINPUT65), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n247), .B(new_n253), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n242), .A2(new_n264), .A3(KEYINPUT25), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n239), .A2(new_n224), .A3(new_n241), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n243), .A2(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(new_n246), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n265), .B1(new_n268), .B2(KEYINPUT25), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT68), .B1(new_n269), .B2(new_n238), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n216), .B1(new_n260), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G227gat), .A2(G233gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n238), .B1(new_n251), .B2(new_n258), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n215), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n271), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT34), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT34), .B1(new_n277), .B2(new_n278), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT72), .ZN(new_n281));
  INV_X1    g080(.A(new_n272), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n215), .B1(new_n275), .B2(new_n259), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n270), .A2(new_n216), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT69), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n287), .B(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT33), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT32), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n290), .B1(new_n286), .B2(new_n288), .ZN(new_n291));
  XNOR2_X1  g090(.A(G15gat), .B(G43gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT70), .ZN(new_n293));
  XNOR2_X1  g092(.A(G71gat), .B(G99gat), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n293), .B(new_n294), .Z(new_n295));
  NOR3_X1   g094(.A1(new_n289), .A2(new_n291), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n295), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT33), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n285), .A2(KEYINPUT69), .ZN(new_n299));
  INV_X1    g098(.A(new_n288), .ZN(new_n300));
  OAI211_X1 g099(.A(KEYINPUT32), .B(new_n298), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT72), .B1(new_n279), .B2(new_n280), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n281), .B1(new_n296), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n289), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT32), .B1(new_n299), .B2(new_n300), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n306), .A3(new_n297), .ZN(new_n307));
  INV_X1    g106(.A(new_n281), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n301), .A4(new_n302), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G8gat), .B(G36gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(G64gat), .B(G92gat), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n311), .B(new_n312), .Z(new_n313));
  XNOR2_X1  g112(.A(G211gat), .B(G218gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(G197gat), .B(G204gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT22), .ZN(new_n316));
  INV_X1    g115(.A(G211gat), .ZN(new_n317));
  INV_X1    g116(.A(G218gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n314), .A2(new_n315), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n314), .B1(new_n319), .B2(new_n315), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G226gat), .ZN(new_n324));
  INV_X1    g123(.A(G233gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n273), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n269), .A2(KEYINPUT73), .A3(new_n238), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n327), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n326), .A2(KEYINPUT29), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n273), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n323), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n269), .A2(new_n326), .A3(new_n238), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n336), .A3(new_n322), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n313), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n334), .A2(new_n337), .A3(new_n313), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n334), .A2(KEYINPUT30), .A3(new_n337), .A4(new_n313), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n342), .A2(new_n343), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n341), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G141gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G148gat), .ZN(new_n348));
  INV_X1    g147(.A(G148gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G141gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n348), .A2(new_n350), .B1(KEYINPUT2), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n353));
  INV_X1    g152(.A(new_n351), .ZN(new_n354));
  NOR2_X1   g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G155gat), .ZN(new_n357));
  INV_X1    g156(.A(G162gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(KEYINPUT75), .A3(new_n351), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n352), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G155gat), .B(G162gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G141gat), .B(G148gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT2), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(G155gat), .B2(G162gat), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n353), .B(new_n362), .C1(new_n363), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n215), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT4), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n215), .A2(new_n370), .A3(new_n367), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n367), .A2(KEYINPUT76), .A3(new_n372), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n210), .B(new_n214), .C1(new_n367), .C2(new_n372), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n369), .A2(new_n371), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n381));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT76), .B1(new_n367), .B2(new_n372), .ZN(new_n386));
  AOI211_X1 g185(.A(new_n374), .B(KEYINPUT3), .C1(new_n361), .C2(new_n366), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n382), .B1(new_n388), .B2(new_n378), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n370), .B1(new_n215), .B2(new_n367), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT77), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(new_n371), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n215), .A2(KEYINPUT77), .A3(new_n370), .A4(new_n367), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n395));
  INV_X1    g194(.A(new_n367), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(new_n210), .A3(new_n214), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n368), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n216), .A2(KEYINPUT78), .A3(new_n396), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n383), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n381), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n385), .B1(new_n394), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G1gat), .B(G29gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT0), .ZN(new_n404));
  XNOR2_X1  g203(.A(G57gat), .B(G85gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(KEYINPUT6), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n402), .A2(new_n407), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n406), .B(new_n385), .C1(new_n394), .C2(new_n401), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n346), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT29), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n414), .B1(new_n386), .B2(new_n387), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n322), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n414), .B1(new_n320), .B2(new_n321), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n367), .B1(new_n417), .B2(new_n372), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(G228gat), .A2(G233gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(G22gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n421), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n416), .A2(new_n424), .A3(new_n419), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT80), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n424), .B1(new_n416), .B2(new_n419), .ZN(new_n428));
  AOI211_X1 g227(.A(new_n421), .B(new_n418), .C1(new_n415), .C2(new_n322), .ZN(new_n429));
  OAI21_X1  g228(.A(G22gat), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT81), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT81), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n432), .B(G22gat), .C1(new_n428), .C2(new_n429), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT80), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n422), .A2(new_n434), .A3(new_n423), .A4(new_n425), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n427), .A2(new_n431), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G78gat), .B(G106gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT31), .B(G50gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT83), .ZN(new_n441));
  INV_X1    g240(.A(new_n439), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n430), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT82), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT82), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n426), .A2(new_n430), .A3(new_n445), .A4(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n440), .A2(new_n441), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n441), .B1(new_n440), .B2(new_n447), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n310), .B(new_n413), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT35), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n440), .A2(new_n447), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT83), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n440), .A2(new_n441), .A3(new_n447), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT86), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT35), .B1(new_n413), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n346), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n412), .A2(new_n408), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT86), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n455), .A2(new_n310), .A3(new_n457), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n451), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n371), .A2(new_n391), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n464), .A2(new_n393), .A3(new_n369), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n400), .B(new_n381), .C1(new_n465), .C2(new_n389), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n406), .B1(new_n466), .B2(new_n385), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n380), .A2(new_n382), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT39), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n407), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n383), .B1(new_n398), .B2(new_n399), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(KEYINPUT84), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT39), .B1(new_n380), .B2(new_n382), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT40), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n467), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n470), .B(KEYINPUT40), .C1(new_n472), .C2(new_n473), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n476), .A2(new_n346), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n459), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n334), .A2(new_n337), .ZN(new_n481));
  INV_X1    g280(.A(new_n313), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(KEYINPUT37), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n483), .A2(new_n484), .B1(KEYINPUT37), .B2(new_n481), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT38), .ZN(new_n487));
  OR3_X1    g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n486), .B1(new_n485), .B2(new_n487), .ZN(new_n489));
  INV_X1    g288(.A(new_n340), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n483), .A2(new_n484), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT37), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n335), .A2(new_n336), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(new_n323), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n322), .B1(new_n331), .B2(new_n333), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT38), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n490), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n480), .A2(new_n488), .A3(new_n489), .A4(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n479), .B(new_n498), .C1(new_n449), .C2(new_n448), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n448), .A2(new_n449), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n460), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n304), .A2(KEYINPUT36), .A3(new_n309), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT36), .B1(new_n304), .B2(new_n309), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n499), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n463), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g305(.A1(KEYINPUT87), .A2(KEYINPUT14), .ZN(new_n507));
  NOR2_X1   g306(.A1(KEYINPUT87), .A2(KEYINPUT14), .ZN(new_n508));
  OAI22_X1  g307(.A1(new_n507), .A2(new_n508), .B1(G29gat), .B2(G36gat), .ZN(new_n509));
  OR2_X1    g308(.A1(G29gat), .A2(G36gat), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(new_n510), .B2(new_n507), .ZN(new_n511));
  NAND2_X1  g310(.A1(G29gat), .A2(G36gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G43gat), .B(G50gat), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n515), .A2(KEYINPUT88), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(KEYINPUT88), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n514), .A2(KEYINPUT15), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n512), .B(KEYINPUT90), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n511), .B(KEYINPUT89), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT17), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT16), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(KEYINPUT91), .ZN(new_n528));
  INV_X1    g327(.A(G1gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n525), .B(KEYINPUT91), .C1(new_n526), .C2(G1gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G8gat), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT92), .Z(new_n534));
  NOR2_X1   g333(.A1(new_n532), .A2(G8gat), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n535), .B(KEYINPUT93), .Z(new_n536));
  NAND3_X1  g335(.A1(new_n524), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n534), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n523), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(KEYINPUT18), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n538), .B(new_n523), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n541), .B(KEYINPUT13), .Z(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n537), .A2(new_n541), .A3(new_n539), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT18), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n542), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G113gat), .B(G141gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(G197gat), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT11), .B(G169gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT12), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n542), .A2(new_n556), .A3(new_n545), .A4(new_n548), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(KEYINPUT94), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n549), .A2(new_n559), .A3(new_n554), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n506), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(G64gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(G57gat), .ZN(new_n566));
  INV_X1    g365(.A(G57gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n567), .A2(G64gat), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT9), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  OR2_X1    g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT95), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(new_n565), .B2(G57gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT96), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(new_n567), .B2(G64gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n567), .A2(KEYINPUT95), .A3(G64gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n565), .A2(KEYINPUT96), .A3(G57gat), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n574), .A2(new_n576), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT9), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n570), .B1(new_n571), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n572), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT21), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G127gat), .B(G155gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G183gat), .B(G211gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT97), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n589), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n583), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n538), .B1(KEYINPUT21), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n594), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n597), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G85gat), .A2(G92gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  NAND2_X1  g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  INV_X1    g403(.A(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(KEYINPUT8), .A2(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G99gat), .B(G106gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  NAND2_X1  g409(.A1(new_n524), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  AND2_X1   g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n612), .A2(new_n523), .B1(KEYINPUT41), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G190gat), .B(G218gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n613), .A2(KEYINPUT41), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT100), .ZN(new_n619));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n617), .B(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT102), .B1(new_n600), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n597), .B(new_n598), .ZN(new_n624));
  INV_X1    g423(.A(new_n622), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT102), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n610), .A2(new_n629), .A3(new_n583), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n583), .B1(new_n632), .B2(new_n608), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n610), .B(new_n633), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n634), .A2(KEYINPUT104), .A3(new_n629), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT104), .B1(new_n634), .B2(new_n629), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n631), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(G230gat), .A2(G233gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n634), .A2(new_n639), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(G120gat), .B(G148gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT105), .ZN(new_n645));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n647), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n640), .A2(new_n642), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n648), .A2(KEYINPUT106), .A3(new_n650), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n628), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n564), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n480), .A2(KEYINPUT107), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n480), .A2(KEYINPUT107), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(new_n529), .ZN(G1324gat));
  INV_X1    g461(.A(new_n657), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n346), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n664), .A2(G8gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT108), .B(KEYINPUT16), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G8gat), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT42), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n669), .B1(KEYINPUT42), .B2(new_n668), .ZN(G1325gat));
  AOI21_X1  g469(.A(G15gat), .B1(new_n663), .B2(new_n310), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n504), .B(KEYINPUT109), .Z(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(G15gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT110), .Z(new_n675));
  AOI21_X1  g474(.A(new_n671), .B1(new_n675), .B2(new_n663), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n657), .A2(new_n455), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NAND4_X1  g478(.A1(new_n600), .A2(new_n654), .A3(new_n653), .A4(new_n622), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT111), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n563), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n684), .A2(G29gat), .A3(new_n660), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT45), .Z(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n478), .B1(new_n453), .B2(new_n454), .ZN(new_n688));
  AOI22_X1  g487(.A1(new_n688), .A2(new_n498), .B1(new_n500), .B2(new_n460), .ZN(new_n689));
  AOI22_X1  g488(.A1(new_n689), .A2(new_n504), .B1(new_n451), .B2(new_n462), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n687), .B1(new_n690), .B2(new_n625), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n506), .A2(KEYINPUT44), .A3(new_n622), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n660), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n655), .A2(new_n624), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT112), .B1(new_n695), .B2(new_n562), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT112), .ZN(new_n697));
  NOR4_X1   g496(.A1(new_n655), .A2(new_n561), .A3(new_n624), .A4(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n693), .A2(new_n694), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(G29gat), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n701), .ZN(G1328gat));
  NOR3_X1   g501(.A1(new_n684), .A2(G36gat), .A3(new_n458), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT46), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n693), .A2(new_n346), .A3(new_n699), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT113), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G36gat), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n705), .A2(KEYINPUT113), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(G1329gat));
  INV_X1    g508(.A(new_n504), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n710), .A3(new_n699), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G43gat), .ZN(new_n712));
  INV_X1    g511(.A(new_n310), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(G43gat), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n563), .A2(new_n682), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n712), .A2(KEYINPUT47), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n691), .A2(new_n673), .A3(new_n692), .A4(new_n699), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G43gat), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n717), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT114), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n716), .B1(new_n719), .B2(G43gat), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT114), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n724), .A2(new_n725), .A3(KEYINPUT47), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n718), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT115), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT115), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n718), .B(new_n729), .C1(new_n723), .C2(new_n726), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1330gat));
  NAND4_X1  g530(.A1(new_n693), .A2(G50gat), .A3(new_n500), .A4(new_n699), .ZN(new_n732));
  INV_X1    g531(.A(G50gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n684), .B2(new_n455), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT48), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n736), .A2(KEYINPUT116), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(KEYINPUT116), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT117), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n732), .A2(new_n734), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(KEYINPUT48), .ZN(new_n741));
  AOI211_X1 g540(.A(KEYINPUT117), .B(new_n735), .C1(new_n732), .C2(new_n734), .ZN(new_n742));
  OAI22_X1  g541(.A1(new_n737), .A2(new_n738), .B1(new_n741), .B2(new_n742), .ZN(G1331gat));
  INV_X1    g542(.A(new_n655), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n628), .A2(new_n562), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n506), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT118), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n660), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(new_n567), .ZN(G1332gat));
  AOI21_X1  g548(.A(new_n458), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  OR3_X1    g550(.A1(new_n747), .A2(KEYINPUT119), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT119), .B1(new_n747), .B2(new_n751), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n753), .B1(new_n752), .B2(new_n754), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(G1333gat));
  OAI21_X1  g556(.A(G71gat), .B1(new_n747), .B2(new_n672), .ZN(new_n758));
  INV_X1    g557(.A(G71gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n310), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n747), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1334gat));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n455), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g564(.A1(new_n744), .A2(new_n562), .A3(new_n624), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n693), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G85gat), .B1(new_n767), .B2(new_n660), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n690), .A2(new_n625), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n562), .A2(new_n624), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT51), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n769), .A2(new_n773), .A3(new_n770), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n655), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n694), .A2(new_n605), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n768), .B1(new_n775), .B2(new_n776), .ZN(G1336gat));
  OAI21_X1  g576(.A(G92gat), .B1(new_n767), .B2(new_n458), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n458), .A2(G92gat), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n772), .A2(new_n655), .A3(new_n774), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n780), .B2(KEYINPUT120), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n781), .B(new_n783), .ZN(G1337gat));
  XNOR2_X1  g583(.A(KEYINPUT121), .B(G99gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n767), .B2(new_n672), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n713), .A2(new_n785), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n775), .B2(new_n787), .ZN(G1338gat));
  NAND4_X1  g587(.A1(new_n772), .A2(new_n500), .A3(new_n655), .A4(new_n774), .ZN(new_n789));
  INV_X1    g588(.A(G106gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n693), .A2(G106gat), .A3(new_n500), .A4(new_n766), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT122), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(G1339gat));
  NOR2_X1   g594(.A1(new_n540), .A2(new_n541), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n543), .A2(new_n544), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n553), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n557), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT123), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n799), .B(new_n800), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n637), .A2(new_n639), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(KEYINPUT54), .A3(new_n640), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n640), .A2(KEYINPUT54), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(new_n647), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n801), .A2(new_n650), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n624), .B1(new_n809), .B2(new_n622), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n655), .A2(new_n557), .A3(new_n798), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n808), .A2(new_n650), .A3(new_n807), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n625), .B(new_n811), .C1(new_n812), .C2(new_n561), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n810), .A2(new_n813), .B1(new_n656), .B2(new_n561), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n814), .A2(new_n500), .A3(new_n713), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n660), .A2(new_n346), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n562), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n655), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(G120gat), .ZN(G1341gat));
  NAND3_X1  g620(.A1(new_n815), .A2(new_n624), .A3(new_n816), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT124), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT124), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n815), .A2(new_n824), .A3(new_n624), .A4(new_n816), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  XOR2_X1   g625(.A(KEYINPUT67), .B(G127gat), .Z(new_n827));
  XNOR2_X1  g626(.A(new_n826), .B(new_n827), .ZN(G1342gat));
  AND3_X1   g627(.A1(new_n815), .A2(new_n622), .A3(new_n816), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n829), .A2(KEYINPUT56), .A3(new_n211), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT56), .B1(new_n829), .B2(new_n211), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n830), .A2(new_n831), .B1(new_n211), .B2(new_n829), .ZN(G1343gat));
  NAND2_X1  g631(.A1(new_n810), .A2(new_n813), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n656), .A2(new_n561), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n455), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT57), .B1(new_n814), .B2(new_n455), .ZN(new_n838));
  INV_X1    g637(.A(new_n816), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n839), .A2(new_n710), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n561), .A2(new_n347), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n837), .A2(new_n838), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n673), .A2(new_n839), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n835), .A2(new_n562), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n347), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n846), .B(KEYINPUT58), .Z(G1344gat));
  AND2_X1   g646(.A1(new_n835), .A2(new_n843), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n349), .A3(new_n655), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n837), .A2(new_n838), .A3(new_n655), .A4(new_n840), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n850), .A2(new_n851), .A3(G148gat), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n850), .B2(G148gat), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n849), .B1(new_n852), .B2(new_n853), .ZN(G1345gat));
  NAND3_X1  g653(.A1(new_n848), .A2(new_n357), .A3(new_n624), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n837), .A2(new_n838), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n856), .A2(new_n624), .A3(new_n840), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n855), .B1(new_n857), .B2(new_n357), .ZN(G1346gat));
  NAND3_X1  g657(.A1(new_n848), .A2(new_n358), .A3(new_n622), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n856), .A2(new_n622), .A3(new_n840), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n859), .B1(new_n860), .B2(new_n358), .ZN(G1347gat));
  INV_X1    g660(.A(KEYINPUT125), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n694), .A2(new_n458), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n815), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n562), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n862), .B1(new_n866), .B2(G169gat), .ZN(new_n867));
  OR4_X1    g666(.A1(new_n862), .A2(new_n864), .A3(G169gat), .A4(new_n561), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(G169gat), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(G1348gat));
  NAND2_X1  g669(.A1(new_n865), .A2(new_n655), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(G176gat), .ZN(G1349gat));
  OAI21_X1  g671(.A(new_n217), .B1(new_n864), .B2(new_n600), .ZN(new_n873));
  NAND2_X1  g672(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n874));
  INV_X1    g673(.A(new_n235), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n815), .A2(new_n875), .A3(new_n624), .A4(new_n863), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n874), .B1(new_n873), .B2(new_n876), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(G1350gat));
  OAI22_X1  g678(.A1(new_n864), .A2(new_n625), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n880));
  NAND2_X1  g679(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n880), .B(new_n881), .ZN(G1351gat));
  AND2_X1   g681(.A1(new_n672), .A2(new_n863), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n837), .A2(new_n838), .A3(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(G197gat), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n884), .A2(new_n885), .A3(new_n561), .ZN(new_n886));
  NOR4_X1   g685(.A1(new_n814), .A2(new_n458), .A3(new_n455), .A4(new_n694), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n887), .A2(new_n672), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n562), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n886), .B1(new_n885), .B2(new_n889), .ZN(G1352gat));
  NOR2_X1   g689(.A1(new_n744), .A2(G204gat), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n887), .A2(new_n672), .A3(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G204gat), .B1(new_n884), .B2(new_n744), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n893), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(G1353gat));
  NAND3_X1  g696(.A1(new_n888), .A2(new_n317), .A3(new_n624), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n837), .A2(new_n838), .A3(new_n624), .A4(new_n883), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n899), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT63), .B1(new_n899), .B2(G211gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(G1354gat));
  AND2_X1   g701(.A1(new_n884), .A2(KEYINPUT127), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n622), .B1(new_n884), .B2(KEYINPUT127), .ZN(new_n904));
  OAI21_X1  g703(.A(G218gat), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n318), .A3(new_n622), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1355gat));
endmodule


