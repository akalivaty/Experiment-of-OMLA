

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U549 ( .A(n720), .ZN(n586) );
  XNOR2_X1 U550 ( .A(n649), .B(n648), .ZN(n655) );
  INV_X1 U551 ( .A(KEYINPUT29), .ZN(n648) );
  NOR2_X1 U552 ( .A1(n664), .A2(n663), .ZN(n666) );
  XNOR2_X1 U553 ( .A(n670), .B(KEYINPUT89), .ZN(n658) );
  INV_X1 U554 ( .A(KEYINPUT97), .ZN(n707) );
  XNOR2_X1 U555 ( .A(KEYINPUT66), .B(n518), .ZN(n519) );
  AND2_X1 U556 ( .A1(n528), .A2(n527), .ZN(G160) );
  OR2_X1 U557 ( .A1(n716), .A2(n715), .ZN(n516) );
  INV_X1 U558 ( .A(n656), .ZN(n651) );
  INV_X1 U559 ( .A(KEYINPUT28), .ZN(n644) );
  BUF_X1 U560 ( .A(n656), .Z(n672) );
  NAND2_X1 U561 ( .A1(n655), .A2(n654), .ZN(n668) );
  INV_X1 U562 ( .A(G1966), .ZN(n657) );
  AND2_X1 U563 ( .A1(n658), .A2(n657), .ZN(n685) );
  NAND2_X1 U564 ( .A1(n586), .A2(n721), .ZN(n656) );
  OR2_X1 U565 ( .A1(n610), .A2(n543), .ZN(n611) );
  NAND2_X1 U566 ( .A1(n717), .A2(n516), .ZN(n718) );
  OR2_X1 U567 ( .A1(n719), .A2(n718), .ZN(n723) );
  INV_X1 U568 ( .A(KEYINPUT72), .ZN(n621) );
  XNOR2_X1 U569 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X2 U570 ( .A1(G2104), .A2(n521), .ZN(n902) );
  AND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n900) );
  XNOR2_X1 U572 ( .A(n624), .B(n623), .ZN(n971) );
  OR2_X1 U573 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  XOR2_X2 U575 ( .A(KEYINPUT17), .B(n517), .Z(n907) );
  NAND2_X1 U576 ( .A1(G137), .A2(n907), .ZN(n520) );
  INV_X1 U577 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n900), .A2(G113), .ZN(n518) );
  AND2_X1 U579 ( .A1(n520), .A2(n519), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n902), .A2(G125), .ZN(n522) );
  XNOR2_X1 U581 ( .A(n522), .B(KEYINPUT64), .ZN(n525) );
  AND2_X2 U582 ( .A1(n521), .A2(G2104), .ZN(n906) );
  NAND2_X1 U583 ( .A1(n906), .A2(G101), .ZN(n523) );
  XOR2_X1 U584 ( .A(KEYINPUT23), .B(n523), .Z(n524) );
  NAND2_X1 U585 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U586 ( .A(n526), .B(KEYINPUT65), .ZN(n527) );
  NAND2_X1 U587 ( .A1(G102), .A2(n906), .ZN(n530) );
  NAND2_X1 U588 ( .A1(G138), .A2(n907), .ZN(n529) );
  NAND2_X1 U589 ( .A1(n530), .A2(n529), .ZN(n534) );
  NAND2_X1 U590 ( .A1(G126), .A2(n902), .ZN(n532) );
  NAND2_X1 U591 ( .A1(G114), .A2(n900), .ZN(n531) );
  NAND2_X1 U592 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U593 ( .A1(n534), .A2(n533), .ZN(G164) );
  NOR2_X1 U594 ( .A1(G651), .A2(G543), .ZN(n814) );
  NAND2_X1 U595 ( .A1(G90), .A2(n814), .ZN(n538) );
  INV_X1 U596 ( .A(G543), .ZN(n535) );
  NAND2_X1 U597 ( .A1(KEYINPUT0), .A2(n535), .ZN(n613) );
  INV_X1 U598 ( .A(KEYINPUT0), .ZN(n536) );
  NAND2_X1 U599 ( .A1(n536), .A2(G543), .ZN(n540) );
  NAND2_X1 U600 ( .A1(n613), .A2(n540), .ZN(n612) );
  INV_X1 U601 ( .A(G651), .ZN(n543) );
  NOR2_X1 U602 ( .A1(n612), .A2(n543), .ZN(n815) );
  NAND2_X1 U603 ( .A1(G77), .A2(n815), .ZN(n537) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n539), .B(KEYINPUT9), .ZN(n542) );
  AND2_X1 U606 ( .A1(n540), .A2(n543), .ZN(n615) );
  AND2_X1 U607 ( .A1(n613), .A2(n615), .ZN(n811) );
  NAND2_X1 U608 ( .A1(G52), .A2(n811), .ZN(n541) );
  NAND2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n547) );
  NOR2_X1 U610 ( .A1(G543), .A2(n543), .ZN(n544) );
  XOR2_X1 U611 ( .A(KEYINPUT1), .B(n544), .Z(n607) );
  BUF_X1 U612 ( .A(n607), .Z(n810) );
  NAND2_X1 U613 ( .A1(n810), .A2(G64), .ZN(n545) );
  XOR2_X1 U614 ( .A(KEYINPUT68), .B(n545), .Z(n546) );
  NOR2_X1 U615 ( .A1(n547), .A2(n546), .ZN(G171) );
  NAND2_X1 U616 ( .A1(n810), .A2(G63), .ZN(n548) );
  XOR2_X1 U617 ( .A(KEYINPUT73), .B(n548), .Z(n550) );
  NAND2_X1 U618 ( .A1(n811), .A2(G51), .ZN(n549) );
  NAND2_X1 U619 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U620 ( .A(KEYINPUT6), .B(n551), .ZN(n557) );
  NAND2_X1 U621 ( .A1(n814), .A2(G89), .ZN(n552) );
  XNOR2_X1 U622 ( .A(n552), .B(KEYINPUT4), .ZN(n554) );
  NAND2_X1 U623 ( .A1(G76), .A2(n815), .ZN(n553) );
  NAND2_X1 U624 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U625 ( .A(n555), .B(KEYINPUT5), .Z(n556) );
  NOR2_X1 U626 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U627 ( .A(KEYINPUT7), .B(n558), .Z(n559) );
  XNOR2_X1 U628 ( .A(KEYINPUT74), .B(n559), .ZN(G168) );
  XOR2_X1 U629 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U630 ( .A1(G88), .A2(n814), .ZN(n561) );
  NAND2_X1 U631 ( .A1(G75), .A2(n815), .ZN(n560) );
  NAND2_X1 U632 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U633 ( .A1(G62), .A2(n810), .ZN(n563) );
  NAND2_X1 U634 ( .A1(G50), .A2(n811), .ZN(n562) );
  NAND2_X1 U635 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U636 ( .A1(n565), .A2(n564), .ZN(G166) );
  NAND2_X1 U637 ( .A1(G87), .A2(n612), .ZN(n567) );
  NAND2_X1 U638 ( .A1(G74), .A2(G651), .ZN(n566) );
  NAND2_X1 U639 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U640 ( .A1(n810), .A2(n568), .ZN(n571) );
  NAND2_X1 U641 ( .A1(G49), .A2(n811), .ZN(n569) );
  XOR2_X1 U642 ( .A(KEYINPUT79), .B(n569), .Z(n570) );
  NAND2_X1 U643 ( .A1(n571), .A2(n570), .ZN(G288) );
  INV_X1 U644 ( .A(G166), .ZN(G303) );
  NAND2_X1 U645 ( .A1(G86), .A2(n814), .ZN(n573) );
  NAND2_X1 U646 ( .A1(G61), .A2(n810), .ZN(n572) );
  NAND2_X1 U647 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n815), .A2(G73), .ZN(n574) );
  XOR2_X1 U649 ( .A(KEYINPUT2), .B(n574), .Z(n575) );
  NOR2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n811), .A2(G48), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n578), .A2(n577), .ZN(G305) );
  NAND2_X1 U653 ( .A1(G85), .A2(n814), .ZN(n580) );
  NAND2_X1 U654 ( .A1(G72), .A2(n815), .ZN(n579) );
  NAND2_X1 U655 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U656 ( .A(KEYINPUT67), .B(n581), .ZN(n585) );
  NAND2_X1 U657 ( .A1(G60), .A2(n810), .ZN(n583) );
  NAND2_X1 U658 ( .A1(G47), .A2(n811), .ZN(n582) );
  AND2_X1 U659 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n585), .A2(n584), .ZN(G290) );
  NAND2_X1 U661 ( .A1(G160), .A2(G40), .ZN(n720) );
  NOR2_X1 U662 ( .A1(G164), .A2(G1384), .ZN(n721) );
  NAND2_X1 U663 ( .A1(n651), .A2(G2072), .ZN(n587) );
  XNOR2_X1 U664 ( .A(KEYINPUT27), .B(n587), .ZN(n590) );
  NAND2_X1 U665 ( .A1(G1956), .A2(n672), .ZN(n588) );
  XNOR2_X1 U666 ( .A(KEYINPUT91), .B(n588), .ZN(n589) );
  NOR2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n643) );
  NAND2_X1 U668 ( .A1(G91), .A2(n814), .ZN(n592) );
  NAND2_X1 U669 ( .A1(G78), .A2(n815), .ZN(n591) );
  NAND2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U671 ( .A1(G65), .A2(n810), .ZN(n594) );
  NAND2_X1 U672 ( .A1(G53), .A2(n811), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U674 ( .A1(n596), .A2(n595), .ZN(n955) );
  NAND2_X1 U675 ( .A1(n643), .A2(n955), .ZN(n642) );
  XNOR2_X1 U676 ( .A(KEYINPUT69), .B(KEYINPUT13), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n814), .A2(G81), .ZN(n597) );
  XNOR2_X1 U678 ( .A(n597), .B(KEYINPUT12), .ZN(n599) );
  NAND2_X1 U679 ( .A1(G68), .A2(n815), .ZN(n598) );
  NAND2_X1 U680 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U681 ( .A(n601), .B(n600), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n810), .A2(G56), .ZN(n602) );
  XOR2_X1 U683 ( .A(KEYINPUT14), .B(n602), .Z(n603) );
  NOR2_X1 U684 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n811), .A2(G43), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n606), .A2(n605), .ZN(n957) );
  NAND2_X1 U687 ( .A1(G92), .A2(n814), .ZN(n609) );
  NAND2_X1 U688 ( .A1(G66), .A2(n607), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(n620) );
  INV_X1 U690 ( .A(G79), .ZN(n610) );
  OR2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n617) );
  AND2_X1 U692 ( .A1(n613), .A2(G54), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U695 ( .A(n618), .B(KEYINPUT71), .Z(n619) );
  NOR2_X1 U696 ( .A1(n620), .A2(n619), .ZN(n624) );
  INV_X1 U697 ( .A(KEYINPUT15), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n971), .A2(G1348), .ZN(n625) );
  NAND2_X1 U699 ( .A1(n625), .A2(KEYINPUT26), .ZN(n626) );
  NOR2_X1 U700 ( .A1(G1341), .A2(n626), .ZN(n627) );
  NOR2_X1 U701 ( .A1(n627), .A2(n651), .ZN(n629) );
  NOR2_X1 U702 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n628) );
  NOR2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n634) );
  NAND2_X1 U704 ( .A1(KEYINPUT26), .A2(G1996), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n971), .A2(G2067), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n651), .A2(n632), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U709 ( .A1(n957), .A2(n635), .ZN(n640) );
  NAND2_X1 U710 ( .A1(G1348), .A2(n672), .ZN(n637) );
  NAND2_X1 U711 ( .A1(G2067), .A2(n651), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U713 ( .A1(n971), .A2(n638), .ZN(n639) );
  NOR2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U715 ( .A1(n642), .A2(n641), .ZN(n647) );
  NOR2_X1 U716 ( .A1(n643), .A2(n955), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n649) );
  NOR2_X1 U719 ( .A1(n651), .A2(G1961), .ZN(n650) );
  XOR2_X1 U720 ( .A(KEYINPUT90), .B(n650), .Z(n653) );
  XNOR2_X1 U721 ( .A(G2078), .B(KEYINPUT25), .ZN(n935) );
  NAND2_X1 U722 ( .A1(n651), .A2(n935), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n662) );
  NAND2_X1 U724 ( .A1(n662), .A2(G171), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n656), .A2(G8), .ZN(n670) );
  NOR2_X1 U726 ( .A1(G2084), .A2(n672), .ZN(n681) );
  NOR2_X1 U727 ( .A1(n685), .A2(n681), .ZN(n659) );
  NAND2_X1 U728 ( .A1(G8), .A2(n659), .ZN(n660) );
  XNOR2_X1 U729 ( .A(KEYINPUT30), .B(n660), .ZN(n661) );
  NOR2_X1 U730 ( .A1(n661), .A2(G168), .ZN(n664) );
  NOR2_X1 U731 ( .A1(G171), .A2(n662), .ZN(n663) );
  XOR2_X1 U732 ( .A(KEYINPUT31), .B(KEYINPUT92), .Z(n665) );
  XNOR2_X1 U733 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n683) );
  AND2_X1 U735 ( .A1(G286), .A2(G8), .ZN(n669) );
  NAND2_X1 U736 ( .A1(n683), .A2(n669), .ZN(n679) );
  INV_X1 U737 ( .A(G8), .ZN(n677) );
  XOR2_X1 U738 ( .A(KEYINPUT89), .B(n670), .Z(n716) );
  NOR2_X1 U739 ( .A1(G1971), .A2(n716), .ZN(n671) );
  XNOR2_X1 U740 ( .A(KEYINPUT93), .B(n671), .ZN(n675) );
  NOR2_X1 U741 ( .A1(G2090), .A2(n672), .ZN(n673) );
  NOR2_X1 U742 ( .A1(G166), .A2(n673), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n676) );
  OR2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U746 ( .A(n680), .B(KEYINPUT32), .ZN(n687) );
  NAND2_X1 U747 ( .A1(G8), .A2(n681), .ZN(n682) );
  NAND2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U749 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U750 ( .A1(n687), .A2(n686), .ZN(n689) );
  INV_X1 U751 ( .A(KEYINPUT94), .ZN(n688) );
  XNOR2_X1 U752 ( .A(n689), .B(n688), .ZN(n711) );
  NOR2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n693) );
  NOR2_X1 U754 ( .A1(G1971), .A2(G303), .ZN(n690) );
  NOR2_X1 U755 ( .A1(n693), .A2(n690), .ZN(n975) );
  NAND2_X1 U756 ( .A1(n711), .A2(n975), .ZN(n691) );
  NAND2_X1 U757 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NAND2_X1 U758 ( .A1(n691), .A2(n974), .ZN(n692) );
  XNOR2_X1 U759 ( .A(n692), .B(KEYINPUT95), .ZN(n700) );
  INV_X1 U760 ( .A(n716), .ZN(n696) );
  INV_X1 U761 ( .A(KEYINPUT33), .ZN(n702) );
  NAND2_X1 U762 ( .A1(n696), .A2(n693), .ZN(n694) );
  NOR2_X1 U763 ( .A1(n702), .A2(n694), .ZN(n695) );
  XOR2_X1 U764 ( .A(n695), .B(KEYINPUT96), .Z(n701) );
  AND2_X1 U765 ( .A1(n696), .A2(n701), .ZN(n698) );
  XNOR2_X1 U766 ( .A(G1981), .B(G305), .ZN(n967) );
  INV_X1 U767 ( .A(n967), .ZN(n697) );
  AND2_X1 U768 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U769 ( .A1(n700), .A2(n699), .ZN(n706) );
  INV_X1 U770 ( .A(n701), .ZN(n703) );
  OR2_X1 U771 ( .A1(n703), .A2(n702), .ZN(n704) );
  OR2_X1 U772 ( .A1(n967), .A2(n704), .ZN(n705) );
  NAND2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n708) );
  XNOR2_X1 U774 ( .A(n708), .B(n707), .ZN(n719) );
  NOR2_X1 U775 ( .A1(G2090), .A2(G303), .ZN(n709) );
  NAND2_X1 U776 ( .A1(G8), .A2(n709), .ZN(n710) );
  XNOR2_X1 U777 ( .A(n710), .B(KEYINPUT98), .ZN(n712) );
  NAND2_X1 U778 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U779 ( .A1(n713), .A2(n716), .ZN(n717) );
  NOR2_X1 U780 ( .A1(G1981), .A2(G305), .ZN(n714) );
  XOR2_X1 U781 ( .A(n714), .B(KEYINPUT24), .Z(n715) );
  NOR2_X1 U782 ( .A1(n721), .A2(n720), .ZN(n767) );
  XNOR2_X1 U783 ( .A(G1986), .B(G290), .ZN(n959) );
  NAND2_X1 U784 ( .A1(n767), .A2(n959), .ZN(n722) );
  NAND2_X1 U785 ( .A1(n723), .A2(n722), .ZN(n755) );
  XNOR2_X1 U786 ( .A(KEYINPUT37), .B(G2067), .ZN(n765) );
  NAND2_X1 U787 ( .A1(G104), .A2(n906), .ZN(n725) );
  NAND2_X1 U788 ( .A1(G140), .A2(n907), .ZN(n724) );
  NAND2_X1 U789 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U790 ( .A(KEYINPUT34), .B(n726), .ZN(n731) );
  NAND2_X1 U791 ( .A1(G128), .A2(n902), .ZN(n728) );
  NAND2_X1 U792 ( .A1(G116), .A2(n900), .ZN(n727) );
  NAND2_X1 U793 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U794 ( .A(KEYINPUT35), .B(n729), .Z(n730) );
  NOR2_X1 U795 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U796 ( .A(KEYINPUT36), .B(n732), .ZN(n920) );
  NOR2_X1 U797 ( .A1(n765), .A2(n920), .ZN(n1024) );
  NAND2_X1 U798 ( .A1(n1024), .A2(n767), .ZN(n764) );
  NAND2_X1 U799 ( .A1(G117), .A2(n900), .ZN(n733) );
  XNOR2_X1 U800 ( .A(n733), .B(KEYINPUT86), .ZN(n742) );
  NAND2_X1 U801 ( .A1(G105), .A2(n906), .ZN(n734) );
  XOR2_X1 U802 ( .A(KEYINPUT87), .B(n734), .Z(n735) );
  XNOR2_X1 U803 ( .A(n735), .B(KEYINPUT38), .ZN(n737) );
  NAND2_X1 U804 ( .A1(G129), .A2(n902), .ZN(n736) );
  NAND2_X1 U805 ( .A1(n737), .A2(n736), .ZN(n740) );
  NAND2_X1 U806 ( .A1(n907), .A2(G141), .ZN(n738) );
  XOR2_X1 U807 ( .A(KEYINPUT88), .B(n738), .Z(n739) );
  NOR2_X1 U808 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U809 ( .A1(n742), .A2(n741), .ZN(n915) );
  AND2_X1 U810 ( .A1(n915), .A2(G1996), .ZN(n751) );
  NAND2_X1 U811 ( .A1(n906), .A2(G95), .ZN(n745) );
  NAND2_X1 U812 ( .A1(G119), .A2(n902), .ZN(n743) );
  XOR2_X1 U813 ( .A(KEYINPUT85), .B(n743), .Z(n744) );
  NAND2_X1 U814 ( .A1(n745), .A2(n744), .ZN(n749) );
  NAND2_X1 U815 ( .A1(G107), .A2(n900), .ZN(n747) );
  NAND2_X1 U816 ( .A1(G131), .A2(n907), .ZN(n746) );
  NAND2_X1 U817 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U818 ( .A1(n749), .A2(n748), .ZN(n897) );
  INV_X1 U819 ( .A(G1991), .ZN(n938) );
  NOR2_X1 U820 ( .A1(n897), .A2(n938), .ZN(n750) );
  NOR2_X1 U821 ( .A1(n751), .A2(n750), .ZN(n1013) );
  INV_X1 U822 ( .A(n767), .ZN(n752) );
  NOR2_X1 U823 ( .A1(n1013), .A2(n752), .ZN(n758) );
  INV_X1 U824 ( .A(n758), .ZN(n753) );
  NAND2_X1 U825 ( .A1(n764), .A2(n753), .ZN(n754) );
  NOR2_X1 U826 ( .A1(n755), .A2(n754), .ZN(n771) );
  NOR2_X1 U827 ( .A1(G1996), .A2(n915), .ZN(n1017) );
  NOR2_X1 U828 ( .A1(G1986), .A2(G290), .ZN(n756) );
  AND2_X1 U829 ( .A1(n938), .A2(n897), .ZN(n1015) );
  NOR2_X1 U830 ( .A1(n756), .A2(n1015), .ZN(n757) );
  NOR2_X1 U831 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U832 ( .A(KEYINPUT99), .B(n759), .Z(n760) );
  NOR2_X1 U833 ( .A1(n1017), .A2(n760), .ZN(n761) );
  XOR2_X1 U834 ( .A(KEYINPUT39), .B(n761), .Z(n762) );
  XOR2_X1 U835 ( .A(KEYINPUT100), .B(n762), .Z(n763) );
  NAND2_X1 U836 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U837 ( .A1(n765), .A2(n920), .ZN(n1026) );
  NAND2_X1 U838 ( .A1(n766), .A2(n1026), .ZN(n768) );
  NAND2_X1 U839 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U840 ( .A(n769), .B(KEYINPUT101), .ZN(n770) );
  XNOR2_X1 U841 ( .A(n772), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U842 ( .A(G2451), .B(G2454), .Z(n774) );
  XNOR2_X1 U843 ( .A(G2430), .B(KEYINPUT102), .ZN(n773) );
  XNOR2_X1 U844 ( .A(n774), .B(n773), .ZN(n775) );
  XOR2_X1 U845 ( .A(n775), .B(G2446), .Z(n777) );
  XNOR2_X1 U846 ( .A(G1348), .B(G1341), .ZN(n776) );
  XNOR2_X1 U847 ( .A(n777), .B(n776), .ZN(n781) );
  XOR2_X1 U848 ( .A(G2438), .B(G2427), .Z(n779) );
  XNOR2_X1 U849 ( .A(G2443), .B(G2435), .ZN(n778) );
  XNOR2_X1 U850 ( .A(n779), .B(n778), .ZN(n780) );
  XOR2_X1 U851 ( .A(n781), .B(n780), .Z(n782) );
  AND2_X1 U852 ( .A1(G14), .A2(n782), .ZN(G401) );
  AND2_X1 U853 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U854 ( .A1(G123), .A2(n902), .ZN(n783) );
  XNOR2_X1 U855 ( .A(n783), .B(KEYINPUT18), .ZN(n791) );
  NAND2_X1 U856 ( .A1(n906), .A2(G99), .ZN(n784) );
  XNOR2_X1 U857 ( .A(n784), .B(KEYINPUT78), .ZN(n786) );
  NAND2_X1 U858 ( .A1(G135), .A2(n907), .ZN(n785) );
  NAND2_X1 U859 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U860 ( .A1(G111), .A2(n900), .ZN(n787) );
  XNOR2_X1 U861 ( .A(KEYINPUT77), .B(n787), .ZN(n788) );
  NOR2_X1 U862 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U863 ( .A1(n791), .A2(n790), .ZN(n1012) );
  XNOR2_X1 U864 ( .A(G2096), .B(n1012), .ZN(n792) );
  OR2_X1 U865 ( .A1(G2100), .A2(n792), .ZN(G156) );
  INV_X1 U866 ( .A(G132), .ZN(G219) );
  INV_X1 U867 ( .A(G82), .ZN(G220) );
  INV_X1 U868 ( .A(G96), .ZN(G221) );
  INV_X1 U869 ( .A(G57), .ZN(G237) );
  INV_X1 U870 ( .A(G120), .ZN(G236) );
  NAND2_X1 U871 ( .A1(G7), .A2(G661), .ZN(n793) );
  XNOR2_X1 U872 ( .A(n793), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U873 ( .A(G223), .ZN(n849) );
  NAND2_X1 U874 ( .A1(n849), .A2(G567), .ZN(n794) );
  XOR2_X1 U875 ( .A(KEYINPUT11), .B(n794), .Z(G234) );
  INV_X1 U876 ( .A(G860), .ZN(n802) );
  OR2_X1 U877 ( .A1(n957), .A2(n802), .ZN(G153) );
  XOR2_X1 U878 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  INV_X1 U879 ( .A(G868), .ZN(n795) );
  NOR2_X1 U880 ( .A1(G301), .A2(n795), .ZN(n797) );
  NOR2_X1 U881 ( .A1(n971), .A2(G868), .ZN(n796) );
  NOR2_X1 U882 ( .A1(n797), .A2(n796), .ZN(G284) );
  INV_X1 U883 ( .A(n955), .ZN(G299) );
  XNOR2_X1 U884 ( .A(KEYINPUT75), .B(G868), .ZN(n798) );
  NOR2_X1 U885 ( .A1(G286), .A2(n798), .ZN(n800) );
  NOR2_X1 U886 ( .A1(G868), .A2(G299), .ZN(n799) );
  NOR2_X1 U887 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U888 ( .A(KEYINPUT76), .B(n801), .ZN(G297) );
  NAND2_X1 U889 ( .A1(n802), .A2(G559), .ZN(n803) );
  INV_X1 U890 ( .A(n971), .ZN(n808) );
  NAND2_X1 U891 ( .A1(n803), .A2(n808), .ZN(n804) );
  XNOR2_X1 U892 ( .A(n804), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U893 ( .A1(G868), .A2(n957), .ZN(n807) );
  NAND2_X1 U894 ( .A1(n808), .A2(G868), .ZN(n805) );
  NOR2_X1 U895 ( .A1(G559), .A2(n805), .ZN(n806) );
  NOR2_X1 U896 ( .A1(n807), .A2(n806), .ZN(G282) );
  NAND2_X1 U897 ( .A1(n808), .A2(G559), .ZN(n809) );
  XNOR2_X1 U898 ( .A(n809), .B(n957), .ZN(n826) );
  NOR2_X1 U899 ( .A1(n826), .A2(G860), .ZN(n820) );
  NAND2_X1 U900 ( .A1(G67), .A2(n810), .ZN(n813) );
  NAND2_X1 U901 ( .A1(G55), .A2(n811), .ZN(n812) );
  NAND2_X1 U902 ( .A1(n813), .A2(n812), .ZN(n819) );
  NAND2_X1 U903 ( .A1(G93), .A2(n814), .ZN(n817) );
  NAND2_X1 U904 ( .A1(G80), .A2(n815), .ZN(n816) );
  NAND2_X1 U905 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U906 ( .A1(n819), .A2(n818), .ZN(n828) );
  XNOR2_X1 U907 ( .A(n820), .B(n828), .ZN(G145) );
  XNOR2_X1 U908 ( .A(G166), .B(KEYINPUT19), .ZN(n825) );
  XNOR2_X1 U909 ( .A(n955), .B(n828), .ZN(n823) );
  XNOR2_X1 U910 ( .A(G305), .B(G288), .ZN(n821) );
  XNOR2_X1 U911 ( .A(n821), .B(G290), .ZN(n822) );
  XNOR2_X1 U912 ( .A(n823), .B(n822), .ZN(n824) );
  XNOR2_X1 U913 ( .A(n825), .B(n824), .ZN(n922) );
  XNOR2_X1 U914 ( .A(n826), .B(n922), .ZN(n827) );
  NAND2_X1 U915 ( .A1(n827), .A2(G868), .ZN(n830) );
  OR2_X1 U916 ( .A1(n828), .A2(G868), .ZN(n829) );
  NAND2_X1 U917 ( .A1(n830), .A2(n829), .ZN(G295) );
  NAND2_X1 U918 ( .A1(G2084), .A2(G2078), .ZN(n831) );
  XOR2_X1 U919 ( .A(KEYINPUT20), .B(n831), .Z(n832) );
  NAND2_X1 U920 ( .A1(G2090), .A2(n832), .ZN(n833) );
  XNOR2_X1 U921 ( .A(KEYINPUT21), .B(n833), .ZN(n834) );
  NAND2_X1 U922 ( .A1(n834), .A2(G2072), .ZN(n835) );
  XNOR2_X1 U923 ( .A(KEYINPUT80), .B(n835), .ZN(G158) );
  XNOR2_X1 U924 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U925 ( .A1(G236), .A2(G237), .ZN(n836) );
  NAND2_X1 U926 ( .A1(G69), .A2(n836), .ZN(n837) );
  XNOR2_X1 U927 ( .A(KEYINPUT83), .B(n837), .ZN(n838) );
  NAND2_X1 U928 ( .A1(n838), .A2(G108), .ZN(n855) );
  NAND2_X1 U929 ( .A1(G567), .A2(n855), .ZN(n839) );
  XOR2_X1 U930 ( .A(KEYINPUT84), .B(n839), .Z(n846) );
  NOR2_X1 U931 ( .A1(G220), .A2(G219), .ZN(n840) );
  XOR2_X1 U932 ( .A(KEYINPUT22), .B(n840), .Z(n841) );
  NOR2_X1 U933 ( .A1(G218), .A2(n841), .ZN(n842) );
  XNOR2_X1 U934 ( .A(n842), .B(KEYINPUT81), .ZN(n843) );
  NOR2_X1 U935 ( .A1(G221), .A2(n843), .ZN(n844) );
  XOR2_X1 U936 ( .A(KEYINPUT82), .B(n844), .Z(n854) );
  AND2_X1 U937 ( .A1(n854), .A2(G2106), .ZN(n845) );
  NOR2_X1 U938 ( .A1(n846), .A2(n845), .ZN(G319) );
  INV_X1 U939 ( .A(G319), .ZN(n848) );
  NAND2_X1 U940 ( .A1(G661), .A2(G483), .ZN(n847) );
  NOR2_X1 U941 ( .A1(n848), .A2(n847), .ZN(n851) );
  NAND2_X1 U942 ( .A1(n851), .A2(G36), .ZN(G176) );
  NAND2_X1 U943 ( .A1(G2106), .A2(n849), .ZN(G217) );
  AND2_X1 U944 ( .A1(G15), .A2(G2), .ZN(n850) );
  NAND2_X1 U945 ( .A1(G661), .A2(n850), .ZN(G259) );
  NAND2_X1 U946 ( .A1(G3), .A2(G1), .ZN(n852) );
  NAND2_X1 U947 ( .A1(n852), .A2(n851), .ZN(n853) );
  XOR2_X1 U948 ( .A(KEYINPUT103), .B(n853), .Z(G188) );
  INV_X1 U950 ( .A(G108), .ZN(G238) );
  NOR2_X1 U951 ( .A1(n855), .A2(n854), .ZN(G325) );
  INV_X1 U952 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U953 ( .A(G1961), .B(KEYINPUT41), .ZN(n865) );
  XOR2_X1 U954 ( .A(G1986), .B(G1976), .Z(n857) );
  XNOR2_X1 U955 ( .A(G1971), .B(G1981), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U957 ( .A(G1956), .B(G1966), .Z(n859) );
  XNOR2_X1 U958 ( .A(G1996), .B(G1991), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U960 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U961 ( .A(KEYINPUT106), .B(G2474), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(G229) );
  XOR2_X1 U964 ( .A(KEYINPUT105), .B(G2678), .Z(n867) );
  XNOR2_X1 U965 ( .A(KEYINPUT104), .B(KEYINPUT43), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U967 ( .A(KEYINPUT42), .B(G2090), .Z(n869) );
  XNOR2_X1 U968 ( .A(G2067), .B(G2072), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U970 ( .A(n871), .B(n870), .Z(n873) );
  XNOR2_X1 U971 ( .A(G2096), .B(G2100), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(n875) );
  XOR2_X1 U973 ( .A(G2084), .B(G2078), .Z(n874) );
  XNOR2_X1 U974 ( .A(n875), .B(n874), .ZN(G227) );
  NAND2_X1 U975 ( .A1(G100), .A2(n906), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n876), .B(KEYINPUT108), .ZN(n880) );
  XOR2_X1 U977 ( .A(KEYINPUT107), .B(KEYINPUT44), .Z(n878) );
  NAND2_X1 U978 ( .A1(G124), .A2(n902), .ZN(n877) );
  XNOR2_X1 U979 ( .A(n878), .B(n877), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G112), .A2(n900), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G136), .A2(n907), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U984 ( .A1(n884), .A2(n883), .ZN(G162) );
  NAND2_X1 U985 ( .A1(G103), .A2(n906), .ZN(n886) );
  NAND2_X1 U986 ( .A1(G139), .A2(n907), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n892) );
  NAND2_X1 U988 ( .A1(n902), .A2(G127), .ZN(n887) );
  XOR2_X1 U989 ( .A(KEYINPUT111), .B(n887), .Z(n889) );
  NAND2_X1 U990 ( .A1(n900), .A2(G115), .ZN(n888) );
  NAND2_X1 U991 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n890), .Z(n891) );
  NOR2_X1 U993 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U994 ( .A(KEYINPUT112), .B(n893), .Z(n1028) );
  XOR2_X1 U995 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n895) );
  XNOR2_X1 U996 ( .A(G164), .B(KEYINPUT113), .ZN(n894) );
  XNOR2_X1 U997 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n1012), .B(n896), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n897), .B(G162), .ZN(n898) );
  XNOR2_X1 U1000 ( .A(n899), .B(n898), .ZN(n914) );
  NAND2_X1 U1001 ( .A1(G118), .A2(n900), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n901), .B(KEYINPUT110), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(G130), .A2(n902), .ZN(n903) );
  XOR2_X1 U1004 ( .A(KEYINPUT109), .B(n903), .Z(n904) );
  NAND2_X1 U1005 ( .A1(n905), .A2(n904), .ZN(n912) );
  NAND2_X1 U1006 ( .A1(G106), .A2(n906), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(G142), .A2(n907), .ZN(n908) );
  NAND2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1009 ( .A(KEYINPUT45), .B(n910), .Z(n911) );
  NOR2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1011 ( .A(n914), .B(n913), .Z(n917) );
  XOR2_X1 U1012 ( .A(G160), .B(n915), .Z(n916) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1014 ( .A(n1028), .B(n918), .Z(n919) );
  XNOR2_X1 U1015 ( .A(n920), .B(n919), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n921), .ZN(G395) );
  XNOR2_X1 U1017 ( .A(n971), .B(G286), .ZN(n923) );
  XNOR2_X1 U1018 ( .A(n923), .B(n922), .ZN(n925) );
  XNOR2_X1 U1019 ( .A(n957), .B(G171), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(n925), .B(n924), .ZN(n926) );
  NOR2_X1 U1021 ( .A1(G37), .A2(n926), .ZN(G397) );
  NOR2_X1 U1022 ( .A1(G229), .A2(G227), .ZN(n927) );
  XOR2_X1 U1023 ( .A(KEYINPUT114), .B(n927), .Z(n928) );
  XNOR2_X1 U1024 ( .A(KEYINPUT49), .B(n928), .ZN(n933) );
  NOR2_X1 U1025 ( .A1(G395), .A2(G397), .ZN(n929) );
  XOR2_X1 U1026 ( .A(KEYINPUT115), .B(n929), .Z(n930) );
  NAND2_X1 U1027 ( .A1(G319), .A2(n930), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(G401), .A2(n931), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(G225) );
  INV_X1 U1030 ( .A(G225), .ZN(G308) );
  INV_X1 U1031 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1032 ( .A(G2084), .B(G34), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(n934), .B(KEYINPUT54), .ZN(n952) );
  XOR2_X1 U1034 ( .A(G27), .B(n935), .Z(n945) );
  XNOR2_X1 U1035 ( .A(G1996), .B(G32), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(G33), .B(G2072), .ZN(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(G25), .B(n938), .ZN(n939) );
  NAND2_X1 U1039 ( .A1(n939), .A2(G28), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(G26), .B(G2067), .ZN(n940) );
  NOR2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(KEYINPUT53), .B(KEYINPUT118), .ZN(n946) );
  XNOR2_X1 U1045 ( .A(n947), .B(n946), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(G35), .B(G2090), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(n950), .B(KEYINPUT119), .ZN(n951) );
  NOR2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1050 ( .A(KEYINPUT55), .B(n953), .Z(n954) );
  NOR2_X1 U1051 ( .A1(G29), .A2(n954), .ZN(n1009) );
  XNOR2_X1 U1052 ( .A(G16), .B(KEYINPUT56), .ZN(n982) );
  XNOR2_X1 U1053 ( .A(G1956), .B(n955), .ZN(n956) );
  XNOR2_X1 U1054 ( .A(n956), .B(KEYINPUT122), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(G1341), .B(n957), .ZN(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(G1961), .B(G171), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(KEYINPUT121), .B(n962), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n970) );
  XOR2_X1 U1061 ( .A(G1966), .B(KEYINPUT120), .Z(n965) );
  XNOR2_X1 U1062 ( .A(G168), .B(n965), .ZN(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1064 ( .A(KEYINPUT57), .B(n968), .Z(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(G1348), .B(n971), .ZN(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n980) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n977) );
  AND2_X1 U1069 ( .A1(G303), .A2(G1971), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1071 ( .A(KEYINPUT123), .B(n978), .Z(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n1007) );
  INV_X1 U1074 ( .A(G16), .ZN(n1005) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G21), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(G1961), .B(G5), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n995) );
  XNOR2_X1 U1078 ( .A(G1956), .B(G20), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(G19), .B(G1341), .ZN(n985) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n992) );
  XOR2_X1 U1081 ( .A(KEYINPUT124), .B(G4), .Z(n988) );
  XNOR2_X1 U1082 ( .A(G1348), .B(KEYINPUT59), .ZN(n987) );
  XNOR2_X1 U1083 ( .A(n988), .B(n987), .ZN(n990) );
  XNOR2_X1 U1084 ( .A(G1981), .B(G6), .ZN(n989) );
  NOR2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1087 ( .A(KEYINPUT60), .B(n993), .Z(n994) );
  NAND2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(G1971), .B(G22), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(G23), .B(G1976), .ZN(n996) );
  NOR2_X1 U1091 ( .A1(n997), .A2(n996), .ZN(n999) );
  XOR2_X1 U1092 ( .A(G1986), .B(G24), .Z(n998) );
  NAND2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1094 ( .A(KEYINPUT58), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1096 ( .A(KEYINPUT61), .B(n1003), .ZN(n1004) );
  NAND2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(G11), .A2(n1010), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(n1011), .B(KEYINPUT125), .ZN(n1040) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1022) );
  XOR2_X1 U1104 ( .A(G160), .B(G2084), .Z(n1020) );
  XOR2_X1 U1105 ( .A(G2090), .B(G162), .Z(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(KEYINPUT51), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1111 ( .A(n1025), .B(KEYINPUT116), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1034) );
  XOR2_X1 U1113 ( .A(G2072), .B(n1028), .Z(n1030) );
  XNOR2_X1 U1114 ( .A(G164), .B(G2078), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(KEYINPUT50), .B(n1031), .Z(n1032) );
  XNOR2_X1 U1117 ( .A(KEYINPUT117), .B(n1032), .ZN(n1033) );
  NOR2_X1 U1118 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1119 ( .A(KEYINPUT52), .B(n1035), .ZN(n1037) );
  INV_X1 U1120 ( .A(KEYINPUT55), .ZN(n1036) );
  NAND2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1122 ( .A1(n1038), .A2(G29), .ZN(n1039) );
  NAND2_X1 U1123 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1124 ( .A(KEYINPUT62), .B(n1041), .Z(G311) );
  XOR2_X1 U1125 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
endmodule

