//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  OR2_X1    g046(.A1(G100), .A2(G2105), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n472), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G124), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n477), .B1(G136), .B2(new_n463), .ZN(G162));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  OAI211_X1 g055(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n464), .B1(KEYINPUT67), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G114), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n483), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n480), .B1(new_n482), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n483), .ZN(new_n490));
  OAI21_X1  g065(.A(G2105), .B1(new_n486), .B2(G114), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n484), .A2(KEYINPUT67), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(KEYINPUT68), .A3(new_n481), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n474), .A2(G138), .A3(new_n464), .A4(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n464), .C1(new_n460), .C2(new_n461), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT69), .B(KEYINPUT4), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n479), .B1(new_n495), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n493), .A2(KEYINPUT68), .A3(new_n481), .ZN(new_n504));
  AOI21_X1  g079(.A(KEYINPUT68), .B1(new_n493), .B2(new_n481), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n479), .B(new_n502), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT71), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(new_n514), .A3(G651), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(new_n515), .B1(KEYINPUT6), .B2(new_n511), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n519), .A2(new_n521), .B1(new_n518), .B2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n516), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G50), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n510), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n511), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n526), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT74), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n516), .A2(new_n522), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT75), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n533), .A2(new_n535), .A3(KEYINPUT75), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n519), .A2(new_n521), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n518), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT73), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n522), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n547), .A2(G63), .A3(G651), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n516), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G51), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n538), .A2(new_n539), .A3(new_n548), .A4(new_n550), .ZN(G286));
  INV_X1    g126(.A(G286), .ZN(G168));
  AOI22_X1  g127(.A1(new_n547), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n511), .ZN(new_n554));
  AOI22_X1  g129(.A1(G52), .A2(new_n549), .B1(new_n534), .B2(G90), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT76), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n554), .A2(new_n556), .ZN(G171));
  INV_X1    g132(.A(G81), .ZN(new_n558));
  INV_X1    g133(.A(G43), .ZN(new_n559));
  OAI22_X1  g134(.A1(new_n558), .A2(new_n523), .B1(new_n524), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G68), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G56), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n546), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n560), .B1(new_n563), .B2(G651), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G860), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n566), .A2(new_n567), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(new_n549), .A2(G53), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n542), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(new_n534), .B2(G91), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(G299));
  NAND2_X1  g154(.A1(new_n554), .A2(new_n556), .ZN(G301));
  OAI21_X1  g155(.A(G651), .B1(new_n547), .B2(G74), .ZN(new_n581));
  AOI22_X1  g156(.A1(G49), .A2(new_n549), .B1(new_n534), .B2(G87), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(new_n534), .A2(G86), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(KEYINPUT78), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n522), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(new_n511), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n549), .A2(G48), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(KEYINPUT78), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n585), .A2(new_n587), .A3(new_n588), .A4(new_n589), .ZN(G305));
  AND3_X1   g165(.A1(new_n543), .A2(G60), .A3(new_n545), .ZN(new_n591));
  AND2_X1   g166(.A1(G72), .A2(G543), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(G47), .A2(new_n549), .B1(new_n534), .B2(G85), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n593), .A2(new_n594), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n602));
  OR3_X1    g177(.A1(new_n523), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n523), .B2(new_n601), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n522), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G54), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n606), .A2(new_n511), .B1(new_n607), .B2(new_n524), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G171), .B2(new_n610), .ZN(G284));
  XNOR2_X1  g187(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NAND2_X1  g188(.A1(G299), .A2(new_n610), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G168), .B2(new_n610), .ZN(G297));
  XNOR2_X1  g190(.A(G297), .B(KEYINPUT82), .ZN(G280));
  INV_X1    g191(.A(new_n609), .ZN(new_n617));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n566), .A2(new_n610), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n609), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n610), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT83), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g199(.A(new_n475), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G123), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n463), .A2(G135), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n464), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT84), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n474), .A2(new_n465), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2100), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n633), .A2(new_n634), .A3(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT85), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2427), .B(G2430), .Z(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n646), .B(new_n650), .Z(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  AND3_X1   g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT86), .Z(new_n658));
  NOR2_X1   g233(.A1(G2072), .A2(G2078), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n444), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n656), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n660), .B(KEYINPUT17), .Z(new_n663));
  OAI21_X1  g238(.A(new_n662), .B1(new_n663), .B2(new_n658), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n657), .A3(new_n656), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT18), .Z(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(new_n658), .A3(new_n656), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT87), .ZN(new_n669));
  XOR2_X1   g244(.A(G2096), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT20), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n673), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n673), .B2(new_n679), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT88), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n691), .A2(G6), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G305), .B2(G16), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT32), .B(G1981), .Z(new_n694));
  AND2_X1   g269(.A1(new_n691), .A2(G23), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G288), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT33), .B(G1976), .ZN(new_n697));
  AOI22_X1  g272(.A1(new_n693), .A2(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n696), .B2(new_n697), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n691), .A2(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n691), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G1971), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n693), .A2(new_n694), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n699), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT34), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n599), .A2(G16), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G16), .B2(G24), .ZN(new_n707));
  INV_X1    g282(.A(G1986), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n625), .A2(G119), .B1(new_n463), .B2(G131), .ZN(new_n710));
  OAI21_X1  g285(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g287(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n713));
  OAI221_X1 g288(.A(G2104), .B1(G107), .B2(new_n464), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G25), .B(new_n715), .S(G29), .Z(new_n716));
  XOR2_X1   g291(.A(KEYINPUT35), .B(G1991), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT90), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n707), .A2(new_n708), .ZN(new_n720));
  NOR4_X1   g295(.A1(new_n705), .A2(new_n709), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT36), .Z(new_n722));
  NOR2_X1   g297(.A1(G5), .A2(G16), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT95), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G301), .B2(new_n691), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT96), .Z(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(G1961), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n691), .A2(G19), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n566), .B2(G16), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n730), .A2(G1341), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(G1341), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n727), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(G164), .A2(G29), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G27), .B2(G29), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT97), .B(G2078), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n691), .A2(G21), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G168), .B2(new_n691), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n735), .A2(new_n736), .B1(new_n738), .B2(G1966), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G1966), .B2(new_n738), .ZN(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(G162), .A2(G29), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G29), .B2(G35), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT29), .B(G2090), .Z(new_n744));
  OAI22_X1  g319(.A1(new_n632), .A2(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G34), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(G29), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G160), .B2(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G2084), .ZN(new_n750));
  NOR2_X1   g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  AND2_X1   g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n753), .A2(G28), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n741), .B1(new_n753), .B2(G28), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n750), .B1(new_n751), .B2(new_n752), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n741), .A2(G32), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n463), .A2(G141), .B1(G105), .B2(new_n465), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n625), .A2(G129), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT26), .Z(new_n761));
  NAND3_X1  g336(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n757), .B1(new_n762), .B2(G29), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT27), .B(G1996), .ZN(new_n764));
  OAI22_X1  g339(.A1(new_n749), .A2(G2084), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR3_X1   g340(.A1(new_n745), .A2(new_n756), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n691), .A2(G4), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n617), .B2(new_n691), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(G1348), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(G1348), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n766), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n735), .A2(new_n736), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n741), .A2(G26), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n463), .A2(G140), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT91), .Z(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n778));
  INV_X1    g353(.A(G116), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(G2105), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n625), .B2(G128), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n775), .B1(new_n782), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2067), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n763), .A2(new_n764), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT94), .Z(new_n786));
  AND2_X1   g361(.A1(new_n741), .A2(G33), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n474), .A2(G127), .ZN(new_n788));
  AND2_X1   g363(.A1(G115), .A2(G2104), .ZN(new_n789));
  OAI21_X1  g364(.A(G2105), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT25), .ZN(new_n791));
  NAND2_X1  g366(.A1(G103), .A2(G2104), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(G2105), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n463), .A2(G139), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n787), .B1(new_n796), .B2(G29), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(new_n442), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n743), .A2(new_n744), .B1(new_n442), .B2(new_n797), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n784), .A2(new_n786), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NOR4_X1   g375(.A1(new_n740), .A2(new_n771), .A3(new_n772), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n691), .A2(G20), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT23), .Z(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G299), .B2(G16), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT98), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1956), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G1961), .B2(new_n726), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n722), .A2(new_n733), .A3(new_n801), .A4(new_n807), .ZN(G150));
  INV_X1    g383(.A(G150), .ZN(G311));
  AOI22_X1  g384(.A1(new_n547), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n511), .ZN(new_n811));
  INV_X1    g386(.A(G93), .ZN(new_n812));
  INV_X1    g387(.A(G55), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n812), .A2(new_n523), .B1(new_n524), .B2(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n566), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n811), .A2(new_n814), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(new_n564), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n617), .A2(G559), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(KEYINPUT39), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(KEYINPUT39), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n823), .A2(new_n567), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n817), .A2(new_n567), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(G145));
  NAND2_X1  g403(.A1(new_n625), .A2(G130), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n463), .A2(G142), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n464), .A2(G118), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n829), .B(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(new_n636), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n715), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n482), .A2(new_n488), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n502), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n835), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n782), .B(new_n796), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(new_n762), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n838), .B(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n631), .B(G160), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G162), .ZN(new_n843));
  AOI21_X1  g418(.A(G37), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n843), .B2(new_n841), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(G395));
  NAND2_X1  g422(.A1(new_n816), .A2(new_n818), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n621), .ZN(new_n849));
  XOR2_X1   g424(.A(G299), .B(new_n609), .Z(new_n850));
  INV_X1    g425(.A(KEYINPUT41), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n850), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n854), .B2(new_n849), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n855), .A2(KEYINPUT100), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(KEYINPUT100), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n599), .A2(G305), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n599), .A2(G305), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(G288), .B(G303), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n858), .A2(new_n861), .A3(new_n859), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT42), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n856), .A2(new_n857), .A3(new_n866), .ZN(new_n867));
  OR3_X1    g442(.A1(new_n866), .A2(new_n855), .A3(KEYINPUT100), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n868), .A3(G868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT101), .B1(new_n815), .B2(new_n610), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n871), .B1(new_n869), .B2(new_n872), .ZN(G295));
  AOI21_X1  g448(.A(new_n871), .B1(new_n869), .B2(new_n872), .ZN(G331));
  NAND2_X1  g449(.A1(G301), .A2(G286), .ZN(new_n875));
  NAND2_X1  g450(.A1(G171), .A2(G168), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n819), .A2(KEYINPUT102), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n876), .A2(new_n816), .A3(new_n818), .A4(new_n875), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(new_n875), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n848), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n883), .A2(new_n884), .A3(new_n852), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n883), .B2(new_n852), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n882), .A2(new_n850), .A3(new_n878), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n865), .B(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n877), .A2(new_n880), .A3(new_n850), .A4(new_n882), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n882), .A2(new_n878), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n852), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n865), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT43), .B1(new_n891), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n892), .A2(new_n900), .A3(new_n894), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n900), .B1(new_n892), .B2(new_n894), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n901), .A2(new_n890), .A3(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n903), .A2(new_n898), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n899), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT43), .B1(new_n903), .B2(new_n898), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n908));
  AOI21_X1  g483(.A(G37), .B1(new_n895), .B2(new_n865), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n908), .B(new_n909), .C1(new_n888), .C2(new_n890), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n906), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI211_X1 g488(.A(KEYINPUT106), .B(KEYINPUT44), .C1(new_n907), .C2(new_n910), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n905), .B1(new_n913), .B2(new_n914), .ZN(G397));
  XNOR2_X1  g490(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n916));
  AOI21_X1  g491(.A(G1384), .B1(new_n502), .B2(new_n836), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(KEYINPUT107), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(KEYINPUT107), .B2(new_n917), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n466), .A2(new_n470), .A3(G40), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n782), .A2(G2067), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n782), .A2(G2067), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n762), .B(G1996), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n715), .B(new_n717), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n599), .B(new_n708), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n922), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n932), .B(KEYINPUT109), .Z(new_n933));
  INV_X1    g508(.A(KEYINPUT120), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT119), .ZN(new_n935));
  NAND2_X1  g510(.A1(G286), .A2(G8), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT118), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n920), .B1(new_n917), .B2(KEYINPUT45), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT70), .ZN(new_n940));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  INV_X1    g516(.A(new_n916), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n940), .A2(new_n941), .A3(new_n506), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n938), .B1(new_n943), .B2(KEYINPUT114), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT114), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n508), .A2(new_n945), .A3(new_n941), .A4(new_n942), .ZN(new_n946));
  AOI21_X1  g521(.A(G1966), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n940), .A2(new_n941), .A3(new_n506), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n948), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT50), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n950), .B1(new_n917), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n952), .B1(new_n948), .B2(KEYINPUT50), .ZN(new_n953));
  INV_X1    g528(.A(new_n920), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n949), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G2084), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n947), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G8), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n935), .B(new_n937), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G1966), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n943), .A2(KEYINPUT114), .ZN(new_n961));
  INV_X1    g536(.A(new_n938), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n943), .A2(KEYINPUT114), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n948), .A2(KEYINPUT50), .ZN(new_n966));
  INV_X1    g541(.A(new_n952), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n948), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n968), .A2(new_n956), .A3(new_n920), .A4(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n958), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n936), .B(KEYINPUT118), .Z(new_n972));
  OAI21_X1  g547(.A(KEYINPUT119), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n959), .A2(new_n973), .A3(KEYINPUT51), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT119), .B(new_n975), .C1(new_n971), .C2(new_n972), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n957), .A2(new_n937), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n934), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT62), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n959), .A2(new_n973), .A3(KEYINPUT51), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n981), .A2(KEYINPUT120), .A3(new_n977), .A4(new_n976), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT123), .ZN(new_n984));
  NAND2_X1  g559(.A1(G303), .A2(G8), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT55), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n917), .A2(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n920), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n948), .B2(new_n916), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n990), .A2(G1971), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n954), .B1(new_n966), .B2(new_n967), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n969), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n996), .A2(G2090), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n993), .B(new_n994), .C1(new_n997), .C2(KEYINPUT112), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n997), .A2(KEYINPUT112), .ZN(new_n999));
  OAI211_X1 g574(.A(G8), .B(new_n987), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n920), .A2(new_n917), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G8), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1976), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(G288), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n581), .A2(G1976), .A3(new_n582), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1003), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n1007), .B(new_n1010), .Z(new_n1011));
  NAND3_X1  g586(.A1(new_n587), .A2(new_n588), .A3(new_n584), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(G1981), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(G305), .B2(G1981), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1002), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1011), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n917), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n954), .B1(KEYINPUT50), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(KEYINPUT50), .B2(new_n948), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n991), .B1(G2090), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n987), .B1(new_n1023), .B2(G8), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT53), .B1(new_n990), .B2(new_n443), .ZN(new_n1026));
  INV_X1    g601(.A(G1961), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1026), .B1(new_n996), .B2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n944), .A2(new_n946), .A3(KEYINPUT53), .A4(new_n443), .ZN(new_n1029));
  AOI21_X1  g604(.A(G301), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1000), .A2(new_n1025), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n983), .A2(new_n984), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n979), .A2(new_n982), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT62), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n984), .B1(new_n983), .B2(new_n1031), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g612(.A(G1976), .B(G288), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G305), .A2(G1981), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1003), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n1000), .B2(new_n1019), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n998), .B2(new_n999), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n986), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n957), .A2(new_n958), .A3(G286), .ZN(new_n1044));
  AND4_X1   g619(.A1(KEYINPUT63), .A2(new_n1044), .A3(new_n1018), .A4(new_n1011), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1000), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1041), .B1(new_n1046), .B2(KEYINPUT63), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1961), .B1(new_n995), .B2(new_n969), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n920), .B2(KEYINPUT121), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1051), .B(new_n988), .C1(KEYINPUT121), .C2(new_n920), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(new_n919), .ZN(new_n1053));
  NOR4_X1   g628(.A1(new_n1049), .A2(G171), .A3(new_n1026), .A4(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1048), .B1(new_n1030), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT122), .B(new_n1048), .C1(new_n1030), .C2(new_n1054), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1028), .A2(G301), .A3(new_n1029), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1049), .A2(new_n1026), .A3(new_n1053), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1059), .B(KEYINPUT54), .C1(G301), .C2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1057), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G1996), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT58), .B(G1341), .Z(new_n1064));
  AOI22_X1  g639(.A1(new_n990), .A2(new_n1063), .B1(new_n1001), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n1066));
  OR3_X1    g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n566), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n1065), .B2(new_n566), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1001), .A2(G2067), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n955), .B2(G1348), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n617), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1067), .B(new_n1068), .C1(new_n1071), .C2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1348), .B1(new_n995), .B2(new_n969), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n617), .B1(new_n1075), .B2(new_n1069), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n609), .B(new_n1070), .C1(new_n955), .C2(G1348), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1072), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1956), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1022), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n574), .A2(new_n1082), .A3(new_n578), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n574), .B2(new_n578), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT56), .B(G2072), .Z(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT115), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n990), .A2(new_n1087), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1081), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1085), .B1(new_n1081), .B2(new_n1088), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT117), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT61), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(KEYINPUT117), .B(KEYINPUT61), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1089), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1076), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1071), .A2(KEYINPUT116), .A3(new_n617), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1090), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1079), .A2(new_n1095), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1062), .A2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1103), .A2(new_n1033), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1000), .A2(new_n1025), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1047), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n933), .B1(new_n1037), .B2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n928), .A2(new_n714), .A3(new_n710), .A4(new_n717), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n921), .B1(new_n1108), .B2(new_n923), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n930), .A2(new_n922), .ZN(new_n1110));
  XOR2_X1   g685(.A(new_n1110), .B(KEYINPUT125), .Z(new_n1111));
  NOR3_X1   g686(.A1(G290), .A2(G1986), .A3(new_n921), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(KEYINPUT48), .B2(new_n1112), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1112), .A2(KEYINPUT48), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1109), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n922), .A2(new_n1063), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT46), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n922), .B1(new_n926), .B2(new_n762), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT124), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT47), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1115), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1107), .A2(new_n1124), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g700(.A(G319), .ZN(new_n1127));
  OR2_X1    g701(.A1(G227), .A2(new_n1127), .ZN(new_n1128));
  OR2_X1    g702(.A1(new_n1128), .A2(KEYINPUT126), .ZN(new_n1129));
  AOI21_X1  g703(.A(G401), .B1(new_n1128), .B2(KEYINPUT126), .ZN(new_n1130));
  AND4_X1   g704(.A1(new_n689), .A2(new_n845), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  AND3_X1   g705(.A1(new_n911), .A2(KEYINPUT127), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g706(.A(KEYINPUT127), .B1(new_n911), .B2(new_n1131), .ZN(new_n1133));
  NOR2_X1   g707(.A1(new_n1132), .A2(new_n1133), .ZN(G308));
  NAND2_X1  g708(.A1(new_n911), .A2(new_n1131), .ZN(G225));
endmodule


