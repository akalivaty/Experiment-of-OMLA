//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n580, new_n581, new_n582, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n594, new_n595, new_n596,
    new_n597, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT65), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT67), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT68), .Z(new_n452));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n452), .A2(G567), .B1(new_n455), .B2(G2106), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT69), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G125), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT70), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT70), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n461), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT71), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2105), .C1(new_n471), .C2(new_n473), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AND3_X1   g053(.A1(KEYINPUT72), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT3), .B1(KEYINPUT72), .B2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n465), .A2(G2105), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n482), .A2(G137), .B1(G101), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  NAND2_X1  g061(.A1(new_n482), .A2(G136), .ZN(new_n487));
  OAI21_X1  g062(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n487), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n492), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  OAI22_X1  g073(.A1(new_n488), .A2(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n492), .B1(new_n479), .B2(new_n480), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT4), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR3_X1   g077(.A1(new_n501), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT70), .ZN(new_n504));
  AOI21_X1  g079(.A(KEYINPUT70), .B1(new_n468), .B2(new_n469), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n499), .B1(new_n502), .B2(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT73), .B(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n508), .A2(KEYINPUT73), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT74), .A3(G651), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n512), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n510), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(KEYINPUT75), .B1(new_n510), .B2(KEYINPUT5), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G62), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n524), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n516), .A2(new_n521), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT5), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n536), .B2(G543), .ZN(new_n537));
  AOI211_X1 g112(.A(new_n525), .B(new_n509), .C1(new_n537), .C2(new_n527), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n534), .A2(G88), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n523), .A2(new_n533), .A3(new_n539), .ZN(G303));
  INV_X1    g115(.A(G303), .ZN(G166));
  NAND3_X1  g116(.A1(new_n534), .A2(G89), .A3(new_n538), .ZN(new_n542));
  AOI21_X1  g117(.A(KEYINPUT74), .B1(new_n520), .B2(G651), .ZN(new_n543));
  AOI211_X1 g118(.A(new_n513), .B(new_n515), .C1(new_n517), .C2(new_n519), .ZN(new_n544));
  OAI211_X1 g119(.A(G51), .B(new_n511), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n525), .B1(new_n537), .B2(new_n527), .ZN(new_n546));
  AND2_X1   g121(.A1(G63), .A2(G651), .ZN(new_n547));
  NAND3_X1  g122(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(KEYINPUT7), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(KEYINPUT7), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n546), .A2(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n542), .A2(new_n545), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(G168));
  NAND3_X1  g128(.A1(new_n534), .A2(G90), .A3(new_n538), .ZN(new_n554));
  OAI211_X1 g129(.A(G64), .B(new_n526), .C1(new_n528), .C2(new_n529), .ZN(new_n555));
  NAND2_X1  g130(.A1(G77), .A2(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  OAI211_X1 g133(.A(G52), .B(new_n511), .C1(new_n543), .C2(new_n544), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n554), .A2(new_n558), .A3(new_n559), .ZN(G171));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n561));
  OAI211_X1 g136(.A(G56), .B(new_n526), .C1(new_n528), .C2(new_n529), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  AND3_X1   g138(.A1(new_n562), .A2(KEYINPUT76), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(KEYINPUT76), .B1(new_n562), .B2(new_n563), .ZN(new_n565));
  NOR3_X1   g140(.A1(new_n564), .A2(new_n565), .A3(new_n515), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n522), .A2(G43), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n534), .A2(G81), .A3(new_n538), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n561), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n562), .A2(new_n563), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT76), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n562), .A2(KEYINPUT76), .A3(new_n563), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n573), .A2(new_n574), .A3(G651), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n575), .A2(KEYINPUT77), .A3(new_n567), .A4(new_n568), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G860), .ZN(G153));
  NAND4_X1  g153(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g154(.A1(G1), .A2(G3), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT8), .ZN(new_n581));
  NAND4_X1  g156(.A1(G319), .A2(G483), .A3(G661), .A4(new_n581), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT78), .ZN(G188));
  INV_X1    g158(.A(KEYINPUT9), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n534), .A2(new_n511), .ZN(new_n585));
  NAND2_X1  g160(.A1(KEYINPUT79), .A2(G53), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n522), .A2(KEYINPUT79), .A3(KEYINPUT9), .A4(G53), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n534), .A2(G91), .A3(new_n538), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n546), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n515), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n591), .ZN(G299));
  NAND3_X1  g167(.A1(new_n554), .A2(new_n558), .A3(new_n559), .ZN(G301));
  NAND2_X1  g168(.A1(new_n552), .A2(KEYINPUT80), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n542), .A2(new_n545), .A3(new_n595), .A4(new_n551), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G286));
  NAND2_X1  g173(.A1(new_n522), .A2(G49), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n546), .B2(G74), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n509), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n546), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n516), .B2(new_n521), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G87), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(G288));
  AOI22_X1  g181(.A1(new_n546), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(new_n515), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT81), .B1(new_n607), .B2(new_n515), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n604), .A2(G86), .B1(G48), .B2(new_n522), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(G305));
  NAND2_X1  g189(.A1(new_n522), .A2(G47), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n546), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G85), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n534), .A2(new_n538), .ZN(new_n618));
  OAI221_X1 g193(.A(new_n615), .B1(new_n515), .B2(new_n616), .C1(new_n617), .C2(new_n618), .ZN(G290));
  NAND2_X1  g194(.A1(G301), .A2(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n530), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(G54), .A2(new_n522), .B1(new_n623), .B2(G651), .ZN(new_n624));
  AOI21_X1  g199(.A(KEYINPUT10), .B1(new_n604), .B2(G92), .ZN(new_n625));
  AND4_X1   g200(.A1(KEYINPUT10), .A2(new_n534), .A3(G92), .A4(new_n538), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n620), .B1(new_n628), .B2(G868), .ZN(G284));
  OAI21_X1  g204(.A(new_n620), .B1(new_n628), .B2(G868), .ZN(G321));
  NOR2_X1   g205(.A1(G299), .A2(G868), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n597), .B2(G868), .ZN(G297));
  AOI21_X1  g207(.A(new_n631), .B1(new_n597), .B2(G868), .ZN(G280));
  XOR2_X1   g208(.A(KEYINPUT82), .B(G559), .Z(new_n634));
  OAI21_X1  g209(.A(new_n628), .B1(G860), .B2(new_n634), .ZN(G148));
  NAND2_X1  g210(.A1(new_n628), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n577), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n467), .A2(new_n470), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(new_n483), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  INV_X1    g218(.A(G2100), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n482), .A2(G135), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n489), .A2(G123), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n492), .A2(G111), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n647), .B(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n645), .A2(new_n646), .A3(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT85), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2430), .Z(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT84), .B(KEYINPUT14), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2451), .B(G2454), .Z(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(new_n668), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(G14), .A3(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G401));
  XNOR2_X1  g247(.A(G2072), .B(G2078), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT17), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(new_n675), .B2(new_n673), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT86), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n678), .A2(new_n675), .A3(new_n673), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT18), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(new_n675), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n674), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G2096), .B(G2100), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT19), .Z(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1961), .B(G1966), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT87), .ZN(new_n694));
  XOR2_X1   g269(.A(G1956), .B(G2474), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT88), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n692), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n697), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n696), .A2(new_n692), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n694), .A2(new_n695), .ZN(new_n703));
  MUX2_X1   g278(.A(new_n702), .B(new_n692), .S(new_n703), .Z(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n701), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n705), .B1(new_n701), .B2(new_n704), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(G1991), .B(G1996), .Z(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n710), .B1(new_n707), .B2(new_n708), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1981), .B(G1986), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n712), .A2(new_n715), .A3(new_n713), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(G229));
  NOR2_X1   g294(.A1(G27), .A2(G29), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G164), .B2(G29), .ZN(new_n721));
  INV_X1    g296(.A(G2078), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT30), .B(G28), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  OR2_X1    g300(.A1(KEYINPUT31), .A2(G11), .ZN(new_n726));
  NAND2_X1  g301(.A1(KEYINPUT31), .A2(G11), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n724), .A2(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n651), .B2(new_n725), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n482), .A2(G141), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n489), .A2(G129), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT26), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n734), .A2(new_n735), .B1(G105), .B2(new_n483), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n730), .A2(new_n731), .A3(new_n736), .ZN(new_n737));
  MUX2_X1   g312(.A(G32), .B(new_n737), .S(G29), .Z(new_n738));
  XOR2_X1   g313(.A(KEYINPUT27), .B(G1996), .Z(new_n739));
  AOI21_X1  g314(.A(new_n729), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n723), .B(new_n740), .C1(new_n738), .C2(new_n739), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT24), .ZN(new_n742));
  INV_X1    g317(.A(G34), .ZN(new_n743));
  AOI21_X1  g318(.A(G29), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n742), .B2(new_n743), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G160), .B2(new_n725), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n741), .B1(G2084), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n725), .A2(G26), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT28), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n489), .A2(G128), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT93), .Z(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n752));
  INV_X1    g327(.A(G116), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G2105), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n482), .B2(G140), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n749), .B1(new_n756), .B2(G29), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2067), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n725), .A2(G35), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT95), .Z(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n494), .B2(G29), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT29), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G2090), .ZN(new_n763));
  INV_X1    g338(.A(G16), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n764), .ZN(new_n766));
  INV_X1    g341(.A(G1966), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n747), .A2(new_n758), .A3(new_n763), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n764), .A2(G20), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT23), .ZN(new_n771));
  INV_X1    g346(.A(G299), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(new_n764), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1956), .ZN(new_n774));
  NOR2_X1   g349(.A1(G5), .A2(G16), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT94), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G301), .B2(new_n764), .ZN(new_n777));
  INV_X1    g352(.A(G1961), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n492), .A2(G103), .A3(G2104), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT25), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n482), .A2(G139), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n640), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n492), .ZN(new_n786));
  MUX2_X1   g361(.A(G33), .B(new_n786), .S(G29), .Z(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(G2072), .Z(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G2090), .B2(new_n762), .ZN(new_n789));
  OR4_X1    g364(.A1(new_n769), .A2(new_n774), .A3(new_n779), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n764), .A2(G19), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n577), .B2(new_n764), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G1341), .Z(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n628), .A2(new_n764), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G4), .B2(new_n764), .ZN(new_n796));
  INV_X1    g371(.A(G1348), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n798), .B(new_n799), .C1(G2084), .C2(new_n746), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n790), .A2(new_n794), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n725), .A2(G25), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n482), .A2(G131), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n489), .A2(G119), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n492), .A2(G107), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n804), .B(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT90), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n803), .B1(new_n809), .B2(new_n725), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT91), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT35), .B(G1991), .Z(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n811), .A2(new_n813), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n764), .A2(G24), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G290), .B2(G16), .ZN(new_n817));
  INV_X1    g392(.A(G1986), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n814), .A2(new_n815), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n764), .A2(G6), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n522), .A2(G48), .ZN(new_n823));
  INV_X1    g398(.A(G86), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n618), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n611), .B2(new_n610), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n822), .B1(new_n826), .B2(new_n764), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT92), .Z(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT32), .B(G1981), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n764), .A2(G23), .ZN(new_n832));
  INV_X1    g407(.A(G288), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n764), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT33), .B(G1976), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n764), .A2(G22), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G166), .B2(new_n764), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G1971), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n830), .A2(new_n831), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n821), .B1(new_n841), .B2(KEYINPUT34), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT34), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n830), .A2(new_n843), .A3(new_n831), .A4(new_n840), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT36), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT36), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n842), .A2(new_n847), .A3(new_n844), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n802), .B1(new_n846), .B2(new_n848), .ZN(G311));
  NAND2_X1  g424(.A1(new_n846), .A2(new_n848), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n801), .ZN(G150));
  NAND2_X1  g426(.A1(new_n522), .A2(G55), .ZN(new_n852));
  NAND2_X1  g427(.A1(G80), .A2(G543), .ZN(new_n853));
  INV_X1    g428(.A(G67), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n530), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G651), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n534), .A2(G93), .A3(new_n538), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n852), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(KEYINPUT97), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n852), .A2(new_n856), .A3(new_n860), .A4(new_n857), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G860), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT37), .Z(new_n864));
  OAI211_X1 g439(.A(new_n859), .B(new_n861), .C1(new_n566), .C2(new_n569), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n570), .A2(new_n576), .A3(new_n858), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n628), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT39), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT98), .Z(new_n873));
  INV_X1    g448(.A(G860), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n871), .B2(KEYINPUT39), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n864), .B1(new_n873), .B2(new_n875), .ZN(G145));
  XNOR2_X1  g451(.A(new_n485), .B(new_n651), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G162), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n756), .B(G164), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n879), .A2(new_n737), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n737), .ZN(new_n881));
  OR3_X1    g456(.A1(new_n880), .A2(new_n881), .A3(new_n786), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n786), .B1(new_n880), .B2(new_n881), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT100), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  OR3_X1    g464(.A1(new_n492), .A2(KEYINPUT99), .A3(G118), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT99), .B1(new_n492), .B2(G118), .ZN(new_n891));
  AND4_X1   g466(.A1(new_n888), .A2(new_n889), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n489), .A2(G130), .ZN(new_n893));
  AOI211_X1 g468(.A(new_n892), .B(new_n893), .C1(G142), .C2(new_n482), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n642), .ZN(new_n895));
  INV_X1    g470(.A(new_n809), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n885), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n897), .A2(new_n885), .A3(new_n898), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n878), .B1(new_n884), .B2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n882), .A2(new_n900), .A3(new_n883), .A4(new_n901), .ZN(new_n904));
  AOI21_X1  g479(.A(G37), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n884), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n902), .A2(new_n906), .A3(new_n882), .A4(new_n883), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n878), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g487(.A(G868), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n862), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n867), .B(new_n636), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n588), .A2(new_n591), .A3(new_n589), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT10), .ZN(new_n917));
  INV_X1    g492(.A(G92), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n917), .B1(new_n618), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n604), .A2(KEYINPUT10), .A3(G92), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n916), .A2(new_n921), .A3(new_n587), .A4(new_n624), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n627), .A2(G299), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT41), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT41), .B1(new_n922), .B2(new_n923), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n915), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n627), .A2(G299), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n627), .A2(G299), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n928), .B(new_n929), .C1(new_n933), .C2(new_n915), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n915), .A2(KEYINPUT104), .A3(new_n927), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n934), .B2(new_n935), .ZN(new_n938));
  XNOR2_X1  g513(.A(G305), .B(G303), .ZN(new_n939));
  OR2_X1    g514(.A1(G288), .A2(G290), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n941));
  NAND2_X1  g516(.A1(G288), .A2(G290), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n941), .B1(new_n940), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n939), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n944), .A2(new_n939), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT42), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n937), .B1(new_n938), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n947), .B(KEYINPUT42), .Z(new_n950));
  NAND4_X1  g525(.A1(new_n950), .A2(new_n936), .A3(new_n934), .A4(new_n935), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n914), .B1(new_n952), .B2(new_n913), .ZN(G295));
  OAI21_X1  g528(.A(new_n914), .B1(new_n952), .B2(new_n913), .ZN(G331));
  XOR2_X1   g529(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n594), .A2(G171), .A3(new_n596), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(G171), .B2(new_n552), .ZN(new_n959));
  NAND3_X1  g534(.A1(G168), .A2(KEYINPUT108), .A3(G301), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n957), .A2(KEYINPUT109), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n594), .A2(G171), .A3(new_n596), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n961), .A2(new_n964), .B1(new_n866), .B2(new_n865), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n959), .A2(new_n960), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n594), .A2(KEYINPUT109), .A3(G171), .A4(new_n596), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(new_n867), .ZN(new_n969));
  OAI211_X1 g544(.A(KEYINPUT110), .B(new_n927), .C1(new_n965), .C2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n961), .A2(new_n866), .A3(new_n865), .A4(new_n964), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n867), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n932), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(new_n972), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT110), .B1(new_n975), .B2(new_n927), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(G37), .B1(new_n977), .B2(new_n947), .ZN(new_n978));
  INV_X1    g553(.A(new_n947), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n974), .B2(new_n976), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n956), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT41), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n930), .B2(new_n931), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n924), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n971), .B2(new_n972), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n973), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AOI211_X1 g562(.A(KEYINPUT111), .B(new_n984), .C1(new_n971), .C2(new_n972), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n979), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n975), .A2(new_n927), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n992), .A2(new_n947), .A3(new_n973), .A4(new_n970), .ZN(new_n993));
  INV_X1    g568(.A(G37), .ZN(new_n994));
  AND4_X1   g569(.A1(new_n956), .A2(new_n989), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n955), .B1(new_n981), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n989), .A2(new_n993), .A3(new_n994), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n978), .A2(new_n956), .A3(new_n980), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(new_n999), .A3(KEYINPUT44), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(new_n1000), .ZN(G397));
  XNOR2_X1  g576(.A(KEYINPUT113), .B(G40), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n484), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n475), .B2(new_n477), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT112), .B(G1384), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n506), .A2(new_n502), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(new_n499), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1004), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  OR3_X1    g585(.A1(new_n1010), .A2(G1986), .A3(G290), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n756), .A2(G2067), .ZN(new_n1013));
  INV_X1    g588(.A(G2067), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n751), .A2(new_n1014), .A3(new_n755), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1996), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n737), .B(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n896), .A2(new_n813), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n809), .A2(new_n812), .ZN(new_n1020));
  AND4_X1   g595(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  OAI22_X1  g596(.A1(new_n1011), .A2(new_n1012), .B1(new_n1021), .B2(new_n1010), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1009), .A2(new_n1017), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT46), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1016), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1009), .B1(new_n1026), .B2(new_n737), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1028), .B(KEYINPUT47), .Z(new_n1029));
  NAND2_X1  g604(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1015), .B1(new_n1030), .B2(new_n1020), .ZN(new_n1031));
  AOI211_X1 g606(.A(new_n1023), .B(new_n1029), .C1(new_n1009), .C2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1005), .B1(G164), .B2(G1384), .ZN(new_n1033));
  OAI211_X1 g608(.A(KEYINPUT45), .B(new_n1006), .C1(new_n1007), .C2(new_n499), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1004), .A2(new_n722), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1384), .ZN(new_n1038));
  OAI211_X1 g613(.A(KEYINPUT45), .B(new_n1038), .C1(new_n1007), .C2(new_n499), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1036), .A2(G2078), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1004), .A2(new_n1033), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1042), .B(new_n1038), .C1(new_n1007), .C2(new_n499), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1004), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n778), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1037), .A2(new_n1041), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(G171), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1008), .A2(new_n1005), .ZN(new_n1049));
  AND4_X1   g624(.A1(G40), .A2(new_n474), .A3(new_n484), .A4(new_n1040), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1034), .A3(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1037), .A2(new_n1051), .A3(new_n1046), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1048), .B1(G171), .B2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT126), .B(KEYINPUT54), .Z(new_n1054));
  OR2_X1    g629(.A1(new_n1047), .A2(G171), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(new_n1052), .B2(G171), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1053), .A2(new_n1054), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1981), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n612), .A2(new_n1059), .A3(new_n613), .ZN(new_n1060));
  OAI21_X1  g635(.A(G1981), .B1(new_n825), .B2(new_n608), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT49), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1060), .A2(KEYINPUT49), .A3(new_n1061), .ZN(new_n1065));
  INV_X1    g640(.A(G8), .ZN(new_n1066));
  NOR2_X1   g641(.A1(G164), .A2(G1384), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1066), .B1(new_n1004), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1064), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n601), .A2(G1976), .A3(new_n605), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n601), .A2(KEYINPUT117), .A3(G1976), .A4(new_n605), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1068), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT52), .ZN(new_n1075));
  INV_X1    g650(.A(G1976), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT52), .B1(G288), .B2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1077), .A2(new_n1068), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1069), .A2(new_n1075), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1004), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1080));
  INV_X1    g655(.A(G1971), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(G2090), .B2(new_n1045), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n1084));
  AOI22_X1  g659(.A1(G50), .A2(new_n522), .B1(new_n532), .B2(G651), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1066), .B1(new_n1085), .B2(new_n539), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1084), .B1(new_n1086), .B2(KEYINPUT55), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT55), .ZN(new_n1088));
  OAI211_X1 g663(.A(KEYINPUT115), .B(new_n1088), .C1(G166), .C2(new_n1066), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n1086), .B2(KEYINPUT55), .ZN(new_n1091));
  AND4_X1   g666(.A1(new_n1090), .A2(G303), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1087), .B(new_n1089), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1083), .A2(new_n1093), .A3(G8), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1083), .A2(new_n1093), .A3(KEYINPUT116), .A4(G8), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1079), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1093), .ZN(new_n1099));
  AOI21_X1  g674(.A(G2090), .B1(new_n1045), .B2(KEYINPUT118), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1003), .ZN(new_n1101));
  AND4_X1   g676(.A1(new_n478), .A2(new_n1043), .A3(new_n1101), .A4(new_n1044), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1100), .A2(new_n1104), .B1(new_n1081), .B2(new_n1080), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n1106));
  OAI21_X1  g681(.A(G8), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1108), .A2(new_n1106), .A3(new_n1082), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1099), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G2084), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1004), .A2(new_n1033), .A3(new_n1039), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1102), .A2(new_n1111), .B1(new_n1112), .B2(new_n767), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(G168), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n767), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1004), .A2(new_n1111), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(G168), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(G8), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT51), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1066), .B1(new_n1113), .B2(G168), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT51), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1058), .A2(new_n1098), .A3(new_n1110), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1956), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1045), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT56), .B(G2072), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1004), .A2(new_n1033), .A3(new_n1034), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(KEYINPUT121), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(KEYINPUT121), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1133), .A2(KEYINPUT57), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(KEYINPUT57), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n916), .A2(new_n587), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(G299), .A2(new_n1133), .A3(KEYINPUT57), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1132), .A2(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1139), .A2(KEYINPUT123), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1139), .A2(KEYINPUT123), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT124), .B1(new_n1144), .B2(new_n1132), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1045), .A2(new_n797), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1004), .A2(new_n1014), .A3(new_n1067), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1147), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n628), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1145), .A2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1144), .A2(new_n1132), .A3(KEYINPUT124), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1141), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n628), .B2(KEYINPUT125), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1151), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1157), .B1(new_n1158), .B2(new_n1149), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n628), .A2(KEYINPUT125), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI221_X1 g736(.A(new_n1157), .B1(KEYINPUT125), .B2(new_n628), .C1(new_n1158), .C2(new_n1149), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1150), .A2(new_n1156), .A3(new_n1151), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1004), .A2(new_n1067), .ZN(new_n1165));
  XOR2_X1   g740(.A(KEYINPUT58), .B(G1341), .Z(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1004), .A2(new_n1017), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1169), .A2(new_n1170), .A3(new_n577), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1170), .B1(new_n1169), .B2(new_n577), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1174), .B1(new_n1132), .B2(new_n1140), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1173), .B1(new_n1175), .B2(new_n1141), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1132), .A2(new_n1174), .A3(new_n1140), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1164), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1124), .B1(new_n1155), .B2(new_n1178), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1079), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1069), .A2(new_n1076), .A3(new_n833), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1060), .ZN(new_n1183));
  AOI22_X1  g758(.A1(new_n1180), .A2(new_n1181), .B1(new_n1068), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n552), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1121), .B1(new_n1120), .B2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1118), .A2(KEYINPUT51), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT62), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1048), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1119), .A2(new_n1191), .A3(new_n1122), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1110), .A2(new_n1098), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1184), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NOR3_X1   g770(.A1(new_n1113), .A2(new_n1066), .A3(G286), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1110), .A2(new_n1098), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1196), .A2(KEYINPUT63), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1093), .B1(new_n1083), .B2(G8), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AOI22_X1  g776(.A1(new_n1197), .A2(new_n1198), .B1(new_n1098), .B2(new_n1201), .ZN(new_n1202));
  NOR3_X1   g777(.A1(new_n1179), .A2(new_n1195), .A3(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(G290), .B(new_n818), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1010), .B1(new_n1021), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1032), .B1(new_n1203), .B2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g781(.A1(new_n981), .A2(new_n995), .ZN(new_n1208));
  OR3_X1    g782(.A1(G401), .A2(G227), .A3(new_n459), .ZN(new_n1209));
  AOI21_X1  g783(.A(new_n1209), .B1(new_n717), .B2(new_n718), .ZN(new_n1210));
  NAND2_X1  g784(.A1(new_n911), .A2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g785(.A1(new_n1208), .A2(new_n1211), .ZN(G308));
  OAI211_X1 g786(.A(new_n911), .B(new_n1210), .C1(new_n981), .C2(new_n995), .ZN(G225));
endmodule


