

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599;

  XOR2_X1 U323 ( .A(n369), .B(n368), .Z(n291) );
  XOR2_X1 U324 ( .A(n387), .B(n386), .Z(n590) );
  XOR2_X1 U325 ( .A(KEYINPUT41), .B(n590), .Z(n546) );
  INV_X1 U326 ( .A(G190GAT), .ZN(n467) );
  XNOR2_X1 U327 ( .A(n467), .B(KEYINPUT58), .ZN(n468) );
  XNOR2_X1 U328 ( .A(n469), .B(n468), .ZN(G1351GAT) );
  XOR2_X1 U329 ( .A(KEYINPUT14), .B(G64GAT), .Z(n293) );
  XNOR2_X1 U330 ( .A(G22GAT), .B(G78GAT), .ZN(n292) );
  XNOR2_X1 U331 ( .A(n293), .B(n292), .ZN(n312) );
  XNOR2_X1 U332 ( .A(G8GAT), .B(G183GAT), .ZN(n294) );
  XNOR2_X1 U333 ( .A(n294), .B(KEYINPUT79), .ZN(n335) );
  INV_X1 U334 ( .A(KEYINPUT13), .ZN(n295) );
  NAND2_X1 U335 ( .A1(KEYINPUT71), .A2(n295), .ZN(n298) );
  INV_X1 U336 ( .A(KEYINPUT71), .ZN(n296) );
  NAND2_X1 U337 ( .A1(n296), .A2(KEYINPUT13), .ZN(n297) );
  NAND2_X1 U338 ( .A1(n298), .A2(n297), .ZN(n300) );
  XNOR2_X1 U339 ( .A(G71GAT), .B(G57GAT), .ZN(n299) );
  XNOR2_X1 U340 ( .A(n300), .B(n299), .ZN(n370) );
  XNOR2_X1 U341 ( .A(n335), .B(n370), .ZN(n310) );
  XOR2_X1 U342 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n302) );
  XNOR2_X1 U343 ( .A(KEYINPUT12), .B(KEYINPUT81), .ZN(n301) );
  XNOR2_X1 U344 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U345 ( .A(G155GAT), .B(G211GAT), .Z(n304) );
  XOR2_X1 U346 ( .A(G1GAT), .B(KEYINPUT70), .Z(n349) );
  XOR2_X1 U347 ( .A(G15GAT), .B(G127GAT), .Z(n453) );
  XNOR2_X1 U348 ( .A(n349), .B(n453), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U350 ( .A(n306), .B(n305), .Z(n308) );
  NAND2_X1 U351 ( .A1(G231GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U352 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U353 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U354 ( .A(n312), .B(n311), .Z(n594) );
  INV_X1 U355 ( .A(n594), .ZN(n567) );
  XOR2_X1 U356 ( .A(G141GAT), .B(G22GAT), .Z(n359) );
  XNOR2_X1 U357 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n313) );
  XNOR2_X1 U358 ( .A(n313), .B(KEYINPUT2), .ZN(n420) );
  XNOR2_X1 U359 ( .A(n359), .B(n420), .ZN(n314) );
  XOR2_X1 U360 ( .A(G148GAT), .B(G78GAT), .Z(n372) );
  XNOR2_X1 U361 ( .A(n314), .B(n372), .ZN(n320) );
  XOR2_X1 U362 ( .A(G162GAT), .B(KEYINPUT75), .Z(n316) );
  XNOR2_X1 U363 ( .A(G50GAT), .B(G218GAT), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n395) );
  XOR2_X1 U365 ( .A(n395), .B(KEYINPUT24), .Z(n318) );
  NAND2_X1 U366 ( .A1(G228GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U368 ( .A(n320), .B(n319), .Z(n328) );
  XOR2_X1 U369 ( .A(KEYINPUT90), .B(G211GAT), .Z(n322) );
  XNOR2_X1 U370 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U372 ( .A(G197GAT), .B(n323), .Z(n333) );
  XOR2_X1 U373 ( .A(KEYINPUT91), .B(KEYINPUT23), .Z(n325) );
  XNOR2_X1 U374 ( .A(G106GAT), .B(KEYINPUT22), .ZN(n324) );
  XNOR2_X1 U375 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U376 ( .A(n333), .B(n326), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n479) );
  XOR2_X1 U378 ( .A(KEYINPUT88), .B(KEYINPUT17), .Z(n330) );
  XNOR2_X1 U379 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n330), .B(n329), .ZN(n332) );
  XOR2_X1 U381 ( .A(KEYINPUT18), .B(KEYINPUT87), .Z(n331) );
  XOR2_X1 U382 ( .A(n332), .B(n331), .Z(n460) );
  INV_X1 U383 ( .A(n460), .ZN(n334) );
  XOR2_X1 U384 ( .A(n334), .B(n333), .Z(n343) );
  XOR2_X1 U385 ( .A(G176GAT), .B(G64GAT), .Z(n371) );
  XOR2_X1 U386 ( .A(n371), .B(n335), .Z(n337) );
  NAND2_X1 U387 ( .A1(G226GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U389 ( .A(n338), .B(KEYINPUT95), .Z(n341) );
  XNOR2_X1 U390 ( .A(G36GAT), .B(G190GAT), .ZN(n339) );
  XNOR2_X1 U391 ( .A(n339), .B(G92GAT), .ZN(n393) );
  XNOR2_X1 U392 ( .A(G218GAT), .B(n393), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U394 ( .A(n343), .B(n342), .ZN(n533) );
  XOR2_X1 U395 ( .A(KEYINPUT68), .B(KEYINPUT66), .Z(n345) );
  XNOR2_X1 U396 ( .A(G8GAT), .B(KEYINPUT30), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n345), .B(n344), .ZN(n363) );
  XOR2_X1 U398 ( .A(G113GAT), .B(G15GAT), .Z(n347) );
  XNOR2_X1 U399 ( .A(G50GAT), .B(G36GAT), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U401 ( .A(n348), .B(G197GAT), .Z(n351) );
  XNOR2_X1 U402 ( .A(G169GAT), .B(n349), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U404 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n353) );
  NAND2_X1 U405 ( .A1(G229GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U406 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U407 ( .A(n355), .B(n354), .Z(n361) );
  XOR2_X1 U408 ( .A(KEYINPUT69), .B(KEYINPUT7), .Z(n357) );
  XNOR2_X1 U409 ( .A(G43GAT), .B(G29GAT), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U411 ( .A(KEYINPUT8), .B(n358), .Z(n396) );
  XNOR2_X1 U412 ( .A(n396), .B(n359), .ZN(n360) );
  XNOR2_X1 U413 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n363), .B(n362), .ZN(n587) );
  INV_X1 U415 ( .A(G92GAT), .ZN(n364) );
  NAND2_X1 U416 ( .A1(KEYINPUT31), .A2(n364), .ZN(n367) );
  INV_X1 U417 ( .A(KEYINPUT31), .ZN(n365) );
  NAND2_X1 U418 ( .A1(n365), .A2(G92GAT), .ZN(n366) );
  NAND2_X1 U419 ( .A1(n367), .A2(n366), .ZN(n369) );
  XNOR2_X1 U420 ( .A(G120GAT), .B(G204GAT), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n291), .B(n370), .ZN(n374) );
  XNOR2_X1 U422 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U423 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U424 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n376) );
  NAND2_X1 U425 ( .A1(G230GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U426 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U427 ( .A(n378), .B(n377), .Z(n387) );
  INV_X1 U428 ( .A(KEYINPUT73), .ZN(n379) );
  NAND2_X1 U429 ( .A1(KEYINPUT72), .A2(n379), .ZN(n382) );
  INV_X1 U430 ( .A(KEYINPUT72), .ZN(n380) );
  NAND2_X1 U431 ( .A1(n380), .A2(KEYINPUT73), .ZN(n381) );
  NAND2_X1 U432 ( .A1(n382), .A2(n381), .ZN(n384) );
  XNOR2_X1 U433 ( .A(G106GAT), .B(G85GAT), .ZN(n383) );
  XNOR2_X1 U434 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U435 ( .A(G99GAT), .B(n385), .Z(n394) );
  XNOR2_X1 U436 ( .A(n394), .B(KEYINPUT33), .ZN(n386) );
  NAND2_X1 U437 ( .A1(n587), .A2(n546), .ZN(n388) );
  XNOR2_X1 U438 ( .A(n388), .B(KEYINPUT46), .ZN(n404) );
  XOR2_X1 U439 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n390) );
  XNOR2_X1 U440 ( .A(G134GAT), .B(KEYINPUT77), .ZN(n389) );
  XNOR2_X1 U441 ( .A(n390), .B(n389), .ZN(n392) );
  XOR2_X1 U442 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n391) );
  XNOR2_X1 U443 ( .A(n392), .B(n391), .ZN(n400) );
  XOR2_X1 U444 ( .A(n394), .B(n393), .Z(n398) );
  XNOR2_X1 U445 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U446 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U447 ( .A(n400), .B(n399), .ZN(n402) );
  NAND2_X1 U448 ( .A1(G232GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U449 ( .A(n402), .B(n401), .ZN(n571) );
  NOR2_X1 U450 ( .A1(n594), .A2(n571), .ZN(n403) );
  AND2_X1 U451 ( .A1(n404), .A2(n403), .ZN(n406) );
  XNOR2_X1 U452 ( .A(KEYINPUT47), .B(KEYINPUT113), .ZN(n405) );
  XNOR2_X1 U453 ( .A(n406), .B(n405), .ZN(n413) );
  XNOR2_X1 U454 ( .A(n571), .B(KEYINPUT78), .ZN(n466) );
  XNOR2_X1 U455 ( .A(KEYINPUT36), .B(KEYINPUT101), .ZN(n407) );
  XNOR2_X1 U456 ( .A(n466), .B(n407), .ZN(n496) );
  NOR2_X1 U457 ( .A1(n567), .A2(n496), .ZN(n409) );
  XNOR2_X1 U458 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n408) );
  XNOR2_X1 U459 ( .A(n409), .B(n408), .ZN(n411) );
  OR2_X1 U460 ( .A1(n590), .A2(n587), .ZN(n410) );
  NOR2_X1 U461 ( .A1(n411), .A2(n410), .ZN(n412) );
  NOR2_X1 U462 ( .A1(n413), .A2(n412), .ZN(n414) );
  XNOR2_X1 U463 ( .A(n414), .B(KEYINPUT48), .ZN(n558) );
  NOR2_X1 U464 ( .A1(n533), .A2(n558), .ZN(n415) );
  XNOR2_X1 U465 ( .A(n415), .B(KEYINPUT54), .ZN(n436) );
  XOR2_X1 U466 ( .A(G57GAT), .B(KEYINPUT1), .Z(n417) );
  XNOR2_X1 U467 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n416) );
  XNOR2_X1 U468 ( .A(n417), .B(n416), .ZN(n435) );
  XOR2_X1 U469 ( .A(G120GAT), .B(KEYINPUT0), .Z(n419) );
  XNOR2_X1 U470 ( .A(G113GAT), .B(G134GAT), .ZN(n418) );
  XNOR2_X1 U471 ( .A(n419), .B(n418), .ZN(n452) );
  XNOR2_X1 U472 ( .A(n452), .B(n420), .ZN(n433) );
  XOR2_X1 U473 ( .A(G85GAT), .B(G162GAT), .Z(n422) );
  XNOR2_X1 U474 ( .A(G29GAT), .B(G127GAT), .ZN(n421) );
  XNOR2_X1 U475 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U476 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n424) );
  XNOR2_X1 U477 ( .A(G141GAT), .B(G148GAT), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U479 ( .A(n426), .B(n425), .Z(n431) );
  XOR2_X1 U480 ( .A(KEYINPUT92), .B(KEYINPUT6), .Z(n428) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U483 ( .A(G1GAT), .B(n429), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U485 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U486 ( .A(n435), .B(n434), .Z(n477) );
  INV_X1 U487 ( .A(n477), .ZN(n530) );
  NAND2_X1 U488 ( .A1(n436), .A2(n530), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n437), .B(KEYINPUT64), .ZN(n585) );
  NOR2_X1 U490 ( .A1(n479), .A2(n585), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n438), .B(KEYINPUT122), .ZN(n440) );
  INV_X1 U492 ( .A(KEYINPUT55), .ZN(n439) );
  NAND2_X1 U493 ( .A1(n440), .A2(n439), .ZN(n443) );
  INV_X1 U494 ( .A(n440), .ZN(n441) );
  NAND2_X1 U495 ( .A1(KEYINPUT55), .A2(n441), .ZN(n442) );
  NAND2_X1 U496 ( .A1(n443), .A2(n442), .ZN(n462) );
  XOR2_X1 U497 ( .A(G176GAT), .B(G190GAT), .Z(n445) );
  XNOR2_X1 U498 ( .A(G43GAT), .B(G99GAT), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U500 ( .A(G71GAT), .B(G183GAT), .Z(n447) );
  XNOR2_X1 U501 ( .A(KEYINPUT89), .B(KEYINPUT86), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U503 ( .A(n449), .B(n448), .Z(n459) );
  XOR2_X1 U504 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n451) );
  XNOR2_X1 U505 ( .A(KEYINPUT20), .B(KEYINPUT85), .ZN(n450) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n457) );
  XOR2_X1 U507 ( .A(n453), .B(n452), .Z(n455) );
  NAND2_X1 U508 ( .A1(G227GAT), .A2(G233GAT), .ZN(n454) );
  XNOR2_X1 U509 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U511 ( .A(n459), .B(n458), .ZN(n461) );
  XOR2_X1 U512 ( .A(n461), .B(n460), .Z(n542) );
  NAND2_X1 U513 ( .A1(n462), .A2(n542), .ZN(n577) );
  NOR2_X1 U514 ( .A1(n567), .A2(n577), .ZN(n465) );
  INV_X1 U515 ( .A(G183GAT), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n463), .B(KEYINPUT124), .ZN(n464) );
  XNOR2_X1 U517 ( .A(n465), .B(n464), .ZN(G1350GAT) );
  INV_X1 U518 ( .A(n466), .ZN(n482) );
  NOR2_X1 U519 ( .A1(n482), .A2(n577), .ZN(n469) );
  INV_X1 U520 ( .A(n587), .ZN(n574) );
  NOR2_X1 U521 ( .A1(n574), .A2(n590), .ZN(n500) );
  INV_X1 U522 ( .A(n542), .ZN(n535) );
  NOR2_X1 U523 ( .A1(n533), .A2(n535), .ZN(n470) );
  NOR2_X1 U524 ( .A1(n479), .A2(n470), .ZN(n471) );
  XOR2_X1 U525 ( .A(n471), .B(KEYINPUT25), .Z(n472) );
  XNOR2_X1 U526 ( .A(KEYINPUT96), .B(n472), .ZN(n475) );
  NAND2_X1 U527 ( .A1(n535), .A2(n479), .ZN(n473) );
  XNOR2_X1 U528 ( .A(n473), .B(KEYINPUT26), .ZN(n584) );
  XNOR2_X1 U529 ( .A(n533), .B(KEYINPUT27), .ZN(n478) );
  NOR2_X1 U530 ( .A1(n584), .A2(n478), .ZN(n474) );
  NOR2_X1 U531 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U532 ( .A1(n477), .A2(n476), .ZN(n481) );
  NOR2_X1 U533 ( .A1(n530), .A2(n478), .ZN(n560) );
  XOR2_X1 U534 ( .A(n479), .B(KEYINPUT28), .Z(n538) );
  NAND2_X1 U535 ( .A1(n560), .A2(n538), .ZN(n541) );
  NOR2_X1 U536 ( .A1(n542), .A2(n541), .ZN(n480) );
  NOR2_X1 U537 ( .A1(n481), .A2(n480), .ZN(n497) );
  NAND2_X1 U538 ( .A1(n482), .A2(n594), .ZN(n483) );
  XNOR2_X1 U539 ( .A(n483), .B(KEYINPUT82), .ZN(n484) );
  XNOR2_X1 U540 ( .A(n484), .B(KEYINPUT16), .ZN(n485) );
  NOR2_X1 U541 ( .A1(n497), .A2(n485), .ZN(n518) );
  NAND2_X1 U542 ( .A1(n500), .A2(n518), .ZN(n493) );
  NOR2_X1 U543 ( .A1(n530), .A2(n493), .ZN(n487) );
  XNOR2_X1 U544 ( .A(KEYINPUT34), .B(KEYINPUT97), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U546 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  NOR2_X1 U547 ( .A1(n533), .A2(n493), .ZN(n489) );
  XOR2_X1 U548 ( .A(G8GAT), .B(n489), .Z(G1325GAT) );
  NOR2_X1 U549 ( .A1(n535), .A2(n493), .ZN(n491) );
  XNOR2_X1 U550 ( .A(KEYINPUT98), .B(KEYINPUT35), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U552 ( .A(G15GAT), .B(n492), .ZN(G1326GAT) );
  NOR2_X1 U553 ( .A1(n538), .A2(n493), .ZN(n495) );
  XNOR2_X1 U554 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(G1327GAT) );
  NOR2_X1 U556 ( .A1(n497), .A2(n496), .ZN(n498) );
  NAND2_X1 U557 ( .A1(n498), .A2(n567), .ZN(n499) );
  XNOR2_X1 U558 ( .A(KEYINPUT37), .B(n499), .ZN(n529) );
  NAND2_X1 U559 ( .A1(n500), .A2(n529), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n501), .B(KEYINPUT102), .ZN(n502) );
  XNOR2_X1 U561 ( .A(KEYINPUT38), .B(n502), .ZN(n514) );
  NOR2_X1 U562 ( .A1(n514), .A2(n530), .ZN(n506) );
  XOR2_X1 U563 ( .A(KEYINPUT100), .B(KEYINPUT103), .Z(n504) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n506), .B(n505), .ZN(G1328GAT) );
  NOR2_X1 U567 ( .A1(n533), .A2(n514), .ZN(n508) );
  XNOR2_X1 U568 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(n509), .ZN(G1329GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n511) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(KEYINPUT106), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(n513) );
  NOR2_X1 U574 ( .A1(n535), .A2(n514), .ZN(n512) );
  XOR2_X1 U575 ( .A(n513), .B(n512), .Z(G1330GAT) );
  NOR2_X1 U576 ( .A1(n538), .A2(n514), .ZN(n515) );
  XOR2_X1 U577 ( .A(G50GAT), .B(n515), .Z(G1331GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n517) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n517), .B(n516), .ZN(n520) );
  INV_X1 U581 ( .A(n546), .ZN(n576) );
  NOR2_X1 U582 ( .A1(n576), .A2(n587), .ZN(n528) );
  NAND2_X1 U583 ( .A1(n528), .A2(n518), .ZN(n524) );
  NOR2_X1 U584 ( .A1(n530), .A2(n524), .ZN(n519) );
  XOR2_X1 U585 ( .A(n520), .B(n519), .Z(n521) );
  XNOR2_X1 U586 ( .A(KEYINPUT108), .B(n521), .ZN(G1332GAT) );
  NOR2_X1 U587 ( .A1(n533), .A2(n524), .ZN(n522) );
  XOR2_X1 U588 ( .A(G64GAT), .B(n522), .Z(G1333GAT) );
  NOR2_X1 U589 ( .A1(n535), .A2(n524), .ZN(n523) );
  XOR2_X1 U590 ( .A(G71GAT), .B(n523), .Z(G1334GAT) );
  NOR2_X1 U591 ( .A1(n538), .A2(n524), .ZN(n526) );
  XNOR2_X1 U592 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U594 ( .A(G78GAT), .B(n527), .Z(G1335GAT) );
  NAND2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n537) );
  NOR2_X1 U596 ( .A1(n530), .A2(n537), .ZN(n531) );
  XOR2_X1 U597 ( .A(G85GAT), .B(n531), .Z(n532) );
  XNOR2_X1 U598 ( .A(KEYINPUT112), .B(n532), .ZN(G1336GAT) );
  NOR2_X1 U599 ( .A1(n533), .A2(n537), .ZN(n534) );
  XOR2_X1 U600 ( .A(G92GAT), .B(n534), .Z(G1337GAT) );
  NOR2_X1 U601 ( .A1(n535), .A2(n537), .ZN(n536) );
  XOR2_X1 U602 ( .A(G99GAT), .B(n536), .Z(G1338GAT) );
  NOR2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U604 ( .A(KEYINPUT44), .B(n539), .Z(n540) );
  XNOR2_X1 U605 ( .A(G106GAT), .B(n540), .ZN(G1339GAT) );
  NOR2_X1 U606 ( .A1(n558), .A2(n541), .ZN(n543) );
  NAND2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U608 ( .A(KEYINPUT114), .B(n544), .Z(n555) );
  NAND2_X1 U609 ( .A1(n587), .A2(n555), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G113GAT), .B(n545), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n548) );
  NAND2_X1 U612 ( .A1(n555), .A2(n546), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(n550) );
  XOR2_X1 U614 ( .A(G120GAT), .B(KEYINPUT115), .Z(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(G1341GAT) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n554) );
  XOR2_X1 U617 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n552) );
  NAND2_X1 U618 ( .A1(n594), .A2(n555), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1342GAT) );
  XOR2_X1 U621 ( .A(G134GAT), .B(KEYINPUT51), .Z(n557) );
  NAND2_X1 U622 ( .A1(n555), .A2(n466), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1343GAT) );
  NOR2_X1 U624 ( .A1(n584), .A2(n558), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n570) );
  NOR2_X1 U626 ( .A1(n574), .A2(n570), .ZN(n561) );
  XOR2_X1 U627 ( .A(G141GAT), .B(n561), .Z(G1344GAT) );
  NOR2_X1 U628 ( .A1(n576), .A2(n570), .ZN(n566) );
  XOR2_X1 U629 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n563) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U632 ( .A(KEYINPUT52), .B(n564), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(G1345GAT) );
  NOR2_X1 U634 ( .A1(n567), .A2(n570), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1346GAT) );
  INV_X1 U637 ( .A(n570), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U640 ( .A1(n574), .A2(n577), .ZN(n575) );
  XOR2_X1 U641 ( .A(G169GAT), .B(n575), .Z(G1348GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT56), .B(KEYINPUT123), .Z(n579) );
  XNOR2_X1 U644 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1349GAT) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT59), .ZN(n583) );
  XOR2_X1 U649 ( .A(KEYINPUT60), .B(n583), .Z(n589) );
  NOR2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(KEYINPUT125), .B(n586), .ZN(n597) );
  INV_X1 U652 ( .A(n597), .ZN(n595) );
  NAND2_X1 U653 ( .A1(n595), .A2(n587), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1352GAT) );
  XOR2_X1 U655 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n592) );
  NAND2_X1 U656 ( .A1(n595), .A2(n590), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(n593) );
  XOR2_X1 U658 ( .A(G204GAT), .B(n593), .Z(G1353GAT) );
  NAND2_X1 U659 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U660 ( .A(n596), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U661 ( .A1(n496), .A2(n597), .ZN(n598) );
  XOR2_X1 U662 ( .A(KEYINPUT62), .B(n598), .Z(n599) );
  XNOR2_X1 U663 ( .A(G218GAT), .B(n599), .ZN(G1355GAT) );
endmodule

