//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n211), .A2(new_n212), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT64), .B(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G77), .A2(G244), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n218), .B1(new_n212), .B2(new_n211), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G58), .Z(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT65), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G58), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n215), .B1(new_n219), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  AOI22_X1  g0049(.A1(new_n248), .A2(G20), .B1(G159), .B2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT7), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n255), .A2(new_n256), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT74), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n253), .A2(KEYINPUT74), .A3(new_n254), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n262), .A3(new_n207), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n257), .B1(new_n256), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G68), .ZN(new_n265));
  OAI211_X1 g0065(.A(KEYINPUT16), .B(new_n250), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT16), .ZN(new_n267));
  XOR2_X1   g0067(.A(KEYINPUT64), .B(G68), .Z(new_n268));
  AOI21_X1  g0068(.A(new_n201), .B1(new_n268), .B2(G58), .ZN(new_n269));
  INV_X1    g0069(.A(G159), .ZN(new_n270));
  INV_X1    g0070(.A(new_n249), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n269), .A2(new_n207), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n256), .B1(new_n255), .B2(G20), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n259), .A2(new_n260), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n219), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n267), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n213), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n266), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  XOR2_X1   g0080(.A(KEYINPUT8), .B(G58), .Z(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n213), .A3(new_n278), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n206), .B2(G20), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n284), .B1(new_n286), .B2(new_n282), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G274), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G1), .A3(G13), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n289), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n291), .B1(new_n294), .B2(new_n233), .ZN(new_n295));
  OAI211_X1 g0095(.A(G226), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT75), .ZN(new_n297));
  AOI21_X1  g0097(.A(G1698), .B1(new_n253), .B2(new_n254), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G223), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT75), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n255), .A2(new_n300), .A3(G226), .A4(G1698), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G87), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n297), .A2(new_n299), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n293), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n295), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(G169), .ZN(new_n306));
  AOI211_X1 g0106(.A(G179), .B(new_n295), .C1(new_n303), .C2(new_n304), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n288), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT18), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT18), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n288), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n303), .A2(new_n304), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  INV_X1    g0114(.A(new_n295), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(G200), .B2(new_n305), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n317), .A2(new_n280), .A3(new_n287), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT17), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n317), .A2(KEYINPUT17), .A3(new_n280), .A4(new_n287), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n310), .A2(new_n312), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n279), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n207), .A2(G33), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT67), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n281), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n249), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT68), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n330), .A2(new_n285), .B1(G50), .B2(new_n283), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n298), .A2(G222), .B1(new_n274), .B2(G77), .ZN(new_n333));
  INV_X1    g0133(.A(G223), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n255), .A2(G1698), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n304), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT66), .ZN(new_n338));
  AND3_X1   g0138(.A1(new_n293), .A2(new_n338), .A3(new_n289), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n338), .B1(new_n293), .B2(new_n289), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G226), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n337), .A2(new_n291), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G179), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(G169), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n332), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n332), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT9), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(KEYINPUT70), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT70), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n332), .B2(KEYINPUT9), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n351), .B(new_n353), .C1(new_n314), .C2(new_n343), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n332), .A2(KEYINPUT9), .ZN(new_n355));
  INV_X1    g0155(.A(G200), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n355), .B1(new_n344), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT10), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n354), .A2(KEYINPUT10), .A3(new_n357), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n348), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n282), .A2(new_n271), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT15), .B(G87), .ZN(new_n363));
  INV_X1    g0163(.A(G77), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n363), .A2(new_n324), .B1(new_n207), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n279), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n283), .A2(G77), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n286), .B2(G77), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n298), .A2(G232), .B1(new_n274), .B2(G107), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n220), .B2(new_n335), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n304), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n341), .A2(G244), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n291), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT69), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n374), .A2(KEYINPUT69), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n314), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n374), .A2(KEYINPUT69), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(new_n356), .A3(new_n375), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n369), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n369), .ZN(new_n382));
  OAI21_X1  g0182(.A(G179), .B1(new_n376), .B2(new_n377), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n379), .A2(G169), .A3(new_n375), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OR4_X1    g0185(.A1(new_n322), .A2(new_n361), .A3(new_n381), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT12), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n268), .A2(new_n387), .A3(new_n283), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n387), .B2(new_n283), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n286), .B2(new_n387), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n325), .A2(G77), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n219), .A2(G20), .B1(G50), .B2(new_n249), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n279), .ZN(new_n395));
  XOR2_X1   g0195(.A(KEYINPUT72), .B(KEYINPUT11), .Z(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n396), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n394), .A2(new_n279), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n391), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(G232), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n401));
  INV_X1    g0201(.A(G1698), .ZN(new_n402));
  OAI211_X1 g0202(.A(G226), .B(new_n402), .C1(new_n259), .C2(new_n260), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G97), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n401), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n304), .ZN(new_n406));
  OAI21_X1  g0206(.A(G238), .B1(new_n339), .B2(new_n340), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n407), .A3(new_n291), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(KEYINPUT13), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(KEYINPUT13), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(G190), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(KEYINPUT71), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT71), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n408), .A2(new_n414), .A3(KEYINPUT13), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n409), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n400), .B(new_n412), .C1(new_n416), .C2(new_n356), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(KEYINPUT73), .A2(G169), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT14), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n408), .A2(new_n414), .A3(KEYINPUT13), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n414), .B1(new_n408), .B2(KEYINPUT13), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n410), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT14), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n423), .A2(KEYINPUT73), .A3(new_n424), .A4(G169), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n410), .A2(G179), .A3(new_n411), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n420), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n400), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n418), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G116), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(G20), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT23), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n207), .B2(G107), .ZN(new_n434));
  INV_X1    g0234(.A(G107), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(KEYINPUT23), .A3(G20), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n432), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n255), .A2(new_n207), .A3(G87), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT22), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT22), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n255), .A2(new_n441), .A3(new_n207), .A4(G87), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n438), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n443), .A2(KEYINPUT24), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n323), .B1(new_n443), .B2(KEYINPUT24), .ZN(new_n445));
  INV_X1    g0245(.A(G13), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G1), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(G20), .A3(new_n435), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n448), .B(KEYINPUT25), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT76), .B1(new_n252), .B2(G1), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT76), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(new_n206), .A3(G33), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n453), .A2(new_n285), .A3(new_n435), .ZN(new_n454));
  OR3_X1    g0254(.A1(new_n449), .A2(KEYINPUT84), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT84), .B1(new_n449), .B2(new_n454), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n444), .A2(new_n445), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G45), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(G1), .ZN(new_n459));
  NAND2_X1  g0259(.A1(KEYINPUT5), .A2(G41), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(G264), .A3(new_n293), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n459), .B(G274), .C1(new_n462), .C2(new_n461), .ZN(new_n465));
  INV_X1    g0265(.A(G294), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n252), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G257), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(new_n253), .B2(new_n254), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n467), .B1(new_n469), .B2(G1698), .ZN(new_n470));
  OAI211_X1 g0270(.A(G250), .B(new_n402), .C1(new_n259), .C2(new_n260), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT85), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(G257), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n473));
  INV_X1    g0273(.A(new_n467), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n471), .A2(new_n473), .A3(KEYINPUT85), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n304), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n464), .B(new_n465), .C1(new_n472), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT86), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT85), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(new_n304), .A3(new_n475), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT86), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(new_n464), .A4(new_n465), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n478), .A2(G169), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n477), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G179), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n457), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n486), .A2(G200), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n478), .A2(new_n484), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(G190), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n488), .B1(new_n492), .B2(new_n457), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  INV_X1    g0294(.A(G97), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n494), .B(new_n207), .C1(G33), .C2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT83), .ZN(new_n497));
  INV_X1    g0297(.A(G116), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G20), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n279), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n497), .B1(new_n279), .B2(new_n499), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT20), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(KEYINPUT20), .B(new_n496), .C1(new_n500), .C2(new_n501), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n453), .A2(new_n285), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G116), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n283), .A2(new_n498), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n504), .A2(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n463), .A2(G270), .A3(new_n293), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n465), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT82), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n510), .A2(new_n465), .A3(KEYINPUT82), .ZN(new_n514));
  OAI211_X1 g0314(.A(G264), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n515));
  OAI211_X1 g0315(.A(G257), .B(new_n402), .C1(new_n259), .C2(new_n260), .ZN(new_n516));
  INV_X1    g0316(.A(G303), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n515), .B(new_n516), .C1(new_n517), .C2(new_n255), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n304), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n513), .A2(new_n514), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(G190), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n511), .A2(new_n512), .B1(new_n518), .B2(new_n304), .ZN(new_n522));
  AOI21_X1  g0322(.A(G200), .B1(new_n522), .B2(new_n514), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n509), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT21), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n520), .A2(G169), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n526), .B2(new_n509), .ZN(new_n527));
  INV_X1    g0327(.A(G169), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n522), .B2(new_n514), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n513), .A2(new_n514), .A3(new_n519), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n529), .A2(KEYINPUT21), .B1(new_n530), .B2(G179), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n524), .B(new_n527), .C1(new_n531), .C2(new_n509), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT4), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(G1698), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n534), .B(G244), .C1(new_n260), .C2(new_n259), .ZN(new_n535));
  INV_X1    g0335(.A(G244), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n253), .B2(new_n254), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n535), .B(new_n494), .C1(new_n537), .C2(KEYINPUT4), .ZN(new_n538));
  OAI21_X1  g0338(.A(G250), .B1(new_n259), .B2(new_n260), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n402), .B1(new_n539), .B2(KEYINPUT4), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n304), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT77), .ZN(new_n542));
  INV_X1    g0342(.A(G179), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n463), .A2(G257), .A3(new_n293), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n465), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT77), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n547), .B(new_n304), .C1(new_n538), .C2(new_n540), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n542), .A2(new_n543), .A3(new_n546), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n541), .A2(new_n546), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n528), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT6), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n552), .A2(new_n495), .A3(G107), .ZN(new_n553));
  XNOR2_X1  g0353(.A(G97), .B(G107), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n555), .A2(new_n207), .B1(new_n364), .B2(new_n271), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n435), .B1(new_n273), .B2(new_n275), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n279), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  MUX2_X1   g0358(.A(new_n283), .B(new_n506), .S(G97), .Z(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n549), .A2(new_n551), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n545), .B1(new_n541), .B2(KEYINPUT77), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n356), .B1(new_n562), .B2(new_n548), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n558), .B(new_n559), .C1(new_n550), .C2(new_n314), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n532), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(G250), .B1(new_n458), .B2(G1), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n293), .ZN(new_n570));
  OAI211_X1 g0370(.A(G244), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n571));
  OAI211_X1 g0371(.A(G238), .B(new_n402), .C1(new_n259), .C2(new_n260), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n572), .A3(new_n431), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n573), .A2(KEYINPUT78), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT78), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n571), .A2(new_n572), .A3(new_n575), .A4(new_n431), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n304), .ZN(new_n577));
  OAI211_X1 g0377(.A(G190), .B(new_n570), .C1(new_n574), .C2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n363), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(new_n283), .ZN(new_n580));
  INV_X1    g0380(.A(G87), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n453), .A2(new_n285), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n207), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(new_n495), .A3(new_n435), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT80), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n584), .A2(KEYINPUT80), .A3(new_n585), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n255), .A2(new_n207), .A3(G68), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n404), .B2(G20), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n588), .A2(new_n589), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  AOI211_X1 g0393(.A(new_n580), .B(new_n582), .C1(new_n593), .C2(new_n279), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n576), .A2(new_n304), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n573), .A2(KEYINPUT78), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n595), .A2(new_n596), .B1(new_n293), .B2(new_n569), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n578), .B(new_n594), .C1(new_n597), .C2(new_n356), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n593), .A2(new_n279), .ZN(new_n600));
  INV_X1    g0400(.A(new_n580), .ZN(new_n601));
  OR3_X1    g0401(.A1(new_n453), .A2(new_n285), .A3(new_n363), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT81), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT81), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n600), .A2(new_n605), .A3(new_n601), .A4(new_n602), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n543), .B(new_n570), .C1(new_n574), .C2(new_n577), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n597), .B2(G169), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n607), .B1(KEYINPUT79), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT79), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n608), .B(new_n611), .C1(new_n597), .C2(G169), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n599), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n493), .A2(new_n566), .A3(new_n613), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n386), .A2(new_n430), .A3(new_n614), .ZN(G372));
  AND2_X1   g0415(.A1(new_n320), .A2(new_n321), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n427), .A2(new_n428), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n385), .A2(new_n417), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n288), .A2(new_n308), .A3(new_n311), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n311), .B1(new_n288), .B2(new_n308), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI22_X1  g0424(.A1(new_n620), .A2(new_n624), .B1(new_n359), .B2(new_n360), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n348), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n386), .A2(new_n430), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT87), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n569), .A2(new_n628), .A3(new_n293), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n628), .B1(new_n569), .B2(new_n293), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n595), .B2(new_n596), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n594), .B(new_n578), .C1(new_n632), .C2(new_n356), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n608), .B(new_n603), .C1(new_n632), .C2(G169), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT88), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n549), .B2(new_n551), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n549), .A2(new_n636), .A3(new_n551), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n635), .B(new_n560), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT89), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT89), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n639), .A2(new_n643), .A3(new_n640), .ZN(new_n644));
  INV_X1    g0444(.A(new_n561), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n613), .A2(KEYINPUT26), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n642), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(G190), .B1(new_n478), .B2(new_n484), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n457), .B1(new_n648), .B2(new_n489), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n563), .A2(new_n564), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n649), .A2(new_n561), .A3(new_n650), .A4(new_n635), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n527), .B1(new_n531), .B2(new_n509), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(new_n488), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n634), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n647), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n627), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n626), .B1(new_n658), .B2(KEYINPUT90), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(KEYINPUT90), .B2(new_n658), .ZN(G369));
  INV_X1    g0460(.A(new_n652), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n447), .A2(new_n207), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n509), .A2(new_n668), .ZN(new_n669));
  MUX2_X1   g0469(.A(new_n532), .B(new_n661), .S(new_n669), .Z(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n493), .B1(new_n457), .B2(new_n668), .ZN(new_n674));
  INV_X1    g0474(.A(new_n488), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n668), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n488), .A2(new_n668), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n652), .A2(new_n668), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(G399));
  INV_X1    g0481(.A(KEYINPUT91), .ZN(new_n682));
  INV_X1    g0482(.A(new_n210), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n683), .B2(G41), .ZN(new_n684));
  INV_X1    g0484(.A(G41), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n210), .A2(KEYINPUT91), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NOR4_X1   g0487(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n216), .B2(new_n687), .ZN(new_n690));
  XOR2_X1   g0490(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n691));
  XNOR2_X1  g0491(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n656), .A2(new_n668), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT93), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT29), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n667), .B1(new_n647), .B2(new_n655), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT93), .B1(new_n697), .B2(KEYINPUT29), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n609), .A2(KEYINPUT79), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(new_n612), .A3(new_n604), .A4(new_n606), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n702), .A2(new_n645), .A3(new_n640), .A4(new_n598), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n668), .B1(new_n704), .B2(new_n654), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n699), .B1(new_n705), .B2(new_n695), .ZN(new_n706));
  OR3_X1    g0506(.A1(new_n705), .A2(new_n699), .A3(new_n695), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n696), .A2(new_n698), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n493), .A2(new_n566), .A3(new_n613), .A4(new_n668), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n513), .A2(G179), .A3(new_n514), .A4(new_n519), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n570), .B1(new_n574), .B2(new_n577), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n464), .B1(new_n472), .B2(new_n476), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n550), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n713), .A2(new_n715), .A3(KEYINPUT30), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT30), .B1(new_n713), .B2(new_n715), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n530), .A2(G179), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n562), .A2(new_n548), .ZN(new_n720));
  INV_X1    g0520(.A(new_n632), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n719), .A2(new_n477), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n668), .B1(new_n718), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n713), .A2(new_n715), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n713), .A2(new_n715), .A3(KEYINPUT30), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n722), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n667), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n724), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(G330), .B1(new_n710), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n708), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n692), .B1(new_n736), .B2(G1), .ZN(G364));
  NOR2_X1   g0537(.A1(new_n446), .A2(G20), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G45), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n687), .A2(G1), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n213), .B1(G20), .B2(new_n528), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n207), .A2(new_n314), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n356), .A2(G179), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G87), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n543), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n747), .B1(new_n247), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n543), .A2(new_n356), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n207), .A2(G190), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n274), .B(new_n750), .C1(G68), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n207), .B1(new_n756), .B2(G190), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G97), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n752), .A2(new_n756), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n270), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT32), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n744), .A2(new_n752), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n435), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n752), .A2(new_n748), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n364), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n751), .A2(new_n743), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n764), .B(new_n766), .C1(G50), .C2(new_n768), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n755), .A2(new_n759), .A3(new_n762), .A4(new_n769), .ZN(new_n770));
  XOR2_X1   g0570(.A(KEYINPUT33), .B(G317), .Z(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n753), .ZN(new_n772));
  INV_X1    g0572(.A(G322), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n274), .B1(new_n749), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n760), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n772), .B(new_n774), .C1(G329), .C2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G326), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n767), .A2(new_n777), .B1(new_n757), .B2(new_n466), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT97), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  INV_X1    g0581(.A(G283), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n782), .A2(new_n763), .B1(new_n765), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(G303), .B2(new_n746), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n776), .A2(new_n780), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n742), .B1(new_n770), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT96), .Z(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n741), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n683), .A2(new_n274), .ZN(new_n792));
  XOR2_X1   g0592(.A(G355), .B(KEYINPUT95), .Z(new_n793));
  AOI22_X1  g0593(.A1(new_n792), .A2(new_n793), .B1(new_n498), .B2(new_n683), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n217), .A2(G45), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(new_n241), .B2(G45), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n261), .A2(new_n262), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n683), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n794), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n740), .B(new_n787), .C1(new_n791), .C2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT98), .Z(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(new_n670), .B2(new_n790), .ZN(new_n803));
  INV_X1    g0603(.A(new_n740), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n673), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n671), .A2(G330), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n803), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  NAND2_X1  g0609(.A1(new_n383), .A2(new_n384), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n369), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n382), .A2(new_n668), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n381), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n385), .A2(new_n668), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n693), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n813), .A2(new_n814), .ZN(new_n817));
  AND3_X1   g0617(.A1(new_n639), .A2(new_n643), .A3(new_n640), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n643), .B1(new_n639), .B2(new_n640), .ZN(new_n819));
  AND4_X1   g0619(.A1(KEYINPUT26), .A2(new_n702), .A3(new_n598), .A4(new_n645), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n668), .B(new_n817), .C1(new_n821), .C2(new_n654), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n816), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n734), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n816), .A2(new_n735), .A3(new_n822), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n824), .A2(new_n740), .A3(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n763), .A2(new_n581), .B1(new_n760), .B2(new_n783), .ZN(new_n827));
  INV_X1    g0627(.A(new_n749), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n255), .B(new_n827), .C1(G294), .C2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n765), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G107), .A2(new_n746), .B1(new_n830), .B2(G116), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G303), .A2(new_n768), .B1(new_n754), .B2(G283), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n829), .A2(new_n759), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G143), .ZN(new_n834));
  INV_X1    g0634(.A(G150), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n834), .A2(new_n749), .B1(new_n753), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n767), .A2(new_n837), .B1(new_n765), .B2(new_n270), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n839), .A2(KEYINPUT34), .ZN(new_n840));
  INV_X1    g0640(.A(new_n797), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G58), .B2(new_n758), .ZN(new_n842));
  INV_X1    g0642(.A(G132), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n745), .A2(new_n202), .B1(new_n760), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n763), .A2(new_n265), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n842), .B(new_n846), .C1(new_n839), .C2(KEYINPUT34), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n833), .B1(new_n840), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n741), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n741), .A2(new_n788), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n740), .B1(new_n364), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n849), .B(new_n851), .C1(new_n817), .C2(new_n789), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n826), .A2(new_n852), .ZN(G384));
  INV_X1    g0653(.A(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n555), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n855), .A2(G116), .A3(new_n214), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n856), .A2(KEYINPUT99), .B1(new_n854), .B2(new_n555), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(KEYINPUT99), .B2(new_n856), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT36), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n217), .B(G77), .C1(new_n247), .C2(new_n219), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n202), .A2(G68), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n206), .B(G13), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  INV_X1    g0664(.A(new_n665), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n288), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n309), .A2(new_n866), .A3(new_n318), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n866), .B1(new_n616), .B2(new_n623), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n864), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n250), .B1(new_n264), .B2(new_n265), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n267), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(new_n279), .A3(new_n266), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n665), .B1(new_n874), .B2(new_n287), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n322), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n305), .A2(new_n543), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(G169), .B2(new_n305), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n287), .A2(new_n874), .B1(new_n878), .B2(new_n665), .ZN(new_n879));
  INV_X1    g0679(.A(new_n318), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT37), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n309), .A2(new_n866), .A3(new_n868), .A4(new_n318), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n876), .A2(KEYINPUT38), .A3(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n871), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n876), .A2(new_n883), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n864), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n886), .B1(new_n889), .B2(new_n884), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n618), .A2(new_n667), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n892), .A2(new_n893), .B1(new_n624), .B2(new_n665), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n428), .A2(new_n667), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n618), .A2(new_n417), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n427), .A2(new_n428), .A3(new_n667), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT100), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n427), .A2(KEYINPUT100), .A3(new_n428), .A4(new_n667), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n822), .B2(new_n814), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n889), .A2(new_n884), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n894), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n626), .B1(new_n708), .B2(new_n627), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n906), .B(new_n907), .Z(new_n908));
  AOI22_X1  g0708(.A1(new_n429), .A2(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n815), .B1(new_n909), .B2(new_n900), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT102), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n723), .B2(KEYINPUT31), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n730), .A2(KEYINPUT102), .A3(new_n731), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n912), .A2(new_n709), .A3(new_n724), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n910), .A2(new_n904), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n901), .A2(new_n914), .A3(new_n817), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n871), .B2(new_n884), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n915), .A2(new_n916), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n627), .A2(new_n914), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n920), .B(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(G330), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n908), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n206), .B2(new_n738), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n908), .A2(new_n923), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n863), .B1(new_n925), .B2(new_n926), .ZN(G367));
  INV_X1    g0727(.A(new_n791), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n683), .B2(new_n579), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n798), .A2(new_n237), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n740), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT104), .Z(new_n932));
  OAI22_X1  g0732(.A1(new_n753), .A2(new_n270), .B1(new_n765), .B2(new_n202), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT105), .ZN(new_n934));
  INV_X1    g0734(.A(new_n763), .ZN(new_n935));
  AOI22_X1  g0735(.A1(G58), .A2(new_n746), .B1(new_n935), .B2(G77), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n768), .A2(G143), .B1(new_n775), .B2(G137), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n757), .A2(new_n265), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n274), .B(new_n938), .C1(G150), .C2(new_n828), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n934), .A2(new_n936), .A3(new_n937), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n746), .A2(G116), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT46), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n758), .A2(G107), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n767), .A2(new_n783), .B1(new_n763), .B2(new_n495), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n797), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n753), .A2(new_n466), .B1(new_n765), .B2(new_n782), .ZN(new_n946));
  INV_X1    g0746(.A(G317), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n749), .A2(new_n517), .B1(new_n760), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n942), .A2(new_n943), .A3(new_n945), .A4(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT47), .B1(new_n940), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n940), .A2(new_n950), .A3(KEYINPUT47), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n741), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n932), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT106), .Z(new_n955));
  INV_X1    g0755(.A(new_n790), .ZN(new_n956));
  INV_X1    g0756(.A(new_n635), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n594), .A2(new_n668), .ZN(new_n958));
  MUX2_X1   g0758(.A(new_n634), .B(new_n957), .S(new_n958), .Z(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n955), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n739), .A2(G1), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n560), .B(new_n667), .C1(new_n638), .C2(new_n637), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n560), .A2(new_n667), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n650), .A2(new_n561), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n680), .A2(new_n678), .A3(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT45), .Z(new_n968));
  AOI21_X1  g0768(.A(new_n966), .B1(new_n680), .B2(new_n678), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n677), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n673), .A2(KEYINPUT103), .ZN(new_n974));
  INV_X1    g0774(.A(new_n679), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n680), .B1(new_n676), .B2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n974), .B(new_n976), .Z(new_n977));
  NAND2_X1  g0777(.A1(new_n736), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n736), .B1(new_n973), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n687), .B(KEYINPUT41), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n962), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n966), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n680), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n561), .B1(new_n983), .B2(new_n675), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n984), .A2(KEYINPUT42), .B1(new_n985), .B2(new_n668), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(KEYINPUT42), .B2(new_n984), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n677), .A2(new_n983), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n991), .B(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n961), .B1(new_n982), .B2(new_n994), .ZN(G387));
  NAND2_X1  g0795(.A1(new_n977), .A2(new_n962), .ZN(new_n996));
  INV_X1    g0796(.A(new_n688), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n792), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(G107), .B2(new_n210), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n234), .A2(G45), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT107), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n281), .A2(new_n202), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT50), .Z(new_n1003));
  AOI211_X1 g0803(.A(G45), .B(new_n997), .C1(G68), .C2(G77), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n799), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n999), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n804), .B1(new_n1006), .B2(new_n928), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n745), .A2(new_n466), .B1(new_n757), .B2(new_n782), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G322), .A2(new_n768), .B1(new_n830), .B2(G303), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n783), .B2(new_n753), .C1(new_n947), .C2(new_n749), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT108), .Z(new_n1011));
  AOI21_X1  g0811(.A(new_n1008), .B1(new_n1011), .B2(KEYINPUT48), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(KEYINPUT48), .B2(new_n1011), .ZN(new_n1013));
  XOR2_X1   g0813(.A(KEYINPUT109), .B(KEYINPUT49), .Z(new_n1014));
  XNOR2_X1  g0814(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G116), .A2(new_n935), .B1(new_n775), .B2(G326), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n841), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n746), .A2(G77), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n760), .B2(new_n835), .C1(new_n202), .C2(new_n749), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n758), .A2(new_n579), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n797), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n282), .A2(new_n753), .B1(new_n765), .B2(new_n265), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n767), .A2(new_n270), .B1(new_n763), .B2(new_n495), .ZN(new_n1023));
  OR3_X1    g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1017), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1007), .B1(new_n1025), .B2(new_n741), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n676), .B2(new_n956), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n687), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n978), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n736), .A2(new_n977), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n996), .B(new_n1027), .C1(new_n1029), .C2(new_n1030), .ZN(G393));
  OAI21_X1  g0831(.A(new_n791), .B1(new_n495), .B2(new_n210), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n799), .A2(new_n245), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n804), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n767), .A2(new_n835), .B1(new_n749), .B2(new_n270), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT51), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n282), .A2(new_n765), .B1(new_n219), .B2(new_n745), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G50), .B2(new_n754), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n758), .A2(G77), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n763), .A2(new_n581), .B1(new_n760), .B2(new_n834), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n841), .A2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1036), .A2(new_n1038), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n767), .A2(new_n947), .B1(new_n749), .B2(new_n783), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT52), .Z(new_n1044));
  OAI22_X1  g0844(.A1(new_n745), .A2(new_n782), .B1(new_n760), .B2(new_n773), .ZN(new_n1045));
  OR4_X1    g0845(.A1(new_n255), .A2(new_n1044), .A3(new_n764), .A4(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n753), .A2(new_n517), .B1(new_n765), .B2(new_n466), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G116), .B2(new_n758), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT110), .Z(new_n1049));
  OAI21_X1  g0849(.A(new_n1042), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1034), .B1(new_n1050), .B2(new_n741), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n966), .B2(new_n956), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n962), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n973), .A2(new_n978), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1028), .B1(new_n973), .B2(new_n978), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1052), .B1(new_n973), .B2(new_n1053), .C1(new_n1054), .C2(new_n1055), .ZN(G390));
  NAND3_X1  g0856(.A1(new_n627), .A2(G330), .A3(new_n914), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n814), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n697), .B2(new_n817), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n902), .B1(new_n734), .B2(new_n815), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n901), .A2(new_n914), .A3(new_n817), .A4(G330), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n914), .A2(new_n817), .A3(G330), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n735), .A2(new_n910), .B1(new_n1065), .B2(new_n902), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n668), .B(new_n813), .C1(new_n704), .C2(new_n654), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n814), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT111), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1067), .A2(KEYINPUT111), .A3(new_n814), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1066), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1064), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n907), .A2(new_n1057), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n890), .B1(new_n886), .B2(new_n885), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n903), .B2(new_n893), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1070), .A2(new_n901), .A3(new_n1071), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n885), .A2(new_n893), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n735), .A2(new_n910), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1077), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n893), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1059), .B2(new_n902), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1084), .A2(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1082), .B1(new_n1085), .B2(new_n1062), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n687), .B1(new_n1075), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1086), .B2(new_n1075), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1086), .A2(new_n1053), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n850), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n804), .B1(new_n281), .B2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n767), .A2(new_n782), .B1(new_n749), .B2(new_n498), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n845), .B(new_n1092), .C1(G294), .C2(new_n775), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1093), .A2(new_n274), .A3(new_n747), .A4(new_n1039), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n753), .A2(new_n435), .B1(new_n765), .B2(new_n495), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT112), .Z(new_n1096));
  XNOR2_X1  g0896(.A(KEYINPUT54), .B(G143), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n768), .A2(G128), .B1(new_n830), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n274), .B1(new_n828), .B2(G132), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(new_n270), .C2(new_n757), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n745), .A2(new_n835), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT53), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G137), .A2(new_n754), .B1(new_n935), .B2(G50), .ZN(new_n1104));
  INV_X1    g0904(.A(G125), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1103), .B(new_n1104), .C1(new_n1105), .C2(new_n760), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1094), .A2(new_n1096), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1091), .B1(new_n1107), .B2(new_n741), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n892), .B2(new_n789), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1088), .A2(new_n1089), .A3(new_n1109), .ZN(G378));
  NOR2_X1   g0910(.A1(new_n332), .A2(new_n665), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n361), .A2(new_n1111), .ZN(new_n1112));
  OR3_X1    g0912(.A1(new_n354), .A2(KEYINPUT10), .A3(new_n357), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n347), .B1(new_n1113), .B2(new_n358), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1111), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1112), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT116), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n920), .B2(G330), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n901), .A2(new_n914), .A3(new_n817), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n884), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT38), .B1(new_n876), .B2(new_n883), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n916), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n919), .A2(new_n910), .A3(new_n914), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1128), .A2(new_n1129), .A3(new_n1122), .A4(G330), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1121), .B1(new_n1123), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n906), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1128), .A2(new_n1129), .A3(G330), .ZN(new_n1134));
  OAI21_X1  g0934(.A(KEYINPUT115), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1117), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT115), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1112), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1134), .B1(new_n1135), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1132), .A2(new_n1133), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1121), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1134), .A2(KEYINPUT116), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n1130), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n906), .B1(new_n1146), .B2(new_n1141), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1053), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1135), .A2(new_n1140), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1149), .A2(new_n789), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n252), .A2(new_n685), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT113), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n202), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n685), .B2(new_n841), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G116), .A2(new_n768), .B1(new_n828), .B2(G107), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n938), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n935), .A2(G58), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1018), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n775), .A2(G283), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n495), .B2(new_n753), .C1(new_n363), .C2(new_n765), .ZN(new_n1160));
  NOR4_X1   g0960(.A1(new_n1158), .A2(new_n1160), .A3(G41), .A4(new_n797), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1154), .B1(new_n1161), .B2(KEYINPUT58), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n767), .A2(new_n1105), .B1(new_n753), .B2(new_n843), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1098), .A2(new_n746), .B1(new_n828), .B2(G128), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n837), .B2(new_n765), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(G150), .C2(new_n758), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1167), .A2(KEYINPUT59), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n763), .A2(new_n270), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1169), .B(new_n1152), .C1(G124), .C2(new_n775), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT59), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n1166), .B2(new_n1171), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1162), .B1(KEYINPUT58), .B2(new_n1161), .C1(new_n1168), .C2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n741), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT114), .Z(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n804), .C1(G50), .C2(new_n1090), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1150), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1148), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n707), .A2(new_n706), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n694), .B1(new_n693), .B2(new_n695), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n697), .A2(KEYINPUT93), .A3(KEYINPUT29), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1179), .B(new_n627), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1182), .A2(new_n348), .A3(new_n625), .A4(new_n1057), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1074), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1184), .B1(new_n1086), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1133), .B1(new_n1132), .B2(new_n1142), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1146), .A2(new_n906), .A3(new_n1141), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1186), .B(KEYINPUT57), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(KEYINPUT117), .A3(new_n1028), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT57), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT117), .B1(new_n1189), .B2(new_n1028), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1178), .B1(new_n1194), .B2(new_n1195), .ZN(G375));
  NAND3_X1  g0996(.A1(new_n1183), .A2(new_n1185), .A3(KEYINPUT118), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT118), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n981), .A3(new_n1075), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n804), .B1(G68), .B2(new_n1090), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n498), .A2(new_n753), .B1(new_n749), .B2(new_n782), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n255), .B(new_n1203), .C1(G77), .C2(new_n935), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G97), .A2(new_n746), .B1(new_n775), .B2(G303), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G294), .A2(new_n768), .B1(new_n830), .B2(G107), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1204), .A2(new_n1020), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G58), .A2(new_n935), .B1(new_n775), .B2(G128), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n835), .B2(new_n765), .C1(new_n270), .C2(new_n745), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n841), .B(new_n1209), .C1(G50), .C2(new_n758), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT119), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G132), .A2(new_n768), .B1(new_n754), .B2(new_n1098), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n837), .B2(new_n749), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1207), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1202), .B1(new_n1214), .B2(new_n741), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n788), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1215), .B1(new_n901), .B2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n1185), .B2(new_n1053), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1201), .A2(new_n1219), .ZN(G381));
  XNOR2_X1  g1020(.A(G375), .B(KEYINPUT121), .ZN(new_n1221));
  INV_X1    g1021(.A(G378), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(G387), .A2(G390), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  OR3_X1    g1025(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1226));
  AOI21_X1  g1026(.A(G381), .B1(new_n1226), .B2(KEYINPUT120), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(KEYINPUT120), .B2(new_n1226), .ZN(new_n1228));
  OR3_X1    g1028(.A1(new_n1223), .A2(new_n1225), .A3(new_n1228), .ZN(G407));
  OAI211_X1 g1029(.A(G407), .B(G213), .C1(G343), .C2(new_n1223), .ZN(G409));
  NAND2_X1  g1030(.A1(new_n666), .A2(G213), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT118), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1075), .A2(KEYINPUT60), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1236), .A3(new_n1197), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT60), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1028), .B1(new_n1233), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1237), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1219), .ZN(new_n1242));
  INV_X1    g1042(.A(G384), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1241), .A2(G384), .A3(new_n1219), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  OAI211_X1 g1046(.A(G378), .B(new_n1178), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n962), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1177), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(KEYINPUT122), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT122), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1148), .B2(new_n1177), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1250), .B(new_n1252), .C1(new_n980), .C2(new_n1191), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1222), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1232), .B(new_n1246), .C1(new_n1247), .C2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(KEYINPUT123), .B1(new_n1255), .B2(KEYINPUT63), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1247), .A2(new_n1254), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1246), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1231), .A3(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT123), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT63), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1256), .A2(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(G393), .B(new_n808), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G387), .A2(G390), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(new_n1266), .B2(new_n1224), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1264), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1225), .A2(new_n1268), .A3(new_n1265), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT61), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1267), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1257), .A2(new_n1231), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT124), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1232), .A2(G2897), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1244), .A2(new_n1245), .A3(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1241), .B2(new_n1219), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1243), .B(new_n1218), .C1(new_n1237), .C2(new_n1240), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1275), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1232), .B1(new_n1247), .B2(new_n1254), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n1282), .B2(KEYINPUT124), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1271), .B1(new_n1274), .B2(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1257), .A2(KEYINPUT63), .A3(new_n1258), .A4(new_n1231), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1282), .A2(KEYINPUT125), .A3(KEYINPUT63), .A4(new_n1258), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1263), .A2(new_n1284), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT126), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1263), .A2(new_n1284), .A3(KEYINPUT126), .A4(new_n1289), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  OAI221_X1 g1096(.A(new_n1270), .B1(new_n1282), .B2(new_n1281), .C1(new_n1259), .C2(KEYINPUT62), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1259), .A2(KEYINPUT62), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1294), .A2(new_n1299), .ZN(G405));
  NAND2_X1  g1100(.A1(G375), .A2(new_n1222), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1247), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1246), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n1258), .A3(new_n1247), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1295), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1295), .B1(new_n1304), .B2(new_n1303), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1305), .B1(new_n1306), .B2(KEYINPUT127), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(KEYINPUT127), .B2(new_n1306), .ZN(G402));
endmodule


