

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  INV_X1 U324 ( .A(n440), .ZN(n441) );
  XNOR2_X1 U325 ( .A(n434), .B(n402), .ZN(n403) );
  XNOR2_X1 U326 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U327 ( .A(n480), .B(KEYINPUT120), .ZN(n565) );
  XOR2_X1 U328 ( .A(n475), .B(KEYINPUT28), .Z(n527) );
  XOR2_X1 U329 ( .A(G92GAT), .B(G218GAT), .Z(n292) );
  OR2_X1 U330 ( .A1(n550), .A2(n566), .ZN(n457) );
  INV_X1 U331 ( .A(KEYINPUT95), .ZN(n420) );
  XNOR2_X1 U332 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U333 ( .A(KEYINPUT96), .B(KEYINPUT25), .ZN(n423) );
  XNOR2_X1 U334 ( .A(n424), .B(n423), .ZN(n425) );
  INV_X1 U335 ( .A(KEYINPUT91), .ZN(n400) );
  XNOR2_X1 U336 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U337 ( .A(G176GAT), .B(G64GAT), .Z(n404) );
  XNOR2_X1 U338 ( .A(n317), .B(n316), .ZN(n321) );
  NOR2_X1 U339 ( .A1(n475), .A2(n575), .ZN(n477) );
  INV_X1 U340 ( .A(n405), .ZN(n406) );
  XNOR2_X1 U341 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U342 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U343 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U344 ( .A(n409), .B(n408), .ZN(n414) );
  XOR2_X1 U345 ( .A(KEYINPUT41), .B(n465), .Z(n566) );
  INV_X1 U346 ( .A(G43GAT), .ZN(n452) );
  XNOR2_X1 U347 ( .A(n451), .B(KEYINPUT38), .ZN(n502) );
  XNOR2_X1 U348 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n483) );
  XNOR2_X1 U349 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U350 ( .A(n484), .B(n483), .ZN(G1351GAT) );
  XNOR2_X1 U351 ( .A(n455), .B(n454), .ZN(G1330GAT) );
  XOR2_X1 U352 ( .A(G141GAT), .B(G113GAT), .Z(n294) );
  XNOR2_X1 U353 ( .A(G169GAT), .B(G15GAT), .ZN(n293) );
  XNOR2_X1 U354 ( .A(n294), .B(n293), .ZN(n309) );
  XOR2_X1 U355 ( .A(KEYINPUT69), .B(G1GAT), .Z(n332) );
  XOR2_X1 U356 ( .A(G29GAT), .B(G43GAT), .Z(n296) );
  XNOR2_X1 U357 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n295) );
  XNOR2_X1 U358 ( .A(n296), .B(n295), .ZN(n435) );
  XOR2_X1 U359 ( .A(n332), .B(n435), .Z(n298) );
  XNOR2_X1 U360 ( .A(G36GAT), .B(G50GAT), .ZN(n297) );
  XNOR2_X1 U361 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U362 ( .A(KEYINPUT68), .B(G8GAT), .Z(n300) );
  NAND2_X1 U363 ( .A1(G229GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U364 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U365 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U366 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n304) );
  XNOR2_X1 U367 ( .A(G22GAT), .B(G197GAT), .ZN(n303) );
  XNOR2_X1 U368 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U369 ( .A(n305), .B(KEYINPUT67), .ZN(n306) );
  XNOR2_X1 U370 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U371 ( .A(n309), .B(n308), .Z(n550) );
  XOR2_X1 U372 ( .A(n404), .B(G92GAT), .Z(n311) );
  XOR2_X1 U373 ( .A(G148GAT), .B(G78GAT), .Z(n387) );
  XNOR2_X1 U374 ( .A(G120GAT), .B(n387), .ZN(n310) );
  XNOR2_X1 U375 ( .A(n311), .B(n310), .ZN(n317) );
  XOR2_X1 U376 ( .A(KEYINPUT31), .B(KEYINPUT71), .Z(n313) );
  XNOR2_X1 U377 ( .A(KEYINPUT32), .B(KEYINPUT70), .ZN(n312) );
  XOR2_X1 U378 ( .A(n313), .B(n312), .Z(n315) );
  NAND2_X1 U379 ( .A1(G230GAT), .A2(G233GAT), .ZN(n314) );
  XOR2_X1 U380 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n319) );
  XNOR2_X1 U381 ( .A(G204GAT), .B(KEYINPUT72), .ZN(n318) );
  XNOR2_X1 U382 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n325) );
  XNOR2_X1 U384 ( .A(G99GAT), .B(G106GAT), .ZN(n322) );
  XNOR2_X1 U385 ( .A(n322), .B(G85GAT), .ZN(n440) );
  XNOR2_X1 U386 ( .A(G71GAT), .B(G57GAT), .ZN(n323) );
  XNOR2_X1 U387 ( .A(n323), .B(KEYINPUT13), .ZN(n340) );
  XOR2_X1 U388 ( .A(n440), .B(n340), .Z(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n465) );
  INV_X1 U390 ( .A(n465), .ZN(n580) );
  NOR2_X1 U391 ( .A1(n550), .A2(n580), .ZN(n488) );
  XOR2_X1 U392 ( .A(G64GAT), .B(G78GAT), .Z(n327) );
  XOR2_X1 U393 ( .A(G15GAT), .B(G127GAT), .Z(n373) );
  XOR2_X1 U394 ( .A(G22GAT), .B(G155GAT), .Z(n392) );
  XNOR2_X1 U395 ( .A(n373), .B(n392), .ZN(n326) );
  XNOR2_X1 U396 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U397 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n329) );
  NAND2_X1 U398 ( .A1(G231GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U399 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U400 ( .A(n331), .B(n330), .Z(n334) );
  XNOR2_X1 U401 ( .A(n332), .B(KEYINPUT15), .ZN(n333) );
  XNOR2_X1 U402 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U403 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n336) );
  XNOR2_X1 U404 ( .A(KEYINPUT79), .B(KEYINPUT12), .ZN(n335) );
  XNOR2_X1 U405 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U406 ( .A(n338), .B(n337), .Z(n342) );
  XNOR2_X1 U407 ( .A(G8GAT), .B(G183GAT), .ZN(n339) );
  XNOR2_X1 U408 ( .A(n339), .B(G211GAT), .ZN(n405) );
  XNOR2_X1 U409 ( .A(n340), .B(n405), .ZN(n341) );
  XNOR2_X1 U410 ( .A(n342), .B(n341), .ZN(n584) );
  XOR2_X1 U411 ( .A(G134GAT), .B(KEYINPUT76), .Z(n438) );
  XNOR2_X1 U412 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n343) );
  XNOR2_X1 U413 ( .A(n343), .B(KEYINPUT2), .ZN(n389) );
  XOR2_X1 U414 ( .A(n438), .B(n389), .Z(n345) );
  NAND2_X1 U415 ( .A1(G225GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U416 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U417 ( .A(n346), .B(KEYINPUT5), .Z(n350) );
  XOR2_X1 U418 ( .A(G120GAT), .B(KEYINPUT0), .Z(n348) );
  XNOR2_X1 U419 ( .A(G113GAT), .B(KEYINPUT82), .ZN(n347) );
  XNOR2_X1 U420 ( .A(n348), .B(n347), .ZN(n370) );
  XNOR2_X1 U421 ( .A(n370), .B(KEYINPUT1), .ZN(n349) );
  XNOR2_X1 U422 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U423 ( .A(G85GAT), .B(G162GAT), .Z(n352) );
  XNOR2_X1 U424 ( .A(G29GAT), .B(G127GAT), .ZN(n351) );
  XNOR2_X1 U425 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U426 ( .A(n354), .B(n353), .Z(n362) );
  XOR2_X1 U427 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n356) );
  XNOR2_X1 U428 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n355) );
  XNOR2_X1 U429 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U430 ( .A(G57GAT), .B(G148GAT), .Z(n358) );
  XNOR2_X1 U431 ( .A(G1GAT), .B(G155GAT), .ZN(n357) );
  XNOR2_X1 U432 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U433 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U434 ( .A(n362), .B(n361), .ZN(n547) );
  XOR2_X1 U435 ( .A(KEYINPUT20), .B(G183GAT), .Z(n364) );
  XNOR2_X1 U436 ( .A(G134GAT), .B(G99GAT), .ZN(n363) );
  XNOR2_X1 U437 ( .A(n364), .B(n363), .ZN(n378) );
  XOR2_X1 U438 ( .A(G176GAT), .B(G71GAT), .Z(n366) );
  NAND2_X1 U439 ( .A1(G227GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U440 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U441 ( .A(n367), .B(KEYINPUT83), .Z(n372) );
  XOR2_X1 U442 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n369) );
  XNOR2_X1 U443 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n368) );
  XNOR2_X1 U444 ( .A(n369), .B(n368), .ZN(n412) );
  XNOR2_X1 U445 ( .A(n370), .B(n412), .ZN(n371) );
  XNOR2_X1 U446 ( .A(n372), .B(n371), .ZN(n374) );
  XOR2_X1 U447 ( .A(n374), .B(n373), .Z(n376) );
  XNOR2_X1 U448 ( .A(G43GAT), .B(G190GAT), .ZN(n375) );
  XNOR2_X1 U449 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U450 ( .A(n378), .B(n377), .Z(n478) );
  XOR2_X1 U451 ( .A(KEYINPUT87), .B(G204GAT), .Z(n380) );
  XNOR2_X1 U452 ( .A(G197GAT), .B(KEYINPUT85), .ZN(n379) );
  XNOR2_X1 U453 ( .A(n380), .B(n379), .ZN(n382) );
  XOR2_X1 U454 ( .A(KEYINPUT86), .B(KEYINPUT21), .Z(n381) );
  XNOR2_X1 U455 ( .A(n382), .B(n381), .ZN(n410) );
  XOR2_X1 U456 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n384) );
  XNOR2_X1 U457 ( .A(KEYINPUT24), .B(G211GAT), .ZN(n383) );
  XNOR2_X1 U458 ( .A(n384), .B(n383), .ZN(n397) );
  XOR2_X1 U459 ( .A(KEYINPUT22), .B(KEYINPUT84), .Z(n386) );
  XNOR2_X1 U460 ( .A(G218GAT), .B(G106GAT), .ZN(n385) );
  XNOR2_X1 U461 ( .A(n386), .B(n385), .ZN(n388) );
  XOR2_X1 U462 ( .A(n388), .B(n387), .Z(n395) );
  XOR2_X1 U463 ( .A(G50GAT), .B(G162GAT), .Z(n439) );
  XOR2_X1 U464 ( .A(n389), .B(n439), .Z(n391) );
  NAND2_X1 U465 ( .A1(G228GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U466 ( .A(n391), .B(n390), .ZN(n393) );
  XNOR2_X1 U467 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U468 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U469 ( .A(n397), .B(n396), .Z(n398) );
  XNOR2_X1 U470 ( .A(n410), .B(n398), .ZN(n475) );
  XNOR2_X1 U471 ( .A(G36GAT), .B(G190GAT), .ZN(n399) );
  XNOR2_X1 U472 ( .A(n292), .B(n399), .ZN(n434) );
  NAND2_X1 U473 ( .A1(G226GAT), .A2(G233GAT), .ZN(n401) );
  XOR2_X1 U474 ( .A(n403), .B(KEYINPUT92), .Z(n409) );
  XNOR2_X1 U475 ( .A(n404), .B(KEYINPUT93), .ZN(n407) );
  INV_X1 U476 ( .A(n410), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n522) );
  XOR2_X1 U479 ( .A(n522), .B(KEYINPUT94), .Z(n415) );
  XNOR2_X1 U480 ( .A(KEYINPUT27), .B(n415), .ZN(n418) );
  NAND2_X1 U481 ( .A1(n527), .A2(n418), .ZN(n533) );
  NOR2_X1 U482 ( .A1(n478), .A2(n533), .ZN(n416) );
  NOR2_X1 U483 ( .A1(n547), .A2(n416), .ZN(n428) );
  INV_X1 U484 ( .A(n478), .ZN(n531) );
  NAND2_X1 U485 ( .A1(n531), .A2(n475), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n417), .B(KEYINPUT26), .ZN(n574) );
  INV_X1 U487 ( .A(n418), .ZN(n419) );
  NOR2_X1 U488 ( .A1(n574), .A2(n419), .ZN(n549) );
  NOR2_X1 U489 ( .A1(n522), .A2(n531), .ZN(n421) );
  NOR2_X1 U490 ( .A1(n475), .A2(n422), .ZN(n424) );
  NAND2_X1 U491 ( .A1(n547), .A2(n425), .ZN(n426) );
  NOR2_X1 U492 ( .A1(n549), .A2(n426), .ZN(n427) );
  NOR2_X1 U493 ( .A1(n428), .A2(n427), .ZN(n486) );
  XNOR2_X1 U494 ( .A(KEYINPUT36), .B(KEYINPUT100), .ZN(n447) );
  XOR2_X1 U495 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n430) );
  XNOR2_X1 U496 ( .A(KEYINPUT11), .B(KEYINPUT65), .ZN(n429) );
  XNOR2_X1 U497 ( .A(n430), .B(n429), .ZN(n446) );
  XNOR2_X1 U498 ( .A(KEYINPUT74), .B(KEYINPUT10), .ZN(n432) );
  AND2_X1 U499 ( .A1(G232GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U500 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U501 ( .A(n433), .B(KEYINPUT75), .Z(n437) );
  XNOR2_X1 U502 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U503 ( .A(n437), .B(n436), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n439), .B(n438), .ZN(n442) );
  XOR2_X1 U505 ( .A(n446), .B(n445), .Z(n560) );
  XNOR2_X1 U506 ( .A(n560), .B(KEYINPUT77), .ZN(n543) );
  XNOR2_X1 U507 ( .A(n447), .B(n543), .ZN(n462) );
  NAND2_X1 U508 ( .A1(n486), .A2(n462), .ZN(n448) );
  NOR2_X1 U509 ( .A1(n584), .A2(n448), .ZN(n450) );
  XNOR2_X1 U510 ( .A(KEYINPUT101), .B(KEYINPUT37), .ZN(n449) );
  XNOR2_X1 U511 ( .A(n450), .B(n449), .ZN(n519) );
  NAND2_X1 U512 ( .A1(n488), .A2(n519), .ZN(n451) );
  NOR2_X1 U513 ( .A1(n502), .A2(n531), .ZN(n455) );
  XNOR2_X1 U514 ( .A(KEYINPUT102), .B(KEYINPUT40), .ZN(n453) );
  XOR2_X1 U515 ( .A(KEYINPUT113), .B(KEYINPUT47), .Z(n461) );
  XNOR2_X1 U516 ( .A(KEYINPUT112), .B(n584), .ZN(n570) );
  INV_X1 U517 ( .A(KEYINPUT46), .ZN(n456) );
  XNOR2_X1 U518 ( .A(n457), .B(n456), .ZN(n458) );
  NOR2_X1 U519 ( .A1(n570), .A2(n458), .ZN(n459) );
  NAND2_X1 U520 ( .A1(n459), .A2(n560), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n461), .B(n460), .ZN(n469) );
  NAND2_X1 U522 ( .A1(n462), .A2(n584), .ZN(n464) );
  XOR2_X1 U523 ( .A(KEYINPUT45), .B(KEYINPUT114), .Z(n463) );
  XNOR2_X1 U524 ( .A(n464), .B(n463), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n466), .A2(n465), .ZN(n467) );
  INV_X1 U526 ( .A(n550), .ZN(n576) );
  NOR2_X1 U527 ( .A1(n467), .A2(n576), .ZN(n468) );
  NOR2_X1 U528 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U529 ( .A(KEYINPUT48), .B(n470), .ZN(n532) );
  XNOR2_X1 U530 ( .A(n522), .B(KEYINPUT118), .ZN(n471) );
  NOR2_X1 U531 ( .A1(n532), .A2(n471), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n472), .B(KEYINPUT54), .ZN(n473) );
  NAND2_X1 U533 ( .A1(n473), .A2(n547), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n474), .B(KEYINPUT64), .ZN(n575) );
  XNOR2_X1 U535 ( .A(KEYINPUT119), .B(KEYINPUT55), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(n479) );
  NAND2_X1 U537 ( .A1(n479), .A2(n478), .ZN(n480) );
  NOR2_X1 U538 ( .A1(n565), .A2(n550), .ZN(n482) );
  XNOR2_X1 U539 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n482), .B(n481), .ZN(G1348GAT) );
  INV_X1 U541 ( .A(n565), .ZN(n569) );
  NAND2_X1 U542 ( .A1(n569), .A2(n543), .ZN(n484) );
  INV_X1 U543 ( .A(n584), .ZN(n557) );
  NOR2_X1 U544 ( .A1(n557), .A2(n543), .ZN(n485) );
  XNOR2_X1 U545 ( .A(KEYINPUT16), .B(n485), .ZN(n487) );
  AND2_X1 U546 ( .A1(n487), .A2(n486), .ZN(n505) );
  NAND2_X1 U547 ( .A1(n488), .A2(n505), .ZN(n489) );
  XOR2_X1 U548 ( .A(KEYINPUT97), .B(n489), .Z(n496) );
  NOR2_X1 U549 ( .A1(n547), .A2(n496), .ZN(n490) );
  XOR2_X1 U550 ( .A(KEYINPUT34), .B(n490), .Z(n491) );
  XNOR2_X1 U551 ( .A(G1GAT), .B(n491), .ZN(G1324GAT) );
  NOR2_X1 U552 ( .A1(n522), .A2(n496), .ZN(n492) );
  XOR2_X1 U553 ( .A(G8GAT), .B(n492), .Z(G1325GAT) );
  NOR2_X1 U554 ( .A1(n531), .A2(n496), .ZN(n494) );
  XNOR2_X1 U555 ( .A(KEYINPUT98), .B(KEYINPUT35), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U557 ( .A(G15GAT), .B(n495), .ZN(G1326GAT) );
  NOR2_X1 U558 ( .A1(n527), .A2(n496), .ZN(n498) );
  XNOR2_X1 U559 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1327GAT) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n500) );
  NOR2_X1 U562 ( .A1(n547), .A2(n502), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NOR2_X1 U564 ( .A1(n522), .A2(n502), .ZN(n501) );
  XOR2_X1 U565 ( .A(G36GAT), .B(n501), .Z(G1329GAT) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(KEYINPUT103), .ZN(n504) );
  NOR2_X1 U567 ( .A1(n527), .A2(n502), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1331GAT) );
  NOR2_X1 U569 ( .A1(n566), .A2(n576), .ZN(n518) );
  NAND2_X1 U570 ( .A1(n505), .A2(n518), .ZN(n512) );
  NOR2_X1 U571 ( .A1(n547), .A2(n512), .ZN(n507) );
  XNOR2_X1 U572 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U574 ( .A(G57GAT), .B(n508), .Z(G1332GAT) );
  NOR2_X1 U575 ( .A1(n522), .A2(n512), .ZN(n509) );
  XOR2_X1 U576 ( .A(G64GAT), .B(n509), .Z(G1333GAT) );
  NOR2_X1 U577 ( .A1(n531), .A2(n512), .ZN(n511) );
  XNOR2_X1 U578 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n510) );
  XNOR2_X1 U579 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  NOR2_X1 U580 ( .A1(n527), .A2(n512), .ZN(n517) );
  XOR2_X1 U581 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n514) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n513) );
  XNOR2_X1 U583 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U584 ( .A(KEYINPUT106), .B(n515), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n526) );
  NOR2_X1 U587 ( .A1(n547), .A2(n526), .ZN(n521) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n521), .B(n520), .ZN(G1336GAT) );
  NOR2_X1 U590 ( .A1(n522), .A2(n526), .ZN(n523) );
  XOR2_X1 U591 ( .A(KEYINPUT110), .B(n523), .Z(n524) );
  XNOR2_X1 U592 ( .A(G92GAT), .B(n524), .ZN(G1337GAT) );
  NOR2_X1 U593 ( .A1(n531), .A2(n526), .ZN(n525) );
  XOR2_X1 U594 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U595 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U596 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  NOR2_X1 U599 ( .A1(n547), .A2(n531), .ZN(n535) );
  NOR2_X1 U600 ( .A1(n532), .A2(n533), .ZN(n534) );
  NAND2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n540) );
  NOR2_X1 U602 ( .A1(n550), .A2(n540), .ZN(n536) );
  XOR2_X1 U603 ( .A(G113GAT), .B(n536), .Z(G1340GAT) );
  NOR2_X1 U604 ( .A1(n566), .A2(n540), .ZN(n538) );
  XNOR2_X1 U605 ( .A(KEYINPUT49), .B(KEYINPUT115), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U607 ( .A(G120GAT), .B(n539), .Z(G1341GAT) );
  INV_X1 U608 ( .A(n540), .ZN(n544) );
  NAND2_X1 U609 ( .A1(n570), .A2(n544), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U613 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NOR2_X1 U615 ( .A1(n547), .A2(n532), .ZN(n548) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n559) );
  NOR2_X1 U617 ( .A1(n550), .A2(n559), .ZN(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  NOR2_X1 U621 ( .A1(n566), .A2(n559), .ZN(n555) );
  XNOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n556), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n557), .A2(n559), .ZN(n558) );
  XOR2_X1 U626 ( .A(G155GAT), .B(n558), .Z(G1346GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n561), .Z(G1347GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n563) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U632 ( .A(KEYINPUT56), .B(n564), .ZN(n568) );
  NOR2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  NAND2_X1 U635 ( .A1(n569), .A2(n570), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n578) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n586) );
  NAND2_X1 U641 ( .A1(n576), .A2(n586), .ZN(n577) );
  XOR2_X1 U642 ( .A(n578), .B(n577), .Z(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT59), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n582) );
  NAND2_X1 U645 ( .A1(n586), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n586), .A2(n584), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n588) );
  NAND2_X1 U651 ( .A1(n586), .A2(n462), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

