//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n547, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G101), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(KEYINPUT66), .B1(new_n460), .B2(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(new_n463), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n459), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n460), .A2(KEYINPUT65), .A3(KEYINPUT3), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n463), .A2(G137), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n469), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND4_X1  g056(.A1(new_n468), .A2(new_n470), .A3(G2105), .A4(new_n469), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n463), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI22_X1  g060(.A1(new_n482), .A2(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n471), .A2(new_n463), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(new_n488), .B2(G136), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n468), .A2(new_n470), .A3(new_n491), .A4(new_n469), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n490), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n492), .A2(KEYINPUT4), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(G114), .B2(new_n463), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n482), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n495), .A2(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(KEYINPUT67), .B1(new_n507), .B2(G651), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n507), .A2(KEYINPUT67), .A3(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(G51), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n513), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n510), .A2(G89), .ZN(new_n524));
  NAND2_X1  g099(.A1(G63), .A2(G651), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n505), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G168));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  INV_X1    g103(.A(G52), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n511), .A2(new_n528), .B1(new_n513), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT68), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n531), .A2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  INV_X1    g111(.A(G81), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n511), .A2(new_n537), .B1(new_n513), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n533), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(KEYINPUT69), .B1(new_n539), .B2(new_n541), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n544), .A2(G860), .A3(new_n545), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT70), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  INV_X1    g126(.A(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(KEYINPUT6), .A2(G651), .ZN(new_n553));
  NAND2_X1  g128(.A1(KEYINPUT6), .A2(G651), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n555), .A2(KEYINPUT71), .A3(G53), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n505), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n557), .A2(new_n558), .B1(G651), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n511), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT72), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n562), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G168), .ZN(G286));
  NAND3_X1  g144(.A1(new_n564), .A2(G87), .A3(new_n565), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n509), .A2(G74), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(new_n555), .B2(G49), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n573), .B1(new_n570), .B2(new_n572), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(G288));
  NAND3_X1  g151(.A1(new_n564), .A2(G86), .A3(new_n565), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n505), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G48), .B2(new_n555), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(G305));
  XOR2_X1   g157(.A(KEYINPUT74), .B(G85), .Z(new_n583));
  INV_X1    g158(.A(G47), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n511), .A2(new_n583), .B1(new_n513), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n533), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n588));
  OR3_X1    g163(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n585), .B2(new_n587), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n566), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G54), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n596), .B1(new_n513), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n555), .A2(KEYINPUT76), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n505), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n598), .A2(new_n599), .B1(G651), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n592), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n592), .B1(new_n605), .B2(G868), .ZN(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  INV_X1    g183(.A(G299), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G280));
  XNOR2_X1  g185(.A(G280), .B(KEYINPUT77), .ZN(G297));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n544), .A2(new_n545), .ZN(new_n614));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n604), .A2(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n461), .A2(new_n464), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(new_n493), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT12), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2100), .Z(new_n624));
  INV_X1    g199(.A(G123), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n463), .A2(G111), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  OAI22_X1  g202(.A1(new_n482), .A2(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n488), .B2(G135), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n624), .A2(new_n630), .ZN(G156));
  INV_X1    g206(.A(G14), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT79), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n644), .B(new_n645), .Z(new_n646));
  OR2_X1    g221(.A1(new_n640), .A2(KEYINPUT79), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n640), .A2(KEYINPUT79), .ZN(new_n648));
  INV_X1    g223(.A(new_n642), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n643), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n646), .B1(new_n643), .B2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n634), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT80), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n632), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n652), .A2(new_n634), .A3(new_n653), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT81), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2067), .B(G2678), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT82), .ZN(new_n663));
  NOR2_X1   g238(.A1(G2072), .A2(G2078), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n442), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2084), .B(G2090), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n665), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n665), .B(KEYINPUT17), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n669), .B(new_n666), .C1(new_n663), .C2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n666), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n663), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n668), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n676), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT83), .ZN(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n682), .A2(new_n683), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(new_n686), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n690), .A2(new_n686), .A3(new_n684), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n693), .A2(new_n695), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n680), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(new_n680), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n700), .A2(new_n701), .A3(new_n696), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  AND3_X1   g278(.A1(new_n699), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n703), .B1(new_n699), .B2(new_n702), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(G229));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G23), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n570), .A2(new_n572), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n708), .B1(new_n710), .B2(new_n707), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G6), .B(G305), .S(G16), .Z(new_n714));
  XOR2_X1   g289(.A(KEYINPUT32), .B(G1981), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n707), .A2(G22), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G303), .B2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G1971), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n713), .A2(new_n716), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT86), .B(KEYINPUT34), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(G290), .A2(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n707), .A2(G24), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1986), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n723), .B2(new_n722), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT36), .ZN(new_n731));
  INV_X1    g306(.A(new_n482), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G119), .ZN(new_n733));
  OR2_X1    g308(.A1(G95), .A2(G2105), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n734), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n735));
  INV_X1    g310(.A(G131), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n733), .B(new_n735), .C1(new_n736), .C2(new_n487), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT84), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  MUX2_X1   g316(.A(G25), .B(new_n741), .S(G29), .Z(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT85), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT35), .B(G1991), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(KEYINPUT85), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n743), .A2(new_n745), .ZN(new_n747));
  INV_X1    g322(.A(new_n744), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n730), .A2(new_n731), .A3(new_n746), .A4(new_n749), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n749), .A2(new_n724), .A3(new_n729), .A4(new_n746), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(KEYINPUT36), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n707), .A2(G20), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT23), .Z(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G299), .B2(G16), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1956), .ZN(new_n757));
  INV_X1    g332(.A(G29), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G35), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G162), .B2(new_n758), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT29), .Z(new_n761));
  INV_X1    g336(.A(G2090), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n757), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT94), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G4), .A2(G16), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n605), .B2(G16), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT87), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n604), .A2(new_n707), .ZN(new_n770));
  OAI21_X1  g345(.A(KEYINPUT87), .B1(new_n770), .B2(new_n766), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G1348), .ZN(new_n773));
  INV_X1    g348(.A(G1348), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n769), .A2(new_n774), .A3(new_n771), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n758), .A2(G33), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT90), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT25), .Z(new_n780));
  NAND2_X1  g355(.A1(G115), .A2(G2104), .ZN(new_n781));
  INV_X1    g356(.A(G127), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n476), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n780), .B1(G2105), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n488), .A2(G139), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n777), .B1(new_n786), .B2(new_n758), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(G2072), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(G2072), .ZN(new_n789));
  NOR2_X1   g364(.A1(G27), .A2(G29), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G164), .B2(G29), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(G2078), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n788), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n707), .A2(G5), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G171), .B2(new_n707), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(G1961), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n707), .A2(G19), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n614), .B2(G16), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT88), .B(G1341), .Z(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n795), .A2(G1961), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n791), .A2(G2078), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n796), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n761), .A2(new_n762), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n488), .A2(G141), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n732), .A2(G129), .ZN(new_n806));
  NAND3_X1  g381(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT26), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G105), .B2(new_n620), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n805), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G29), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(KEYINPUT92), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n812), .B(KEYINPUT92), .C1(G29), .C2(G32), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT27), .B(G1996), .Z(new_n815));
  AND3_X1   g390(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n815), .B1(new_n813), .B2(new_n814), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n804), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n793), .A2(new_n803), .A3(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n707), .A2(G21), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G286), .B2(G16), .ZN(new_n821));
  INV_X1    g396(.A(G1966), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT93), .Z(new_n824));
  INV_X1    g399(.A(G2084), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n758), .B1(KEYINPUT24), .B2(G34), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(KEYINPUT24), .B2(G34), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n480), .B2(G29), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n824), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT30), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n830), .A2(G28), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n758), .B1(new_n830), .B2(G28), .ZN(new_n832));
  AND2_X1   g407(.A1(KEYINPUT31), .A2(G11), .ZN(new_n833));
  NOR2_X1   g408(.A1(KEYINPUT31), .A2(G11), .ZN(new_n834));
  OAI22_X1  g409(.A1(new_n831), .A2(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n629), .B2(G29), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n821), .B2(new_n822), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n798), .B2(new_n799), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n828), .A2(new_n825), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT91), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n758), .A2(G26), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT28), .ZN(new_n842));
  OAI21_X1  g417(.A(KEYINPUT89), .B1(G104), .B2(G2105), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NOR3_X1   g419(.A1(KEYINPUT89), .A2(G104), .A3(G2105), .ZN(new_n845));
  OAI221_X1 g420(.A(G2104), .B1(G116), .B2(new_n463), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G128), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n847), .B2(new_n482), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G140), .B2(new_n488), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n842), .B1(new_n849), .B2(new_n758), .ZN(new_n850));
  INV_X1    g425(.A(G2067), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  AND4_X1   g427(.A1(new_n829), .A2(new_n838), .A3(new_n840), .A4(new_n852), .ZN(new_n853));
  AND4_X1   g428(.A1(new_n765), .A2(new_n776), .A3(new_n819), .A4(new_n853), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n753), .A2(new_n854), .A3(KEYINPUT95), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT95), .B1(new_n753), .B2(new_n854), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(G311));
  INV_X1    g432(.A(KEYINPUT96), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n753), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n858), .B1(new_n753), .B2(new_n854), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(G150));
  XOR2_X1   g436(.A(KEYINPUT97), .B(G93), .Z(new_n862));
  INV_X1    g437(.A(G55), .ZN(new_n863));
  OAI22_X1  g438(.A1(new_n511), .A2(new_n862), .B1(new_n513), .B2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT98), .Z(new_n865));
  AOI22_X1  g440(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(new_n533), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n614), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n865), .A2(new_n542), .A3(new_n867), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n605), .A2(G559), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n875));
  AOI21_X1  g450(.A(G860), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n875), .B2(new_n874), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n868), .A2(G860), .ZN(new_n878));
  XOR2_X1   g453(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(G145));
  XNOR2_X1  g456(.A(new_n629), .B(new_n480), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(G162), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n739), .A2(KEYINPUT100), .A3(new_n740), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT100), .B1(new_n739), .B2(new_n740), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n622), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  INV_X1    g463(.A(new_n622), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n889), .A3(new_n884), .ZN(new_n890));
  INV_X1    g465(.A(G130), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n463), .A2(G118), .ZN(new_n892));
  OAI21_X1  g467(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n893));
  OAI22_X1  g468(.A1(new_n482), .A2(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(new_n488), .B2(G142), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n887), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n895), .B1(new_n887), .B2(new_n890), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n786), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n849), .B(G164), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n811), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n900), .A2(new_n811), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n900), .A2(new_n811), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(new_n786), .A3(new_n901), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n883), .B1(new_n898), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n907), .B1(new_n896), .B2(new_n897), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(KEYINPUT101), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT101), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n907), .B(new_n913), .C1(new_n896), .C2(new_n897), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n912), .A2(new_n914), .B1(new_n898), .B2(new_n908), .ZN(new_n915));
  INV_X1    g490(.A(new_n883), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g493(.A1(new_n868), .A2(new_n615), .ZN(new_n919));
  XNOR2_X1  g494(.A(G303), .B(G305), .ZN(new_n920));
  XNOR2_X1  g495(.A(G290), .B(new_n709), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n921), .B2(KEYINPUT102), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(KEYINPUT102), .B2(new_n921), .ZN(new_n923));
  INV_X1    g498(.A(new_n921), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(new_n920), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n928), .A2(KEYINPUT42), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(KEYINPUT42), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n927), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n930), .B1(new_n927), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n605), .A2(new_n609), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n609), .B1(new_n595), .B2(new_n603), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(KEYINPUT41), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n604), .A2(G299), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n939), .B1(new_n940), .B2(new_n936), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n617), .B(new_n871), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n940), .A2(new_n936), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n934), .B(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n919), .B1(new_n948), .B2(new_n615), .ZN(G295));
  OAI21_X1  g524(.A(new_n919), .B1(new_n948), .B2(new_n615), .ZN(G331));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n951));
  NAND2_X1  g526(.A1(G286), .A2(KEYINPUT104), .ZN(new_n952));
  OR2_X1    g527(.A1(G286), .A2(KEYINPUT104), .ZN(new_n953));
  NAND3_X1  g528(.A1(G171), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(G301), .A2(KEYINPUT104), .A3(G286), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n956), .A2(new_n871), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n871), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n938), .B(new_n941), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n958), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n871), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n945), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(G37), .B1(new_n963), .B2(new_n927), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n959), .A2(new_n962), .A3(new_n926), .A4(new_n923), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n965), .B1(new_n964), .B2(new_n966), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n951), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n964), .A2(new_n966), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(KEYINPUT44), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(G397));
  XNOR2_X1  g549(.A(new_n849), .B(new_n851), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT105), .B(G40), .ZN(new_n976));
  INV_X1    g551(.A(new_n474), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n493), .B2(G125), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n976), .B1(new_n978), .B2(new_n463), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n620), .A2(G101), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n472), .A2(new_n468), .A3(new_n469), .A4(new_n470), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT106), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n473), .A2(new_n479), .A3(new_n984), .A4(new_n976), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(new_n495), .B2(new_n500), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n975), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n975), .A2(new_n992), .A3(KEYINPUT109), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n810), .B(G1996), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n992), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n741), .A2(new_n748), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n744), .B1(new_n739), .B2(new_n740), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n992), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G290), .A2(G1986), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT108), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT107), .ZN(new_n1007));
  OR3_X1    g582(.A1(G290), .A2(new_n1007), .A3(G1986), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1007), .B1(G290), .B2(G1986), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1004), .B1(new_n992), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n500), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n493), .A2(new_n494), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n990), .A2(G1384), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n983), .A2(new_n985), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1966), .B1(new_n1019), .B2(new_n991), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n989), .A2(KEYINPUT50), .ZN(new_n1021));
  NOR2_X1   g596(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT114), .B(G2084), .Z(new_n1024));
  AND4_X1   g599(.A1(new_n986), .A2(new_n1021), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT120), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n986), .A2(new_n991), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n822), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n986), .A2(new_n1023), .A3(new_n1021), .A4(new_n1024), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1026), .A2(G168), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G286), .A2(G8), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1034), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(G8), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1037), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT62), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1038), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1041), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT62), .B1(new_n1048), .B2(new_n1045), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n986), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1050));
  INV_X1    g625(.A(G1961), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(G2078), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1052), .B1(new_n1055), .B2(new_n1028), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n991), .A2(KEYINPUT110), .ZN(new_n1057));
  INV_X1    g632(.A(G2078), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n989), .A2(new_n1059), .A3(new_n990), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1019), .A2(new_n1057), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1053), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT121), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1064), .A3(new_n1053), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1056), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(G301), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n989), .B1(new_n983), .B2(new_n985), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n570), .A2(G1976), .A3(new_n572), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1068), .A2(new_n1069), .A3(new_n1035), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT113), .B(G1976), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(G288), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1981), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n577), .A2(new_n581), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n555), .A2(G48), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n509), .A2(new_n510), .A3(G86), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1077), .B(new_n1078), .C1(new_n1079), .C2(new_n533), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G1981), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1076), .A2(KEYINPUT49), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT49), .B1(new_n1076), .B2(new_n1081), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1068), .A2(new_n1035), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1074), .A2(new_n1070), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n986), .A2(new_n1060), .A3(new_n1027), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1059), .B1(new_n989), .B2(new_n990), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n719), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n986), .A2(new_n1023), .A3(new_n1021), .A4(new_n762), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1035), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1035), .B1(new_n516), .B2(new_n517), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n1093));
  OR2_X1    g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1092), .B1(KEYINPUT112), .B2(KEYINPUT55), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1072), .B(new_n1086), .C1(new_n1091), .C2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT111), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1089), .A2(new_n1098), .A3(new_n1090), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1099), .A2(new_n1100), .A3(new_n1035), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1097), .B1(new_n1101), .B2(new_n1096), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1047), .A2(new_n1049), .A3(new_n1067), .A4(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT123), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1084), .A2(G1976), .A3(G288), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1076), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1085), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT111), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1089), .A2(new_n1098), .A3(new_n1090), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1109), .A2(G8), .A3(new_n1096), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1086), .A2(new_n1072), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1107), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1097), .ZN(new_n1114));
  AOI211_X1 g689(.A(new_n1035), .B(G286), .C1(new_n1029), .C2(new_n1031), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(new_n1111), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT63), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1109), .A2(G8), .A3(new_n1110), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1120), .A2(new_n1111), .A3(new_n1115), .A4(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1113), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1067), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1104), .A2(new_n1123), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n1128));
  INV_X1    g703(.A(G40), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n480), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(G160), .A2(KEYINPUT122), .A3(G40), .ZN(new_n1131));
  AND4_X1   g706(.A1(new_n1027), .A2(new_n1130), .A3(new_n1131), .A4(new_n1054), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1132), .A2(new_n991), .B1(new_n1051), .B2(new_n1050), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1065), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1064), .B1(new_n1061), .B2(new_n1053), .ZN(new_n1135));
  OAI211_X1 g710(.A(G301), .B(new_n1133), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1066), .B2(G301), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT54), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1056), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1140), .B(G301), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1132), .A2(new_n991), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1052), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1143), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1141), .B(KEYINPUT54), .C1(new_n1144), .C2(G301), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1139), .A2(new_n1145), .A3(new_n1146), .A4(new_n1102), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1050), .A2(new_n774), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1068), .A2(new_n851), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1150), .A2(KEYINPUT116), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT116), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT60), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1151), .A2(KEYINPUT60), .A3(new_n1153), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1154), .B1(new_n1155), .B2(new_n604), .ZN(new_n1156));
  OAI211_X1 g731(.A(KEYINPUT60), .B(new_n605), .C1(new_n1151), .C2(new_n1153), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(KEYINPUT56), .B(G2072), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1019), .A2(new_n1057), .A3(new_n1060), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(G1956), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1050), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1163), .A2(KEYINPUT117), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1163), .A2(KEYINPUT117), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT57), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT115), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n562), .A2(new_n567), .A3(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1166), .A2(KEYINPUT115), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OR3_X1    g747(.A1(new_n1164), .A2(new_n1165), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT119), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1172), .A2(new_n1162), .A3(new_n1160), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1173), .A2(new_n1174), .A3(KEYINPUT61), .A4(new_n1175), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1164), .A2(new_n1165), .A3(new_n1172), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(KEYINPUT61), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT119), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1163), .B1(new_n1171), .B2(new_n1170), .ZN(new_n1180));
  AOI21_X1  g755(.A(KEYINPUT61), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1019), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1182));
  XNOR2_X1  g757(.A(KEYINPUT58), .B(G1341), .ZN(new_n1183));
  OAI22_X1  g758(.A1(new_n1182), .A2(G1996), .B1(new_n1068), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n614), .B1(KEYINPUT118), .B2(KEYINPUT59), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1186), .B1(KEYINPUT118), .B2(KEYINPUT59), .ZN(new_n1187));
  NOR2_X1   g762(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1184), .A2(new_n1185), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1181), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1158), .A2(new_n1176), .A3(new_n1179), .A4(new_n1190), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n1151), .A2(new_n604), .A3(new_n1153), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1175), .B1(new_n1177), .B2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1147), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1012), .B1(new_n1127), .B2(new_n1194), .ZN(new_n1195));
  NOR3_X1   g770(.A1(new_n987), .A2(G1996), .A3(new_n991), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT46), .Z(new_n1197));
  OAI21_X1  g772(.A(new_n992), .B1(new_n975), .B2(new_n810), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g774(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1199), .B(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1008), .A2(new_n992), .A3(new_n1009), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT48), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1203), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1204));
  AND2_X1   g779(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1205));
  AND3_X1   g780(.A1(new_n997), .A2(new_n1001), .A3(new_n999), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n849), .A2(new_n851), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n992), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(KEYINPUT124), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n1210));
  OAI211_X1 g785(.A(new_n1210), .B(new_n992), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1211));
  NAND4_X1  g786(.A1(new_n1205), .A2(KEYINPUT126), .A3(new_n1209), .A4(new_n1211), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1209), .A2(new_n1211), .A3(new_n1201), .A4(new_n1204), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1195), .A2(new_n1216), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g792(.A1(new_n677), .A2(G319), .A3(new_n678), .ZN(new_n1219));
  XNOR2_X1  g793(.A(new_n1219), .B(KEYINPUT127), .ZN(new_n1220));
  OAI21_X1  g794(.A(new_n1220), .B1(new_n704), .B2(new_n705), .ZN(new_n1221));
  AOI21_X1  g795(.A(new_n1221), .B1(new_n658), .B2(new_n660), .ZN(new_n1222));
  OAI211_X1 g796(.A(new_n917), .B(new_n1222), .C1(new_n967), .C2(new_n968), .ZN(G225));
  INV_X1    g797(.A(G225), .ZN(G308));
endmodule


