//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT32), .ZN(new_n203));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT23), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n210), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT24), .ZN(new_n213));
  NOR2_X1   g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n211), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT25), .B1(new_n209), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n208), .A2(new_n217), .A3(new_n206), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G176gat), .ZN(new_n220));
  INV_X1    g019(.A(G169gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(KEYINPUT23), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT27), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(G183gat), .ZN(new_n225));
  INV_X1    g024(.A(G183gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(KEYINPUT27), .ZN(new_n227));
  INV_X1    g026(.A(G190gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT28), .ZN(new_n229));
  NOR3_X1   g028(.A1(new_n225), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(KEYINPUT27), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT27), .B(G183gat), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n228), .B(new_n233), .C1(new_n234), .C2(new_n232), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT28), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n230), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT26), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n239), .B2(new_n204), .ZN(new_n240));
  INV_X1    g039(.A(G176gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT26), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(new_n212), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n216), .B(new_n223), .C1(new_n237), .C2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247));
  OAI21_X1  g046(.A(G127gat), .B1(new_n247), .B2(KEYINPUT1), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n249));
  INV_X1    g048(.A(G127gat), .ZN(new_n250));
  INV_X1    g049(.A(G113gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(G120gat), .ZN(new_n252));
  INV_X1    g051(.A(G120gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(G113gat), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n249), .B(new_n250), .C1(new_n252), .C2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(G134gat), .B1(new_n248), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n248), .A2(new_n255), .A3(G134gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT67), .B1(new_n246), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n246), .A2(new_n259), .ZN(new_n261));
  INV_X1    g060(.A(new_n258), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(new_n256), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n240), .A2(new_n243), .B1(G183gat), .B2(G190gat), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT66), .B1(new_n225), .B2(new_n227), .ZN(new_n266));
  AOI21_X1  g065(.A(G190gat), .B1(new_n231), .B2(new_n232), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT28), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n265), .B1(new_n268), .B2(new_n230), .ZN(new_n269));
  INV_X1    g068(.A(new_n214), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(KEYINPUT24), .A3(new_n212), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n238), .B1(new_n242), .B2(new_n207), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n211), .A4(new_n205), .ZN(new_n273));
  AOI22_X1  g072(.A1(KEYINPUT25), .A2(new_n273), .B1(new_n219), .B2(new_n222), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n263), .A2(new_n264), .A3(new_n269), .A4(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n260), .A2(new_n261), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G227gat), .A2(G233gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT64), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n203), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT33), .ZN(new_n280));
  XNOR2_X1  g079(.A(G15gat), .B(G43gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT68), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(G71gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(G99gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n279), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT33), .B1(new_n276), .B2(new_n278), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n287));
  NOR4_X1   g086(.A1(new_n279), .A2(new_n286), .A3(new_n287), .A4(new_n284), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n276), .A2(new_n278), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n284), .B1(new_n289), .B2(new_n280), .ZN(new_n290));
  INV_X1    g089(.A(new_n279), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT69), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n285), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT34), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n276), .A2(new_n278), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT34), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n296), .B(new_n285), .C1(new_n288), .C2(new_n292), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n294), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n295), .B1(new_n294), .B2(new_n297), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n202), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n290), .A2(new_n291), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n287), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n290), .A2(KEYINPUT69), .A3(new_n291), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n296), .B1(new_n304), .B2(new_n285), .ZN(new_n305));
  INV_X1    g104(.A(new_n297), .ZN(new_n306));
  OAI22_X1  g105(.A1(new_n305), .A2(new_n306), .B1(new_n278), .B2(new_n276), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n294), .A2(new_n295), .A3(new_n297), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(KEYINPUT95), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT81), .ZN(new_n310));
  INV_X1    g109(.A(G148gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(G141gat), .ZN(new_n312));
  INV_X1    g111(.A(G141gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(KEYINPUT81), .A3(G148gat), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n312), .B(new_n314), .C1(new_n313), .C2(G148gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  INV_X1    g115(.A(G155gat), .ZN(new_n317));
  INV_X1    g116(.A(G162gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n316), .B1(new_n319), .B2(KEYINPUT2), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT79), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT79), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n319), .A2(new_n325), .A3(new_n316), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT80), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n316), .A2(KEYINPUT2), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n311), .A2(G141gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n313), .A2(G148gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n327), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n328), .B1(new_n327), .B2(new_n332), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n321), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G197gat), .ZN(new_n336));
  INV_X1    g135(.A(G204gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G197gat), .A2(G204gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT22), .ZN(new_n340));
  NAND2_X1  g139(.A1(G211gat), .A2(G218gat), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n338), .A2(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(G211gat), .A2(G218gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(G211gat), .A2(G218gat), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT71), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT71), .ZN(new_n346));
  INV_X1    g145(.A(G211gat), .ZN(new_n347));
  INV_X1    g146(.A(G218gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n346), .B1(new_n349), .B2(new_n341), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n342), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n341), .A2(new_n340), .ZN(new_n352));
  NOR2_X1   g151(.A1(G197gat), .A2(G204gat), .ZN(new_n353));
  AND2_X1   g152(.A1(G197gat), .A2(G204gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT71), .B1(new_n343), .B2(new_n344), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n349), .A2(new_n346), .A3(new_n341), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT29), .B1(new_n351), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n335), .B1(KEYINPUT3), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT88), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n363), .B(new_n321), .C1(new_n333), .C2(new_n334), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n358), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n335), .B(KEYINPUT88), .C1(KEYINPUT3), .C2(new_n359), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n362), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT87), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n355), .A2(new_n356), .A3(new_n357), .A4(new_n375), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n376), .A2(new_n365), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n351), .A2(KEYINPUT87), .A3(new_n358), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT3), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n321), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n327), .A2(new_n332), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT80), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n327), .A2(new_n328), .A3(new_n332), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n380), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n372), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n367), .B1(new_n364), .B2(new_n365), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n374), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT31), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT31), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n391), .A3(new_n388), .ZN(new_n392));
  XOR2_X1   g191(.A(G78gat), .B(G106gat), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n390), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n391), .B1(new_n374), .B2(new_n388), .ZN(new_n396));
  AOI211_X1 g195(.A(KEYINPUT31), .B(new_n387), .C1(new_n371), .C2(new_n373), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n393), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G22gat), .B(G50gat), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n395), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n395), .B2(new_n398), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n335), .A2(new_n259), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(KEYINPUT84), .A3(new_n405), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT4), .B1(new_n335), .B2(new_n259), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n335), .A2(KEYINPUT3), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n412), .A2(new_n259), .A3(new_n364), .ZN(new_n413));
  NAND2_X1  g212(.A1(G225gat), .A2(G233gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n415), .B1(new_n406), .B2(new_n410), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n384), .B(new_n259), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n417), .B1(new_n421), .B2(new_n414), .ZN(new_n422));
  OAI22_X1  g221(.A1(new_n411), .A2(new_n419), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G57gat), .B(G85gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(G1gat), .B(G29gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  XOR2_X1   g229(.A(KEYINPUT85), .B(KEYINPUT6), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT86), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n423), .A2(new_n434), .A3(new_n429), .A4(new_n431), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(new_n418), .A3(new_n416), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n437), .B(new_n428), .C1(new_n422), .C2(new_n420), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n430), .A2(new_n432), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n433), .A2(new_n435), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n300), .A2(new_n309), .A3(new_n403), .A4(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT29), .B1(new_n274), .B2(new_n269), .ZN(new_n442));
  INV_X1    g241(.A(G226gat), .ZN(new_n443));
  INV_X1    g242(.A(G233gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT72), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n445), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(new_n274), .B2(new_n269), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n235), .A2(new_n236), .ZN(new_n449));
  INV_X1    g248(.A(new_n230), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n245), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n223), .A2(new_n216), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n365), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n448), .B1(new_n453), .B2(new_n447), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n367), .B(new_n446), .C1(new_n454), .C2(KEYINPUT72), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT73), .ZN(new_n456));
  INV_X1    g255(.A(new_n454), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n368), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT72), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n442), .A2(new_n445), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n459), .B1(new_n460), .B2(new_n448), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT73), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n367), .A4(new_n446), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n456), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT74), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n456), .A2(KEYINPUT74), .A3(new_n463), .A4(new_n458), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(G8gat), .B(G36gat), .Z(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(G64gat), .ZN(new_n470));
  INV_X1    g269(.A(G92gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT75), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n468), .A2(KEYINPUT75), .A3(new_n472), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT89), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT30), .ZN(new_n479));
  INV_X1    g278(.A(new_n472), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n456), .A2(new_n458), .A3(new_n463), .A4(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n481), .A2(KEYINPUT78), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(KEYINPUT78), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n479), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n456), .A2(new_n458), .A3(new_n463), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT76), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT30), .A4(new_n480), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT76), .B1(new_n481), .B2(new_n479), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n477), .A2(new_n478), .A3(new_n484), .A4(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT75), .B1(new_n468), .B2(new_n472), .ZN(new_n491));
  AOI211_X1 g290(.A(new_n474), .B(new_n480), .C1(new_n466), .C2(new_n467), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n484), .B(new_n489), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT89), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n441), .A2(new_n495), .A3(KEYINPUT35), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT35), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n440), .A2(new_n484), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT77), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT77), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n501), .B(new_n489), .C1(new_n491), .C2(new_n492), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n298), .A2(new_n299), .A3(new_n402), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n497), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT70), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT36), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n307), .A2(new_n506), .A3(new_n507), .A4(new_n308), .ZN(new_n508));
  NOR2_X1   g307(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n510), .B(new_n511), .C1(new_n298), .C2(new_n299), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n508), .B(new_n512), .C1(new_n503), .C2(new_n403), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n433), .A2(new_n435), .A3(new_n439), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n482), .A2(new_n483), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n472), .B1(new_n464), .B2(KEYINPUT37), .ZN(new_n518));
  AOI211_X1 g317(.A(new_n517), .B(new_n518), .C1(new_n468), .C2(KEYINPUT37), .ZN(new_n519));
  INV_X1    g318(.A(new_n461), .ZN(new_n520));
  INV_X1    g319(.A(new_n446), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n368), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT93), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT92), .B1(new_n457), .B2(new_n368), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n525), .B(new_n368), .C1(new_n520), .C2(new_n521), .ZN(new_n526));
  OR3_X1    g325(.A1(new_n457), .A2(KEYINPUT92), .A3(new_n368), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n523), .A2(new_n524), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT37), .ZN(new_n529));
  INV_X1    g328(.A(new_n518), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n516), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n514), .B(new_n515), .C1(new_n519), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n403), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT39), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n436), .A2(new_n413), .ZN(new_n535));
  INV_X1    g334(.A(new_n414), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT90), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT90), .ZN(new_n538));
  AOI211_X1 g337(.A(new_n538), .B(new_n414), .C1(new_n436), .C2(new_n413), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n534), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n412), .A2(new_n259), .A3(new_n364), .ZN(new_n541));
  INV_X1    g340(.A(new_n410), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n542), .B1(new_n407), .B2(new_n406), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n541), .B1(new_n543), .B2(new_n409), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n538), .B1(new_n544), .B2(new_n414), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n535), .A2(KEYINPUT90), .A3(new_n536), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n534), .B1(new_n421), .B2(new_n414), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n540), .A2(new_n548), .A3(new_n428), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT40), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(KEYINPUT91), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n430), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n549), .A2(new_n550), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT91), .B1(new_n549), .B2(new_n550), .ZN(new_n554));
  NOR3_X1   g353(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n533), .B1(new_n495), .B2(new_n555), .ZN(new_n556));
  OAI22_X1  g355(.A1(new_n496), .A2(new_n505), .B1(new_n513), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G8gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(G15gat), .B(G22gat), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n559), .A2(G1gat), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n558), .B1(new_n560), .B2(KEYINPUT98), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT16), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n559), .B1(new_n562), .B2(G1gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n561), .B(new_n564), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n567));
  XOR2_X1   g366(.A(G43gat), .B(G50gat), .Z(new_n568));
  INV_X1    g367(.A(KEYINPUT15), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G29gat), .A2(G36gat), .ZN(new_n571));
  NOR3_X1   g370(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n570), .B(new_n571), .C1(new_n572), .C2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n568), .A2(new_n569), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n566), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(KEYINPUT17), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n578), .B1(new_n579), .B2(new_n565), .ZN(new_n580));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT18), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n565), .B(new_n577), .Z(new_n585));
  XOR2_X1   g384(.A(new_n581), .B(KEYINPUT13), .Z(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n580), .A2(KEYINPUT18), .A3(new_n581), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n584), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT96), .B(KEYINPUT11), .ZN(new_n590));
  XNOR2_X1  g389(.A(G113gat), .B(G141gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G169gat), .B(G197gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n594), .B(KEYINPUT12), .Z(new_n595));
  OR2_X1    g394(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n589), .A2(new_n595), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G71gat), .B(G78gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(G57gat), .ZN(new_n602));
  OR3_X1    g401(.A1(new_n602), .A2(KEYINPUT99), .A3(G64gat), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT99), .B1(new_n602), .B2(G64gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n602), .A2(G64gat), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT100), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n601), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT9), .ZN(new_n609));
  INV_X1    g408(.A(G71gat), .ZN(new_n610));
  INV_X1    g409(.A(G78gat), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n608), .B(new_n612), .C1(new_n607), .C2(new_n606), .ZN(new_n613));
  XNOR2_X1  g412(.A(G57gat), .B(G64gat), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n601), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G99gat), .B(G106gat), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n613), .B(new_n615), .C1(KEYINPUT103), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G85gat), .A2(G92gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT7), .ZN(new_n619));
  NAND2_X1  g418(.A1(G99gat), .A2(G106gat), .ZN(new_n620));
  INV_X1    g419(.A(G85gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(KEYINPUT8), .A2(new_n620), .B1(new_n621), .B2(new_n471), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(new_n616), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n617), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n613), .A2(new_n615), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(KEYINPUT10), .ZN(new_n628));
  OAI22_X1  g427(.A1(new_n626), .A2(KEYINPUT10), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n625), .A2(new_n631), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(new_n241), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(new_n337), .ZN(new_n636));
  OR3_X1    g435(.A1(new_n632), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n636), .B1(new_n632), .B2(new_n633), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n599), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n624), .B(KEYINPUT102), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n579), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(G232gat), .A2(G233gat), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n577), .A2(new_n624), .B1(KEYINPUT41), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G134gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G190gat), .B(G218gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n643), .A2(KEYINPUT41), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G162gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n648), .B(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT21), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n627), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n250), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n565), .B1(new_n627), .B2(new_n653), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n658));
  XNOR2_X1  g457(.A(G183gat), .B(G211gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n658), .B(new_n659), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n657), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT101), .B(G155gat), .Z(new_n662));
  NAND2_X1  g461(.A1(G231gat), .A2(G233gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(new_n665), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n652), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n557), .A2(new_n640), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n440), .B(KEYINPUT105), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g475(.A1(new_n562), .A2(new_n558), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n562), .A2(new_n558), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n672), .A2(new_n495), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n672), .A2(new_n495), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(G8gat), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n680), .ZN(new_n683));
  MUX2_X1   g482(.A(new_n680), .B(new_n683), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g483(.A1(new_n300), .A2(new_n309), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(G15gat), .B1(new_n672), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n512), .A2(new_n508), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n672), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(G15gat), .B2(new_n689), .ZN(G1326gat));
  NAND2_X1  g489(.A1(new_n672), .A2(new_n402), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  NAND4_X1  g492(.A1(new_n557), .A2(new_n640), .A3(new_n668), .A4(new_n652), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(G29gat), .A3(new_n673), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT45), .Z(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n513), .A2(new_n556), .ZN(new_n698));
  INV_X1    g497(.A(new_n441), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n490), .A2(new_n494), .A3(new_n497), .ZN(new_n700));
  INV_X1    g499(.A(new_n498), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n501), .B1(new_n477), .B2(new_n489), .ZN(new_n702));
  INV_X1    g501(.A(new_n502), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n504), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  AOI22_X1  g503(.A1(new_n699), .A2(new_n700), .B1(new_n704), .B2(KEYINPUT35), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n652), .B(new_n697), .C1(new_n698), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT108), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n652), .B1(new_n698), .B2(new_n705), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT44), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n557), .A2(new_n710), .A3(new_n652), .A4(new_n697), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n707), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n639), .B(KEYINPUT106), .Z(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n668), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n714), .A2(new_n599), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n712), .A2(new_n674), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G29gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n696), .A2(new_n718), .ZN(G1328gat));
  INV_X1    g518(.A(new_n495), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n694), .A2(G36gat), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT46), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n712), .A2(new_n495), .A3(new_n716), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G36gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1329gat));
  NAND3_X1  g524(.A1(new_n712), .A2(new_n688), .A3(new_n716), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G43gat), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n685), .A2(G43gat), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n694), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT47), .B1(new_n731), .B2(KEYINPUT109), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n729), .B1(new_n726), .B2(G43gat), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT47), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n732), .A2(new_n736), .ZN(G1330gat));
  NAND3_X1  g536(.A1(new_n712), .A2(new_n402), .A3(new_n716), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G50gat), .ZN(new_n739));
  OR3_X1    g538(.A1(new_n694), .A2(G50gat), .A3(new_n403), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1331gat));
  AND2_X1   g542(.A1(new_n557), .A2(new_n714), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n652), .A2(new_n598), .A3(new_n668), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n673), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(new_n602), .ZN(G1332gat));
  NOR2_X1   g547(.A1(new_n746), .A2(new_n720), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  AND2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n749), .B2(new_n750), .ZN(G1333gat));
  INV_X1    g552(.A(new_n688), .ZN(new_n754));
  OAI21_X1  g553(.A(G71gat), .B1(new_n746), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n686), .A2(new_n610), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n746), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g557(.A1(new_n746), .A2(new_n403), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(new_n611), .ZN(G1335gat));
  NAND2_X1  g559(.A1(new_n599), .A2(new_n668), .ZN(new_n761));
  INV_X1    g560(.A(new_n639), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n712), .A2(new_n674), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n761), .B1(KEYINPUT111), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n557), .A2(new_n652), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n765), .A2(KEYINPUT111), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n768), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n557), .A2(new_n652), .A3(new_n770), .A4(new_n766), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n674), .A2(new_n621), .A3(new_n639), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT112), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n764), .A2(new_n621), .B1(new_n772), .B2(new_n774), .ZN(G1336gat));
  NAND3_X1  g574(.A1(new_n712), .A2(new_n495), .A3(new_n763), .ZN(new_n776));
  INV_X1    g575(.A(new_n772), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n720), .A2(new_n713), .A3(G92gat), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n776), .A2(G92gat), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1337gat));
  NAND3_X1  g580(.A1(new_n712), .A2(new_n688), .A3(new_n763), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G99gat), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n685), .A2(G99gat), .A3(new_n762), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n784), .B(KEYINPUT113), .Z(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n772), .B2(new_n785), .ZN(G1338gat));
  NAND3_X1  g585(.A1(new_n712), .A2(new_n402), .A3(new_n763), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G106gat), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n713), .A2(G106gat), .A3(new_n403), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT114), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n769), .A2(new_n771), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n769), .A2(KEYINPUT116), .A3(new_n771), .A4(new_n790), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n788), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n788), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n790), .B(KEYINPUT115), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n777), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT53), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n788), .A2(new_n796), .A3(KEYINPUT117), .A4(new_n793), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n799), .A2(new_n803), .A3(new_n804), .ZN(G1339gat));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n632), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT54), .B1(new_n629), .B2(new_n631), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n807), .B(new_n636), .C1(new_n632), .C2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n632), .A2(new_n808), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n636), .A4(new_n807), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n811), .A2(new_n598), .A3(new_n637), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n580), .A2(new_n581), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n585), .A2(new_n586), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n594), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT118), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n817), .A2(KEYINPUT118), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n639), .A2(new_n596), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT119), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n814), .A2(new_n823), .A3(new_n820), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(new_n651), .A3(new_n824), .ZN(new_n825));
  AND4_X1   g624(.A1(new_n596), .A2(new_n811), .A3(new_n818), .A4(new_n819), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n652), .A2(new_n637), .A3(new_n813), .A4(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n715), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n745), .A2(new_n762), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n685), .A2(new_n402), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n495), .A2(new_n673), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(G113gat), .B1(new_n833), .B2(new_n599), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n828), .A2(new_n829), .ZN(new_n835));
  INV_X1    g634(.A(new_n504), .ZN(new_n836));
  INV_X1    g635(.A(new_n832), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n251), .A3(new_n598), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT120), .ZN(G1340gat));
  OAI21_X1  g640(.A(G120gat), .B1(new_n833), .B2(new_n713), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n253), .A3(new_n639), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1341gat));
  OAI21_X1  g643(.A(G127gat), .B1(new_n833), .B2(new_n668), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n838), .A2(new_n250), .A3(new_n715), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT121), .ZN(G1342gat));
  INV_X1    g647(.A(G134gat), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n838), .A2(new_n849), .A3(new_n652), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n833), .B2(new_n651), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n821), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n814), .A2(KEYINPUT122), .A3(new_n820), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n651), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n715), .B1(new_n859), .B2(new_n827), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n402), .B1(new_n860), .B2(new_n829), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT57), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n837), .A2(new_n688), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n864), .B(new_n402), .C1(new_n828), .C2(new_n829), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n862), .A2(new_n598), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n855), .B1(new_n866), .B2(G141gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n402), .B1(new_n828), .B2(new_n829), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n598), .A2(new_n313), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT123), .ZN(new_n870));
  NOR4_X1   g669(.A1(new_n868), .A2(new_n688), .A3(new_n837), .A4(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n871), .B1(new_n866), .B2(G141gat), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n867), .A2(new_n872), .A3(KEYINPUT58), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  AOI221_X4 g673(.A(new_n871), .B1(new_n855), .B2(new_n874), .C1(new_n866), .C2(G141gat), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n873), .A2(new_n875), .ZN(G1344gat));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  INV_X1    g676(.A(new_n868), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT57), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n861), .A2(new_n864), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n639), .A3(new_n863), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n877), .B1(new_n882), .B2(G148gat), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n877), .B1(new_n884), .B2(new_n762), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n311), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n878), .A2(new_n863), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n639), .A2(new_n311), .ZN(new_n888));
  OAI22_X1  g687(.A1(new_n883), .A2(new_n886), .B1(new_n887), .B2(new_n888), .ZN(G1345gat));
  NOR3_X1   g688(.A1(new_n884), .A2(new_n317), .A3(new_n668), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n878), .A2(new_n715), .A3(new_n863), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n317), .B2(new_n891), .ZN(G1346gat));
  NOR3_X1   g691(.A1(new_n884), .A2(new_n318), .A3(new_n651), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n878), .A2(new_n652), .A3(new_n863), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(new_n318), .B2(new_n894), .ZN(G1347gat));
  NOR2_X1   g694(.A1(new_n720), .A2(new_n674), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n835), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n831), .ZN(new_n899));
  OAI21_X1  g698(.A(G169gat), .B1(new_n899), .B2(new_n599), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n835), .A2(new_n836), .A3(new_n897), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n221), .A3(new_n598), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1348gat));
  NOR3_X1   g702(.A1(new_n899), .A2(new_n220), .A3(new_n713), .ZN(new_n904));
  AOI21_X1  g703(.A(G176gat), .B1(new_n901), .B2(new_n639), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(G1349gat));
  NAND3_X1  g705(.A1(new_n901), .A2(new_n234), .A3(new_n715), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n907), .A2(KEYINPUT125), .ZN(new_n908));
  OAI21_X1  g707(.A(G183gat), .B1(new_n899), .B2(new_n668), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT60), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n908), .A2(new_n912), .A3(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1350gat));
  NAND3_X1  g713(.A1(new_n901), .A2(new_n228), .A3(new_n652), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n831), .A3(new_n652), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n916), .A2(new_n917), .A3(G190gat), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n916), .B2(G190gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(G1351gat));
  AOI21_X1  g719(.A(new_n897), .B1(new_n879), .B2(new_n880), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n598), .A3(new_n754), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G197gat), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n868), .A2(new_n688), .A3(new_n897), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n336), .A3(new_n598), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1352gat));
  NAND4_X1  g725(.A1(new_n881), .A2(new_n754), .A3(new_n714), .A4(new_n896), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT126), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n921), .A2(new_n929), .A3(new_n754), .A4(new_n714), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(G204gat), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n924), .A2(new_n337), .A3(new_n639), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT62), .Z(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1353gat));
  NAND4_X1  g733(.A1(new_n881), .A2(new_n754), .A3(new_n715), .A4(new_n896), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G211gat), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT63), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n924), .A2(new_n347), .A3(new_n715), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT127), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT63), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n935), .A2(new_n940), .A3(G211gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n937), .A2(new_n939), .A3(new_n941), .ZN(G1354gat));
  AOI21_X1  g741(.A(G218gat), .B1(new_n924), .B2(new_n652), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n921), .A2(new_n754), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n651), .A2(new_n348), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(G1355gat));
endmodule


