//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n202));
  XOR2_X1   g001(.A(G141gat), .B(G148gat), .Z(new_n203));
  XNOR2_X1  g002(.A(G155gat), .B(G162gat), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT2), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n204), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT77), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n203), .A2(KEYINPUT77), .A3(new_n204), .A4(new_n207), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(KEYINPUT76), .B(KEYINPUT2), .Z(new_n213));
  NAND2_X1  g012(.A1(new_n203), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n204), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n202), .B1(new_n217), .B2(KEYINPUT3), .ZN(new_n218));
  XNOR2_X1  g017(.A(G197gat), .B(G204gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT71), .B(G211gat), .ZN(new_n220));
  INV_X1    g019(.A(G218gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n219), .B1(new_n222), .B2(KEYINPUT22), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT72), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G211gat), .B(G218gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n223), .B(KEYINPUT72), .ZN(new_n228));
  INV_X1    g027(.A(new_n226), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n230), .A3(KEYINPUT73), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT73), .B1(new_n227), .B2(new_n230), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n218), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n210), .A2(new_n211), .B1(new_n215), .B2(new_n214), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n227), .A2(new_n230), .A3(new_n202), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G228gat), .ZN(new_n240));
  INV_X1    g039(.A(G233gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n234), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n230), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n244), .A2(new_n218), .ZN(new_n245));
  OAI22_X1  g044(.A1(new_n238), .A2(new_n245), .B1(new_n240), .B2(new_n241), .ZN(new_n246));
  XNOR2_X1  g045(.A(G78gat), .B(G106gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT31), .B(G50gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G22gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(KEYINPUT81), .A2(G22gat), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n251), .B1(new_n252), .B2(new_n249), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n243), .A2(new_n246), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n254), .B1(new_n243), .B2(new_n246), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT5), .ZN(new_n258));
  XNOR2_X1  g057(.A(G113gat), .B(G120gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(KEYINPUT1), .ZN(new_n260));
  XNOR2_X1  g059(.A(G127gat), .B(G134gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT69), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n261), .A2(KEYINPUT68), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT1), .B1(new_n259), .B2(KEYINPUT69), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n261), .A2(KEYINPUT68), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n263), .B(new_n264), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n235), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT78), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n235), .A2(KEYINPUT78), .A3(new_n267), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n270), .B(new_n271), .C1(new_n235), .C2(new_n267), .ZN(new_n272));
  NAND2_X1  g071(.A1(G225gat), .A2(G233gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n258), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n217), .A2(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n263), .A2(new_n264), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n265), .A2(new_n266), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(new_n235), .B2(new_n237), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n217), .A2(new_n279), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT4), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n283), .A3(new_n273), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n270), .A2(new_n271), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(KEYINPUT4), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n275), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n282), .A2(KEYINPUT4), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n288), .B1(new_n285), .B2(KEYINPUT4), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT79), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n258), .B(new_n273), .C1(new_n276), .C2(new_n280), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n290), .B1(new_n289), .B2(new_n292), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n287), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G1gat), .B(G29gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT0), .ZN(new_n298));
  XNOR2_X1  g097(.A(G57gat), .B(G85gat), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n298), .B(new_n299), .Z(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n296), .A2(KEYINPUT6), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n289), .A2(new_n292), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT79), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(new_n293), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n300), .B1(new_n306), .B2(new_n287), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n300), .B(new_n287), .C1(new_n294), .C2(new_n295), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT6), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n307), .B1(new_n310), .B2(KEYINPUT80), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n312), .A3(new_n309), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n303), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n244), .ZN(new_n315));
  INV_X1    g114(.A(G226gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(new_n241), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT26), .ZN(new_n320));
  INV_X1    g119(.A(G183gat), .ZN(new_n321));
  INV_X1    g120(.A(G190gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT26), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(new_n319), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT27), .B(G183gat), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n329), .A2(KEYINPUT28), .A3(new_n322), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT28), .B1(new_n329), .B2(new_n322), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT67), .ZN(new_n333));
  XOR2_X1   g132(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT24), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n321), .A2(G190gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n322), .A2(G183gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NOR3_X1   g138(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT24), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT65), .ZN(new_n342));
  OR3_X1    g141(.A1(new_n339), .A2(KEYINPUT65), .A3(new_n340), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n319), .A2(KEYINPUT23), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n346), .B1(G169gat), .B2(G176gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n324), .A3(new_n347), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n348), .A2(KEYINPUT66), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(KEYINPUT66), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n335), .B1(new_n344), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT25), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n341), .A2(new_n353), .A3(new_n348), .ZN(new_n354));
  OAI211_X1 g153(.A(KEYINPUT74), .B(new_n333), .C1(new_n352), .C2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n342), .B(new_n343), .C1(new_n349), .C2(new_n350), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n354), .B1(new_n357), .B2(new_n334), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT67), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n332), .B(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n356), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n318), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n317), .A2(KEYINPUT29), .ZN(new_n363));
  INV_X1    g162(.A(new_n332), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n363), .B1(new_n358), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n315), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n233), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n231), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n355), .A2(new_n361), .A3(new_n363), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n358), .A2(new_n364), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n317), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G64gat), .B(G92gat), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n374), .B(new_n375), .Z(new_n376));
  NAND3_X1  g175(.A1(new_n367), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n377), .A2(KEYINPUT30), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT30), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n367), .A2(new_n373), .A3(new_n379), .A4(new_n376), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT75), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n373), .ZN(new_n383));
  INV_X1    g182(.A(new_n376), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI211_X1 g184(.A(KEYINPUT75), .B(new_n376), .C1(new_n367), .C2(new_n373), .ZN(new_n386));
  OAI22_X1  g185(.A1(new_n378), .A2(new_n381), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n257), .B1(new_n314), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G15gat), .B(G43gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G71gat), .B(G99gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n279), .B(new_n333), .C1(new_n352), .C2(new_n354), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n267), .B1(new_n358), .B2(new_n360), .ZN(new_n393));
  INV_X1    g192(.A(G227gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(new_n241), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n391), .B1(new_n396), .B2(KEYINPUT32), .ZN(new_n397));
  INV_X1    g196(.A(new_n396), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n397), .B1(KEYINPUT33), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n391), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n400), .A2(KEYINPUT70), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(KEYINPUT70), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(KEYINPUT33), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n396), .A2(KEYINPUT32), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT34), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n392), .A2(new_n393), .ZN(new_n407));
  INV_X1    g206(.A(new_n395), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI211_X1 g208(.A(KEYINPUT34), .B(new_n395), .C1(new_n392), .C2(new_n393), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n405), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n399), .A2(new_n404), .A3(new_n411), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n413), .A2(KEYINPUT36), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT36), .B1(new_n413), .B2(new_n414), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT82), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n387), .A2(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(KEYINPUT83), .B(KEYINPUT40), .Z(new_n421));
  NAND2_X1  g220(.A1(new_n285), .A2(KEYINPUT4), .ZN(new_n422));
  INV_X1    g221(.A(new_n288), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n281), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n274), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n300), .B1(new_n425), .B2(KEYINPUT39), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n273), .B1(new_n289), .B2(new_n281), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT39), .B1(new_n272), .B2(new_n274), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n421), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n296), .A2(new_n301), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n429), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT39), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n301), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(KEYINPUT40), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT84), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n433), .A2(new_n435), .A3(KEYINPUT84), .A4(KEYINPUT40), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n432), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n377), .A2(KEYINPUT30), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n380), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n442), .B(KEYINPUT82), .C1(new_n385), .C2(new_n386), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n420), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n255), .A2(new_n256), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n383), .A2(new_n384), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n376), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n446), .A2(new_n449), .B1(KEYINPUT37), .B2(new_n383), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT38), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n355), .A2(new_n361), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n317), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n244), .A3(new_n365), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n370), .A2(new_n372), .ZN(new_n456));
  INV_X1    g255(.A(new_n369), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n454), .A2(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n453), .A2(KEYINPUT85), .A3(new_n244), .A4(new_n365), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n447), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n376), .B1(new_n367), .B2(new_n373), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n451), .B1(new_n461), .B2(new_n448), .ZN(new_n462));
  OAI22_X1  g261(.A1(new_n450), .A2(new_n451), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n302), .B(new_n377), .C1(new_n310), .C2(new_n307), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n445), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n388), .B(new_n418), .C1(new_n444), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n420), .A2(new_n443), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n310), .A2(new_n307), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(new_n303), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n445), .A2(new_n413), .A3(new_n470), .A4(new_n414), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n445), .A2(new_n413), .A3(new_n414), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n314), .A2(new_n387), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n473), .B1(new_n475), .B2(new_n470), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n466), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G232gat), .A2(G233gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT41), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT15), .ZN(new_n481));
  XNOR2_X1  g280(.A(G43gat), .B(G50gat), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n481), .B1(new_n482), .B2(KEYINPUT86), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(KEYINPUT86), .B2(new_n482), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT88), .B(G43gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n485), .A2(G50gat), .ZN(new_n486));
  INV_X1    g285(.A(G50gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n487), .A2(G43gat), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n481), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n490));
  INV_X1    g289(.A(G29gat), .ZN(new_n491));
  INV_X1    g290(.A(G36gat), .ZN(new_n492));
  OR3_X1    g291(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT87), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT87), .B1(new_n491), .B2(new_n492), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n495));
  OR3_X1    g294(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n493), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n484), .A2(new_n489), .A3(new_n490), .A4(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n484), .A2(new_n489), .A3(new_n497), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT89), .B1(new_n484), .B2(new_n497), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT7), .ZN(new_n503));
  OR2_X1    g302(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n504));
  INV_X1    g303(.A(G92gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT8), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n503), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  OR2_X1    g309(.A1(G99gat), .A2(G106gat), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n508), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n503), .A2(new_n513), .A3(new_n507), .A4(new_n509), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n480), .B1(new_n501), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT90), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n501), .A2(new_n517), .A3(KEYINPUT17), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n501), .B2(KEYINPUT17), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n501), .A2(KEYINPUT17), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n515), .B(KEYINPUT99), .Z(new_n522));
  AND2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n516), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G190gat), .B(G218gat), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n526), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(G134gat), .B(G162gat), .Z(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT97), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n479), .A2(KEYINPUT41), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(new_n527), .B2(KEYINPUT100), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT100), .A4(new_n534), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G71gat), .A2(G78gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT9), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT93), .ZN(new_n542));
  INV_X1    g341(.A(G57gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(G64gat), .ZN(new_n544));
  INV_X1    g343(.A(G64gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(G57gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n539), .A2(new_n548), .A3(new_n540), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n542), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n539), .A2(KEYINPUT92), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n539), .A2(KEYINPUT92), .ZN(new_n552));
  INV_X1    g351(.A(G71gat), .ZN(new_n553));
  INV_X1    g352(.A(G78gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n551), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT94), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n555), .A2(new_n539), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n559), .A2(new_n542), .A3(new_n547), .A4(new_n549), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n558), .B1(new_n557), .B2(new_n560), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(KEYINPUT21), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G15gat), .B(G22gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT16), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n570), .B2(G1gat), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(G1gat), .B2(new_n569), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G8gat), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(new_n565), .B2(KEYINPUT21), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n568), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT96), .ZN(new_n577));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(KEYINPUT95), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n577), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G183gat), .B(G211gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n575), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT101), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n515), .B1(new_n561), .B2(new_n563), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n512), .A2(new_n514), .A3(new_n560), .A4(new_n557), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT10), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n512), .A2(KEYINPUT10), .A3(new_n514), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n591), .B1(new_n562), .B2(new_n564), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n587), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n588), .A2(new_n589), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n595), .A2(new_n586), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G120gat), .B(G148gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT102), .ZN(new_n599));
  XOR2_X1   g398(.A(G176gat), .B(G204gat), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n597), .B(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n538), .A2(new_n584), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G113gat), .B(G141gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G197gat), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT11), .B(G169gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n607), .B(KEYINPUT12), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n573), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n610), .B(new_n521), .C1(new_n518), .C2(new_n519), .ZN(new_n611));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n501), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n573), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT18), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n609), .B1(new_n617), .B2(KEYINPUT91), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n611), .A2(KEYINPUT18), .A3(new_n612), .A4(new_n614), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n501), .B(new_n610), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n612), .B(KEYINPUT13), .Z(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g423(.A1(new_n615), .A2(new_n616), .B1(new_n620), .B2(new_n621), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT91), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n626), .B1(new_n615), .B2(new_n616), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n625), .B(new_n619), .C1(new_n627), .C2(new_n609), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n603), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n477), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n314), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G1gat), .ZN(G1324gat));
  INV_X1    g433(.A(new_n632), .ZN(new_n635));
  OAI21_X1  g434(.A(G8gat), .B1(new_n635), .B2(new_n467), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT42), .ZN(new_n637));
  INV_X1    g436(.A(new_n467), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT16), .B(G8gat), .Z(new_n639));
  NAND3_X1  g438(.A1(new_n632), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n637), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n641), .A2(KEYINPUT103), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(KEYINPUT103), .ZN(new_n643));
  OAI221_X1 g442(.A(new_n636), .B1(new_n637), .B2(new_n640), .C1(new_n642), .C2(new_n643), .ZN(G1325gat));
  NAND2_X1  g443(.A1(new_n413), .A2(new_n414), .ZN(new_n645));
  OR3_X1    g444(.A1(new_n635), .A2(G15gat), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(G15gat), .B1(new_n635), .B2(new_n418), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(G1326gat));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n257), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT104), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT43), .B(G22gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  AOI21_X1  g451(.A(new_n538), .B1(new_n466), .B2(new_n476), .ZN(new_n653));
  INV_X1    g452(.A(new_n602), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n630), .A2(new_n584), .A3(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(new_n491), .A3(new_n314), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT45), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n653), .A2(KEYINPUT44), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n653), .A2(KEYINPUT44), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n661), .A2(new_n314), .A3(new_n655), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n658), .B1(new_n662), .B2(new_n491), .ZN(G1328gat));
  NAND4_X1  g462(.A1(new_n659), .A2(new_n638), .A3(new_n660), .A4(new_n655), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(G36gat), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n656), .A2(new_n492), .A3(new_n638), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT46), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT46), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n656), .A2(new_n668), .A3(new_n492), .A4(new_n638), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT105), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n665), .A2(new_n672), .A3(new_n667), .A4(new_n669), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(G1329gat));
  NAND4_X1  g473(.A1(new_n659), .A2(new_n417), .A3(new_n660), .A4(new_n655), .ZN(new_n675));
  INV_X1    g474(.A(new_n485), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n645), .A2(new_n676), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n656), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT47), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n675), .A2(new_n676), .B1(new_n656), .B2(new_n678), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT47), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n683), .A2(KEYINPUT106), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n682), .A2(new_n685), .ZN(G1330gat));
  NAND4_X1  g485(.A1(new_n661), .A2(G50gat), .A3(new_n257), .A4(new_n655), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n656), .A2(new_n257), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n487), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n687), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n690), .B1(new_n687), .B2(new_n689), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(G1331gat));
  NAND2_X1  g492(.A1(new_n458), .A2(new_n459), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT37), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT38), .B1(new_n446), .B2(new_n449), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n383), .A2(KEYINPUT37), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n697), .B1(new_n461), .B2(new_n448), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n695), .A2(new_n696), .B1(new_n698), .B2(KEYINPUT38), .ZN(new_n699));
  INV_X1    g498(.A(new_n464), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n257), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n420), .A2(new_n440), .A3(new_n443), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n417), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n387), .ZN(new_n704));
  INV_X1    g503(.A(new_n474), .ZN(new_n705));
  INV_X1    g504(.A(new_n313), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n312), .B1(new_n308), .B2(new_n309), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n706), .A2(new_n707), .A3(new_n307), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n704), .B(new_n705), .C1(new_n708), .C2(new_n303), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT35), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n703), .A2(new_n388), .B1(new_n710), .B2(new_n473), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n630), .A2(new_n538), .A3(new_n584), .A4(new_n654), .ZN(new_n712));
  OR3_X1    g511(.A1(new_n711), .A2(KEYINPUT108), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT108), .B1(new_n711), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n314), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(new_n543), .ZN(G1332gat));
  NOR2_X1   g517(.A1(new_n715), .A2(new_n467), .ZN(new_n719));
  NOR2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  AND2_X1   g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n719), .B2(new_n720), .ZN(G1333gat));
  OAI21_X1  g522(.A(G71gat), .B1(new_n715), .B2(new_n418), .ZN(new_n724));
  INV_X1    g523(.A(new_n645), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n553), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n715), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n724), .B(KEYINPUT50), .C1(new_n715), .C2(new_n726), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(G1334gat));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n445), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(new_n554), .ZN(G1335gat));
  NOR3_X1   g532(.A1(new_n584), .A2(new_n629), .A3(new_n602), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n661), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n716), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n504), .A2(new_n506), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT109), .B1(new_n711), .B2(new_n538), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n536), .A2(new_n537), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n477), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n584), .A2(new_n629), .ZN(new_n742));
  AND4_X1   g541(.A1(KEYINPUT51), .A2(new_n738), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n742), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n653), .B2(new_n739), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT51), .B1(new_n745), .B2(new_n738), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n654), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n314), .A2(new_n737), .ZN(new_n748));
  OAI22_X1  g547(.A1(new_n736), .A2(new_n737), .B1(new_n747), .B2(new_n748), .ZN(G1336gat));
  NAND3_X1  g548(.A1(new_n638), .A2(new_n505), .A3(new_n654), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT110), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n743), .B2(new_n746), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n659), .A2(new_n638), .A3(new_n660), .A4(new_n734), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G92gat), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT52), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n753), .A2(new_n758), .A3(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(G1337gat));
  OAI21_X1  g559(.A(G99gat), .B1(new_n735), .B2(new_n418), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n743), .A2(new_n746), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n645), .A2(G99gat), .A3(new_n602), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT111), .Z(new_n764));
  OAI21_X1  g563(.A(new_n761), .B1(new_n762), .B2(new_n764), .ZN(G1338gat));
  NOR2_X1   g564(.A1(new_n445), .A2(G106gat), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n654), .B(new_n766), .C1(new_n743), .C2(new_n746), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n659), .A2(new_n257), .A3(new_n660), .A4(new_n734), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G106gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n769), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n767), .B(new_n769), .C1(new_n772), .C2(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(G1339gat));
  NOR2_X1   g575(.A1(new_n603), .A2(new_n629), .ZN(new_n777));
  OR3_X1    g576(.A1(new_n590), .A2(new_n587), .A3(new_n592), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(KEYINPUT54), .A3(new_n593), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n587), .B(new_n780), .C1(new_n590), .C2(new_n592), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n781), .A2(new_n782), .A3(new_n601), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n781), .B2(new_n601), .ZN(new_n784));
  OAI211_X1 g583(.A(KEYINPUT55), .B(new_n779), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  OR3_X1    g584(.A1(new_n594), .A2(new_n596), .A3(new_n601), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n779), .B1(new_n783), .B2(new_n784), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n625), .A2(new_n609), .A3(new_n619), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n612), .B1(new_n611), .B2(new_n614), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n620), .A2(new_n621), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n607), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n740), .A2(new_n793), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n798), .A2(new_n602), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n793), .B2(new_n629), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n802), .B2(new_n740), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n777), .B1(new_n803), .B2(new_n583), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n804), .A2(new_n716), .A3(new_n257), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(new_n725), .A3(new_n467), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n630), .ZN(new_n807));
  NAND2_X1  g606(.A1(KEYINPUT115), .A2(G113gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g608(.A(KEYINPUT115), .B(G113gat), .Z(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n807), .B2(new_n810), .ZN(G1340gat));
  NOR2_X1   g610(.A1(new_n806), .A2(new_n602), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n812), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g612(.A1(new_n806), .A2(new_n583), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n814), .B(G127gat), .Z(G1342gat));
  NAND2_X1  g614(.A1(new_n467), .A2(new_n740), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(G134gat), .A3(new_n645), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n805), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g617(.A(new_n818), .B(KEYINPUT56), .Z(new_n819));
  OAI21_X1  g618(.A(G134gat), .B1(new_n806), .B2(new_n538), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(G1343gat));
  INV_X1    g620(.A(new_n777), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n538), .A2(new_n798), .A3(new_n792), .ZN(new_n823));
  INV_X1    g622(.A(new_n801), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n630), .B2(new_n792), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n823), .B1(new_n825), .B2(new_n538), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n822), .B1(new_n826), .B2(new_n584), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n257), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n418), .A2(new_n467), .A3(new_n314), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n629), .ZN(new_n831));
  INV_X1    g630(.A(G141gat), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n829), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n445), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT55), .B1(new_n789), .B2(KEYINPUT116), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n839), .B(new_n779), .C1(new_n783), .C2(new_n784), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n787), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n629), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI211_X1 g642(.A(KEYINPUT117), .B(new_n787), .C1(new_n840), .C2(new_n838), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n824), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n538), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n584), .B1(new_n846), .B2(new_n800), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n835), .B(new_n837), .C1(new_n847), .C2(new_n777), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n836), .B1(new_n804), .B2(new_n445), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n823), .B1(new_n845), .B2(new_n538), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n822), .B1(new_n851), .B2(new_n584), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n835), .B1(new_n852), .B2(new_n837), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n834), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n630), .A2(new_n832), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n833), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT119), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT58), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n857), .A2(KEYINPUT119), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1344gat));
  NAND2_X1  g661(.A1(new_n828), .A2(KEYINPUT57), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n852), .A2(new_n836), .A3(new_n257), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n834), .A2(new_n654), .ZN(new_n866));
  OAI21_X1  g665(.A(G148gat), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT59), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n654), .B(new_n834), .C1(new_n850), .C2(new_n853), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n870));
  INV_X1    g669(.A(G148gat), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(KEYINPUT59), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n870), .B1(new_n869), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n830), .A2(new_n871), .A3(new_n654), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1345gat));
  OAI21_X1  g676(.A(G155gat), .B1(new_n854), .B2(new_n583), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n830), .A2(new_n205), .A3(new_n584), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1346gat));
  OAI21_X1  g679(.A(G162gat), .B1(new_n854), .B2(new_n538), .ZN(new_n881));
  OR4_X1    g680(.A1(G162gat), .A2(new_n816), .A3(new_n716), .A4(new_n417), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n828), .B2(new_n882), .ZN(G1347gat));
  NOR4_X1   g682(.A1(new_n804), .A2(new_n314), .A3(new_n474), .A4(new_n467), .ZN(new_n884));
  AOI21_X1  g683(.A(G169gat), .B1(new_n884), .B2(new_n629), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n804), .A2(new_n257), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n638), .A2(new_n716), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(new_n645), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT121), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n886), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n629), .A2(G169gat), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n885), .B1(new_n893), .B2(new_n894), .ZN(G1348gat));
  AOI21_X1  g694(.A(G176gat), .B1(new_n884), .B2(new_n654), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT122), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(KEYINPUT122), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n654), .A2(G176gat), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n897), .A2(new_n898), .B1(new_n893), .B2(new_n899), .ZN(G1349gat));
  NAND3_X1  g699(.A1(new_n890), .A2(new_n584), .A3(new_n892), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G183gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n329), .A3(new_n584), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n905));
  NAND2_X1  g704(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n902), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1350gat));
  NAND3_X1  g707(.A1(new_n884), .A2(new_n322), .A3(new_n740), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n890), .A2(new_n740), .A3(new_n892), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n912));
  AND4_X1   g711(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(G190gat), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n322), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n911), .A2(new_n914), .B1(new_n910), .B2(new_n912), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n909), .B1(new_n913), .B2(new_n915), .ZN(G1351gat));
  NAND3_X1  g715(.A1(new_n638), .A2(new_n257), .A3(new_n418), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT125), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n918), .A2(new_n314), .A3(new_n804), .ZN(new_n919));
  XOR2_X1   g718(.A(KEYINPUT126), .B(G197gat), .Z(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n629), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n887), .A2(new_n417), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n863), .A2(new_n864), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(new_n630), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n924), .B2(new_n920), .ZN(G1352gat));
  INV_X1    g724(.A(G204gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n919), .A2(new_n926), .A3(new_n654), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n927), .B(KEYINPUT62), .Z(new_n928));
  OAI21_X1  g727(.A(G204gat), .B1(new_n923), .B2(new_n602), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1353gat));
  NAND3_X1  g729(.A1(new_n919), .A2(new_n220), .A3(new_n584), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n923), .A2(new_n583), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n932), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT63), .B1(new_n932), .B2(G211gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(G1354gat));
  OAI21_X1  g734(.A(G218gat), .B1(new_n923), .B2(new_n538), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n221), .A3(new_n740), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1355gat));
endmodule


