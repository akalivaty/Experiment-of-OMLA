

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781;

  AND2_X2 U374 ( .A1(n433), .A2(n431), .ZN(n741) );
  NAND2_X1 U375 ( .A1(n436), .A2(n435), .ZN(n663) );
  OR2_X1 U376 ( .A1(n643), .A2(n637), .ZN(n374) );
  OR2_X1 U377 ( .A1(n767), .A2(n623), .ZN(n550) );
  XNOR2_X1 U378 ( .A(n535), .B(n352), .ZN(n351) );
  INV_X1 U379 ( .A(n527), .ZN(n352) );
  XNOR2_X1 U380 ( .A(n559), .B(n351), .ZN(n495) );
  XNOR2_X2 U381 ( .A(n606), .B(n520), .ZN(n627) );
  XNOR2_X2 U382 ( .A(n462), .B(n519), .ZN(n606) );
  INV_X1 U383 ( .A(G953), .ZN(n767) );
  NOR2_X2 U384 ( .A1(n466), .A2(n613), .ZN(n440) );
  XNOR2_X2 U385 ( .A(KEYINPUT71), .B(KEYINPUT3), .ZN(n511) );
  XNOR2_X2 U386 ( .A(n636), .B(n402), .ZN(n718) );
  XNOR2_X2 U387 ( .A(n504), .B(n503), .ZN(n751) );
  XNOR2_X2 U388 ( .A(G107), .B(G110), .ZN(n504) );
  INV_X1 U389 ( .A(n687), .ZN(n645) );
  NOR2_X2 U390 ( .A1(n781), .A2(n776), .ZN(n468) );
  NOR2_X1 U391 ( .A1(n688), .A2(n689), .ZN(n641) );
  NOR2_X1 U392 ( .A1(n689), .A2(n605), .ZN(n644) );
  XNOR2_X1 U393 ( .A(n485), .B(KEYINPUT109), .ZN(n701) );
  NAND2_X2 U394 ( .A1(n379), .A2(n376), .ZN(n687) );
  XOR2_X2 U395 ( .A(KEYINPUT4), .B(KEYINPUT68), .Z(n527) );
  XOR2_X1 U396 ( .A(G125), .B(G146), .Z(n535) );
  XNOR2_X1 U397 ( .A(n434), .B(KEYINPUT72), .ZN(n413) );
  AND2_X1 U398 ( .A1(n390), .A2(n616), .ZN(n678) );
  XNOR2_X2 U399 ( .A(n609), .B(KEYINPUT107), .ZN(n614) );
  NAND2_X1 U400 ( .A1(n373), .A2(n372), .ZN(n353) );
  NAND2_X1 U401 ( .A1(n373), .A2(n372), .ZN(n371) );
  XNOR2_X1 U402 ( .A(n353), .B(n442), .ZN(n354) );
  XNOR2_X1 U403 ( .A(n371), .B(n442), .ZN(n777) );
  XNOR2_X1 U404 ( .A(n414), .B(KEYINPUT93), .ZN(n643) );
  XNOR2_X1 U405 ( .A(n517), .B(n516), .ZN(n593) );
  NOR2_X2 U406 ( .A1(n627), .A2(n626), .ZN(n629) );
  NOR2_X2 U407 ( .A1(n414), .A2(n465), .ZN(n404) );
  XNOR2_X2 U408 ( .A(n438), .B(n437), .ZN(n779) );
  XNOR2_X1 U409 ( .A(n619), .B(n486), .ZN(n704) );
  XNOR2_X1 U410 ( .A(KEYINPUT73), .B(KEYINPUT38), .ZN(n486) );
  OR2_X1 U411 ( .A1(n648), .A2(n450), .ZN(n689) );
  XNOR2_X1 U412 ( .A(n446), .B(G131), .ZN(n760) );
  INV_X1 U413 ( .A(G140), .ZN(n446) );
  OR2_X1 U414 ( .A1(G902), .A2(G237), .ZN(n518) );
  AND2_X1 U415 ( .A1(n592), .A2(n355), .ZN(n470) );
  XNOR2_X1 U416 ( .A(n563), .B(n564), .ZN(n605) );
  XNOR2_X1 U417 ( .A(n451), .B(n764), .ZN(n742) );
  XNOR2_X1 U418 ( .A(n541), .B(n452), .ZN(n451) );
  XNOR2_X1 U419 ( .A(n453), .B(n539), .ZN(n452) );
  XNOR2_X1 U420 ( .A(n762), .B(G146), .ZN(n561) );
  AND2_X1 U421 ( .A1(n641), .A2(n635), .ZN(n636) );
  XNOR2_X1 U422 ( .A(n687), .B(n382), .ZN(n630) );
  INV_X1 U423 ( .A(KEYINPUT6), .ZN(n382) );
  NOR2_X1 U424 ( .A1(n678), .A2(n357), .ZN(n469) );
  NAND2_X1 U425 ( .A1(n439), .A2(n474), .ZN(n477) );
  AND2_X1 U426 ( .A1(n651), .A2(n640), .ZN(n474) );
  XNOR2_X1 U427 ( .A(KEYINPUT75), .B(KEYINPUT18), .ZN(n508) );
  XNOR2_X1 U428 ( .A(n515), .B(KEYINPUT76), .ZN(n516) );
  NOR2_X1 U429 ( .A1(G900), .A2(n551), .ZN(n552) );
  XNOR2_X1 U430 ( .A(n574), .B(n384), .ZN(n735) );
  XNOR2_X1 U431 ( .A(n386), .B(n385), .ZN(n384) );
  XNOR2_X1 U432 ( .A(n760), .B(n573), .ZN(n385) );
  INV_X1 U433 ( .A(n443), .ZN(n432) );
  XNOR2_X1 U434 ( .A(n598), .B(KEYINPUT39), .ZN(n599) );
  INV_X1 U435 ( .A(KEYINPUT111), .ZN(n395) );
  INV_X1 U436 ( .A(n610), .ZN(n393) );
  NOR2_X1 U437 ( .A1(n401), .A2(n634), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n546), .B(n545), .ZN(n648) );
  XNOR2_X1 U439 ( .A(n544), .B(n543), .ZN(n545) );
  INV_X1 U440 ( .A(KEYINPUT25), .ZN(n543) );
  AND2_X1 U441 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U442 ( .A1(n383), .A2(G902), .ZN(n380) );
  INV_X1 U443 ( .A(KEYINPUT22), .ZN(n403) );
  NAND2_X1 U444 ( .A1(n702), .A2(n684), .ZN(n465) );
  XNOR2_X1 U445 ( .A(n605), .B(KEYINPUT1), .ZN(n688) );
  INV_X1 U446 ( .A(n742), .ZN(n428) );
  XNOR2_X1 U447 ( .A(n445), .B(n444), .ZN(n560) );
  INV_X1 U448 ( .A(KEYINPUT44), .ZN(n464) );
  NOR2_X1 U449 ( .A1(G953), .A2(G237), .ZN(n571) );
  XOR2_X1 U450 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n570) );
  XNOR2_X1 U451 ( .A(G113), .B(G122), .ZN(n569) );
  XOR2_X1 U452 ( .A(G137), .B(KEYINPUT5), .Z(n524) );
  XOR2_X1 U453 ( .A(KEYINPUT74), .B(G131), .Z(n522) );
  XNOR2_X1 U454 ( .A(n492), .B(n491), .ZN(n514) );
  XNOR2_X1 U455 ( .A(KEYINPUT88), .B(G113), .ZN(n491) );
  XNOR2_X1 U456 ( .A(n511), .B(n512), .ZN(n492) );
  INV_X1 U457 ( .A(G119), .ZN(n512) );
  INV_X1 U458 ( .A(KEYINPUT16), .ZN(n513) );
  XNOR2_X1 U459 ( .A(n538), .B(n537), .ZN(n453) );
  XNOR2_X1 U460 ( .A(G119), .B(G140), .ZN(n537) );
  XNOR2_X1 U461 ( .A(n568), .B(n557), .ZN(n764) );
  XOR2_X1 U462 ( .A(KEYINPUT11), .B(KEYINPUT98), .Z(n573) );
  XNOR2_X1 U463 ( .A(n389), .B(n387), .ZN(n386) );
  XNOR2_X1 U464 ( .A(n569), .B(n388), .ZN(n387) );
  XNOR2_X1 U465 ( .A(n570), .B(n572), .ZN(n389) );
  INV_X1 U466 ( .A(G143), .ZN(n388) );
  XNOR2_X1 U467 ( .A(n535), .B(KEYINPUT10), .ZN(n568) );
  XOR2_X1 U468 ( .A(KEYINPUT69), .B(G137), .Z(n557) );
  NAND2_X1 U469 ( .A1(n704), .A2(n703), .ZN(n485) );
  XNOR2_X1 U470 ( .A(n586), .B(n441), .ZN(n600) );
  XNOR2_X1 U471 ( .A(n587), .B(G478), .ZN(n441) );
  NAND2_X1 U472 ( .A1(G472), .A2(n378), .ZN(n377) );
  INV_X1 U473 ( .A(G902), .ZN(n378) );
  INV_X1 U474 ( .A(n477), .ZN(n482) );
  INV_X1 U475 ( .A(G104), .ZN(n503) );
  XOR2_X1 U476 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n578) );
  XNOR2_X1 U477 ( .A(G107), .B(KEYINPUT100), .ZN(n577) );
  XNOR2_X1 U478 ( .A(n370), .B(G134), .ZN(n580) );
  XNOR2_X1 U479 ( .A(n760), .B(n558), .ZN(n445) );
  INV_X1 U480 ( .A(n557), .ZN(n444) );
  XNOR2_X1 U481 ( .A(n507), .B(n510), .ZN(n494) );
  XNOR2_X1 U482 ( .A(n461), .B(n547), .ZN(n548) );
  NAND2_X1 U483 ( .A1(G237), .A2(G234), .ZN(n547) );
  XNOR2_X1 U484 ( .A(KEYINPUT14), .B(KEYINPUT90), .ZN(n461) );
  NAND2_X1 U485 ( .A1(G214), .A2(n518), .ZN(n703) );
  INV_X1 U486 ( .A(KEYINPUT19), .ZN(n520) );
  OR2_X1 U487 ( .A1(n553), .A2(n625), .ZN(n460) );
  XNOR2_X1 U488 ( .A(n644), .B(KEYINPUT108), .ZN(n592) );
  XNOR2_X1 U489 ( .A(n575), .B(n576), .ZN(n601) );
  XNOR2_X1 U490 ( .A(n483), .B(n604), .ZN(n776) );
  XNOR2_X1 U491 ( .A(n448), .B(n447), .ZN(n781) );
  INV_X1 U492 ( .A(KEYINPUT40), .ZN(n447) );
  XNOR2_X1 U493 ( .A(n392), .B(n391), .ZN(n390) );
  INV_X1 U494 ( .A(KEYINPUT36), .ZN(n391) );
  INV_X1 U495 ( .A(KEYINPUT35), .ZN(n442) );
  INV_X1 U496 ( .A(KEYINPUT32), .ZN(n437) );
  NAND2_X1 U497 ( .A1(n630), .A2(n631), .ZN(n454) );
  INV_X1 U498 ( .A(n673), .ZN(n670) );
  BUF_X1 U499 ( .A(G110), .Z(n406) );
  NOR2_X1 U500 ( .A1(n632), .A2(n645), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n397), .B(n396), .ZN(n673) );
  INV_X1 U502 ( .A(KEYINPUT103), .ZN(n396) );
  NAND2_X1 U503 ( .A1(n601), .A2(n588), .ZN(n397) );
  XNOR2_X1 U504 ( .A(n471), .B(KEYINPUT96), .ZN(n659) );
  AND2_X1 U505 ( .A1(n644), .A2(n687), .ZN(n472) );
  AND2_X1 U506 ( .A1(n398), .A2(n360), .ZN(n657) );
  XNOR2_X1 U507 ( .A(n399), .B(KEYINPUT82), .ZN(n398) );
  INV_X1 U508 ( .A(KEYINPUT122), .ZN(n422) );
  XNOR2_X1 U509 ( .A(n739), .B(n740), .ZN(n415) );
  INV_X1 U510 ( .A(KEYINPUT60), .ZN(n420) );
  XNOR2_X1 U511 ( .A(n732), .B(n733), .ZN(n416) );
  INV_X1 U512 ( .A(KEYINPUT56), .ZN(n417) );
  AND2_X1 U513 ( .A1(n704), .A2(n554), .ZN(n355) );
  INV_X1 U514 ( .A(n684), .ZN(n450) );
  XOR2_X1 U515 ( .A(KEYINPUT30), .B(n590), .Z(n356) );
  XNOR2_X1 U516 ( .A(n460), .B(KEYINPUT77), .ZN(n591) );
  XNOR2_X1 U517 ( .A(KEYINPUT15), .B(G902), .ZN(n531) );
  AND2_X1 U518 ( .A1(n671), .A2(n612), .ZN(n357) );
  INV_X1 U519 ( .A(n648), .ZN(n683) );
  XNOR2_X1 U520 ( .A(G122), .B(G116), .ZN(n359) );
  AND2_X1 U521 ( .A1(n688), .A2(n683), .ZN(n360) );
  INV_X1 U522 ( .A(n630), .ZN(n635) );
  INV_X1 U523 ( .A(G472), .ZN(n383) );
  AND2_X1 U524 ( .A1(n663), .A2(n464), .ZN(n361) );
  AND2_X1 U525 ( .A1(n592), .A2(n554), .ZN(n362) );
  AND2_X1 U526 ( .A1(n620), .A2(n681), .ZN(n363) );
  XNOR2_X1 U527 ( .A(n726), .B(n725), .ZN(n364) );
  XOR2_X1 U528 ( .A(n655), .B(n654), .Z(n365) );
  AND2_X1 U529 ( .A1(n652), .A2(n501), .ZN(n366) );
  XOR2_X1 U530 ( .A(n502), .B(KEYINPUT65), .Z(n367) );
  INV_X1 U531 ( .A(KEYINPUT45), .ZN(n481) );
  XOR2_X1 U532 ( .A(n735), .B(n734), .Z(n368) );
  INV_X1 U533 ( .A(KEYINPUT80), .ZN(n501) );
  INV_X1 U534 ( .A(n743), .ZN(n426) );
  XOR2_X1 U535 ( .A(KEYINPUT87), .B(KEYINPUT63), .Z(n369) );
  INV_X1 U536 ( .A(KEYINPUT2), .ZN(n653) );
  XNOR2_X1 U537 ( .A(n370), .B(n506), .ZN(n507) );
  XNOR2_X2 U538 ( .A(G128), .B(G143), .ZN(n370) );
  NAND2_X1 U539 ( .A1(n400), .A2(n643), .ZN(n372) );
  AND2_X2 U540 ( .A1(n374), .A2(n375), .ZN(n373) );
  OR2_X1 U541 ( .A1(n655), .A2(n377), .ZN(n376) );
  NAND2_X1 U542 ( .A1(n655), .A2(n383), .ZN(n381) );
  AND2_X2 U543 ( .A1(n484), .A2(n363), .ZN(n765) );
  NAND2_X1 U544 ( .A1(n394), .A2(n393), .ZN(n392) );
  XNOR2_X1 U545 ( .A(n614), .B(n395), .ZN(n394) );
  NOR2_X1 U546 ( .A1(n633), .A2(n635), .ZN(n399) );
  AND2_X1 U547 ( .A1(n718), .A2(n637), .ZN(n400) );
  NOR2_X1 U548 ( .A1(n718), .A2(n637), .ZN(n401) );
  INV_X1 U549 ( .A(KEYINPUT33), .ZN(n402) );
  XNOR2_X2 U550 ( .A(n404), .B(n403), .ZN(n633) );
  AND2_X1 U551 ( .A1(n779), .A2(n361), .ZN(n457) );
  BUF_X1 U552 ( .A(n593), .Z(n619) );
  BUF_X1 U553 ( .A(n559), .Z(n405) );
  XNOR2_X1 U554 ( .A(G128), .B(n406), .ZN(n536) );
  BUF_X1 U555 ( .A(n741), .Z(n738) );
  NOR2_X2 U556 ( .A1(n567), .A2(n566), .ZN(n671) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n754), .B(n493), .ZN(n463) );
  BUF_X1 U559 ( .A(n463), .Z(n407) );
  BUF_X1 U560 ( .A(n754), .Z(n408) );
  NAND2_X1 U561 ( .A1(n473), .A2(n751), .ZN(n411) );
  NAND2_X1 U562 ( .A1(n409), .A2(n410), .ZN(n412) );
  NAND2_X1 U563 ( .A1(n412), .A2(n411), .ZN(n559) );
  INV_X1 U564 ( .A(n473), .ZN(n409) );
  INV_X1 U565 ( .A(n751), .ZN(n410) );
  NAND2_X1 U566 ( .A1(n413), .A2(n650), .ZN(n475) );
  AND2_X1 U567 ( .A1(n413), .A2(n476), .ZN(n479) );
  XNOR2_X2 U568 ( .A(n629), .B(n628), .ZN(n414) );
  NOR2_X1 U569 ( .A1(n414), .A2(n694), .ZN(n642) );
  NOR2_X1 U570 ( .A1(n415), .A2(n743), .ZN(G63) );
  NOR2_X1 U571 ( .A1(n416), .A2(n743), .ZN(G54) );
  XNOR2_X1 U572 ( .A(n418), .B(n417), .ZN(G51) );
  NAND2_X1 U573 ( .A1(n425), .A2(n426), .ZN(n418) );
  XNOR2_X1 U574 ( .A(n419), .B(n369), .ZN(G57) );
  NAND2_X1 U575 ( .A1(n429), .A2(n426), .ZN(n419) );
  XNOR2_X1 U576 ( .A(n421), .B(n420), .ZN(G60) );
  NAND2_X1 U577 ( .A1(n424), .A2(n426), .ZN(n421) );
  XNOR2_X1 U578 ( .A(n423), .B(n422), .ZN(G66) );
  NAND2_X1 U579 ( .A1(n427), .A2(n426), .ZN(n423) );
  XNOR2_X1 U580 ( .A(n736), .B(n368), .ZN(n424) );
  XNOR2_X1 U581 ( .A(n727), .B(n364), .ZN(n425) );
  XNOR2_X1 U582 ( .A(n458), .B(n428), .ZN(n427) );
  XNOR2_X1 U583 ( .A(n656), .B(n365), .ZN(n429) );
  NOR2_X1 U584 ( .A1(n657), .A2(n430), .ZN(n650) );
  NOR2_X1 U585 ( .A1(n649), .A2(KEYINPUT64), .ZN(n430) );
  NAND2_X1 U586 ( .A1(n748), .A2(n765), .ZN(n443) );
  NAND2_X2 U587 ( .A1(n455), .A2(n478), .ZN(n748) );
  NAND2_X1 U588 ( .A1(n432), .A2(KEYINPUT2), .ZN(n431) );
  NAND2_X1 U589 ( .A1(n487), .A2(n367), .ZN(n433) );
  NAND2_X1 U590 ( .A1(n457), .A2(n777), .ZN(n434) );
  XNOR2_X1 U591 ( .A(n529), .B(n530), .ZN(n655) );
  XNOR2_X1 U592 ( .A(n449), .B(n599), .ZN(n622) );
  NAND2_X1 U593 ( .A1(n748), .A2(n366), .ZN(n489) );
  INV_X1 U594 ( .A(n633), .ZN(n436) );
  NOR2_X2 U595 ( .A1(n633), .A2(n454), .ZN(n438) );
  NAND2_X1 U596 ( .A1(n639), .A2(KEYINPUT44), .ZN(n439) );
  XNOR2_X1 U597 ( .A(n440), .B(KEYINPUT48), .ZN(n484) );
  XNOR2_X1 U598 ( .A(n443), .B(n653), .ZN(n720) );
  NAND2_X1 U599 ( .A1(n622), .A2(n670), .ZN(n448) );
  NAND2_X1 U600 ( .A1(n470), .A2(n356), .ZN(n449) );
  AND2_X2 U601 ( .A1(n459), .A2(n480), .ZN(n455) );
  NAND2_X1 U602 ( .A1(n456), .A2(n488), .ZN(n487) );
  AND2_X2 U603 ( .A1(n489), .A2(n490), .ZN(n456) );
  NAND2_X1 U604 ( .A1(n463), .A2(n531), .ZN(n517) );
  NAND2_X1 U605 ( .A1(n741), .A2(G217), .ZN(n458) );
  NAND2_X1 U606 ( .A1(n475), .A2(KEYINPUT45), .ZN(n459) );
  NAND2_X1 U607 ( .A1(n593), .A2(n703), .ZN(n462) );
  XNOR2_X1 U608 ( .A(n407), .B(KEYINPUT54), .ZN(n725) );
  NAND2_X1 U609 ( .A1(n779), .A2(n663), .ZN(n649) );
  XNOR2_X1 U610 ( .A(n580), .B(n527), .ZN(n762) );
  NAND2_X1 U611 ( .A1(n469), .A2(n467), .ZN(n466) );
  XNOR2_X1 U612 ( .A(n468), .B(KEYINPUT46), .ZN(n467) );
  NAND2_X1 U613 ( .A1(n356), .A2(n362), .ZN(n597) );
  NAND2_X1 U614 ( .A1(n659), .A2(n675), .ZN(n647) );
  NAND2_X1 U615 ( .A1(n643), .A2(n472), .ZN(n471) );
  XNOR2_X2 U616 ( .A(n505), .B(KEYINPUT67), .ZN(n473) );
  XNOR2_X1 U617 ( .A(n473), .B(G116), .ZN(n521) );
  NAND2_X1 U618 ( .A1(n477), .A2(KEYINPUT45), .ZN(n480) );
  AND2_X1 U619 ( .A1(n650), .A2(n481), .ZN(n476) );
  NAND2_X1 U620 ( .A1(n479), .A2(n482), .ZN(n478) );
  NAND2_X1 U621 ( .A1(n500), .A2(KEYINPUT80), .ZN(n488) );
  INV_X1 U622 ( .A(n514), .ZN(n528) );
  NAND2_X1 U623 ( .A1(n717), .A2(n603), .ZN(n483) );
  XNOR2_X2 U624 ( .A(n602), .B(KEYINPUT41), .ZN(n717) );
  AND2_X2 U625 ( .A1(n765), .A2(n499), .ZN(n490) );
  XNOR2_X2 U626 ( .A(n496), .B(n359), .ZN(n754) );
  NAND2_X1 U627 ( .A1(n498), .A2(n497), .ZN(n496) );
  NAND2_X1 U628 ( .A1(n528), .A2(KEYINPUT16), .ZN(n497) );
  NAND2_X1 U629 ( .A1(n514), .A2(n513), .ZN(n498) );
  INV_X1 U630 ( .A(n748), .ZN(n500) );
  NAND2_X1 U631 ( .A1(n531), .A2(KEYINPUT80), .ZN(n499) );
  XNOR2_X2 U632 ( .A(G101), .B(KEYINPUT66), .ZN(n505) );
  NOR2_X1 U633 ( .A1(G952), .A2(n767), .ZN(n743) );
  INV_X1 U634 ( .A(n682), .ZN(n620) );
  INV_X1 U635 ( .A(KEYINPUT83), .ZN(n519) );
  INV_X1 U636 ( .A(KEYINPUT34), .ZN(n637) );
  INV_X1 U637 ( .A(KEYINPUT81), .ZN(n598) );
  BUF_X1 U638 ( .A(n779), .Z(n780) );
  INV_X1 U639 ( .A(n531), .ZN(n652) );
  NAND2_X1 U640 ( .A1(n652), .A2(KEYINPUT2), .ZN(n502) );
  NAND2_X1 U641 ( .A1(G224), .A2(n767), .ZN(n506) );
  XOR2_X1 U642 ( .A(KEYINPUT89), .B(KEYINPUT17), .Z(n509) );
  XNOR2_X1 U643 ( .A(n509), .B(n508), .ZN(n510) );
  AND2_X1 U644 ( .A1(G210), .A2(n518), .ZN(n515) );
  BUF_X1 U645 ( .A(n627), .Z(n567) );
  XNOR2_X1 U646 ( .A(n522), .B(n521), .ZN(n526) );
  NAND2_X1 U647 ( .A1(n571), .A2(G210), .ZN(n523) );
  XNOR2_X1 U648 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U649 ( .A(n526), .B(n525), .Z(n530) );
  XNOR2_X1 U650 ( .A(n561), .B(n528), .ZN(n529) );
  XOR2_X1 U651 ( .A(KEYINPUT21), .B(KEYINPUT95), .Z(n534) );
  NAND2_X1 U652 ( .A1(n531), .A2(G234), .ZN(n532) );
  XNOR2_X1 U653 ( .A(n532), .B(KEYINPUT20), .ZN(n542) );
  NAND2_X1 U654 ( .A1(n542), .A2(G221), .ZN(n533) );
  XOR2_X1 U655 ( .A(n534), .B(n533), .Z(n684) );
  XNOR2_X1 U656 ( .A(n536), .B(KEYINPUT94), .ZN(n539) );
  XOR2_X1 U657 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n538) );
  NAND2_X1 U658 ( .A1(G234), .A2(n767), .ZN(n540) );
  XOR2_X1 U659 ( .A(KEYINPUT8), .B(n540), .Z(n581) );
  NAND2_X1 U660 ( .A1(G221), .A2(n581), .ZN(n541) );
  NOR2_X1 U661 ( .A1(n742), .A2(G902), .ZN(n546) );
  NAND2_X1 U662 ( .A1(n542), .A2(G217), .ZN(n544) );
  NOR2_X1 U663 ( .A1(n450), .A2(n683), .ZN(n555) );
  NAND2_X1 U664 ( .A1(G952), .A2(n548), .ZN(n716) );
  NOR2_X1 U665 ( .A1(G953), .A2(n716), .ZN(n625) );
  NAND2_X1 U666 ( .A1(n548), .A2(G902), .ZN(n549) );
  XNOR2_X1 U667 ( .A(KEYINPUT92), .B(n549), .ZN(n623) );
  XOR2_X1 U668 ( .A(KEYINPUT105), .B(n550), .Z(n551) );
  XNOR2_X1 U669 ( .A(n552), .B(KEYINPUT106), .ZN(n553) );
  INV_X1 U670 ( .A(n591), .ZN(n554) );
  NAND2_X1 U671 ( .A1(n555), .A2(n554), .ZN(n607) );
  NOR2_X1 U672 ( .A1(n687), .A2(n607), .ZN(n556) );
  XOR2_X1 U673 ( .A(n556), .B(KEYINPUT28), .Z(n565) );
  XNOR2_X1 U674 ( .A(KEYINPUT70), .B(G469), .ZN(n564) );
  NAND2_X1 U675 ( .A1(G227), .A2(n767), .ZN(n558) );
  XNOR2_X1 U676 ( .A(n405), .B(n560), .ZN(n562) );
  XNOR2_X1 U677 ( .A(n562), .B(n561), .ZN(n731) );
  NOR2_X1 U678 ( .A1(G902), .A2(n731), .ZN(n563) );
  NOR2_X1 U679 ( .A1(n565), .A2(n605), .ZN(n603) );
  INV_X1 U680 ( .A(n603), .ZN(n566) );
  XNOR2_X1 U681 ( .A(KEYINPUT13), .B(G475), .ZN(n576) );
  XOR2_X1 U682 ( .A(n568), .B(G104), .Z(n574) );
  NAND2_X1 U683 ( .A1(n571), .A2(G214), .ZN(n572) );
  NOR2_X1 U684 ( .A1(G902), .A2(n735), .ZN(n575) );
  XNOR2_X1 U685 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n587) );
  XNOR2_X1 U686 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U687 ( .A(n580), .B(n579), .ZN(n585) );
  XNOR2_X1 U688 ( .A(n359), .B(KEYINPUT99), .ZN(n583) );
  NAND2_X1 U689 ( .A1(G217), .A2(n581), .ZN(n582) );
  XNOR2_X1 U690 ( .A(n582), .B(n583), .ZN(n584) );
  XNOR2_X1 U691 ( .A(n585), .B(n584), .ZN(n737) );
  NOR2_X1 U692 ( .A1(G902), .A2(n737), .ZN(n586) );
  INV_X1 U693 ( .A(n600), .ZN(n588) );
  NOR2_X1 U694 ( .A1(n601), .A2(n588), .ZN(n664) );
  INV_X1 U695 ( .A(n664), .ZN(n676) );
  XOR2_X1 U696 ( .A(KEYINPUT104), .B(n676), .Z(n621) );
  OR2_X1 U697 ( .A1(n621), .A2(n670), .ZN(n700) );
  NAND2_X1 U698 ( .A1(n671), .A2(n700), .ZN(n589) );
  NAND2_X1 U699 ( .A1(n589), .A2(KEYINPUT47), .ZN(n595) );
  NAND2_X1 U700 ( .A1(n645), .A2(n703), .ZN(n590) );
  NAND2_X1 U701 ( .A1(n601), .A2(n600), .ZN(n634) );
  NOR2_X1 U702 ( .A1(n597), .A2(n634), .ZN(n594) );
  NAND2_X1 U703 ( .A1(n594), .A2(n619), .ZN(n669) );
  NAND2_X1 U704 ( .A1(n595), .A2(n669), .ZN(n596) );
  XNOR2_X1 U705 ( .A(n596), .B(KEYINPUT78), .ZN(n613) );
  XOR2_X1 U706 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n604) );
  NOR2_X1 U707 ( .A1(n601), .A2(n600), .ZN(n702) );
  NAND2_X1 U708 ( .A1(n701), .A2(n702), .ZN(n602) );
  BUF_X1 U709 ( .A(n606), .Z(n610) );
  NOR2_X1 U710 ( .A1(n630), .A2(n607), .ZN(n608) );
  NAND2_X1 U711 ( .A1(n608), .A2(n670), .ZN(n609) );
  XOR2_X1 U712 ( .A(KEYINPUT79), .B(n700), .Z(n646) );
  INV_X1 U713 ( .A(n646), .ZN(n611) );
  NOR2_X1 U714 ( .A1(KEYINPUT47), .A2(n611), .ZN(n612) );
  INV_X1 U715 ( .A(n688), .ZN(n616) );
  NAND2_X1 U716 ( .A1(n614), .A2(n703), .ZN(n615) );
  NOR2_X1 U717 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U718 ( .A(n617), .B(KEYINPUT43), .ZN(n618) );
  NOR2_X1 U719 ( .A1(n619), .A2(n618), .ZN(n682) );
  NAND2_X1 U720 ( .A1(n622), .A2(n621), .ZN(n681) );
  XNOR2_X1 U721 ( .A(KEYINPUT91), .B(G898), .ZN(n746) );
  NAND2_X1 U722 ( .A1(G953), .A2(n746), .ZN(n755) );
  NOR2_X1 U723 ( .A1(n623), .A2(n755), .ZN(n624) );
  NOR2_X1 U724 ( .A1(n625), .A2(n624), .ZN(n626) );
  INV_X1 U725 ( .A(KEYINPUT0), .ZN(n628) );
  NOR2_X1 U726 ( .A1(n683), .A2(n688), .ZN(n631) );
  NAND2_X1 U727 ( .A1(n648), .A2(n688), .ZN(n632) );
  NAND2_X1 U728 ( .A1(n649), .A2(KEYINPUT64), .ZN(n638) );
  NAND2_X1 U729 ( .A1(n638), .A2(n354), .ZN(n639) );
  OR2_X1 U730 ( .A1(KEYINPUT44), .A2(KEYINPUT64), .ZN(n640) );
  NAND2_X1 U731 ( .A1(n645), .A2(n641), .ZN(n694) );
  XNOR2_X1 U732 ( .A(n642), .B(KEYINPUT31), .ZN(n675) );
  NAND2_X1 U733 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U734 ( .A1(n741), .A2(G472), .ZN(n656) );
  XOR2_X1 U735 ( .A(KEYINPUT62), .B(KEYINPUT85), .Z(n654) );
  XOR2_X1 U736 ( .A(n657), .B(G101), .Z(G3) );
  NOR2_X1 U737 ( .A1(n659), .A2(n673), .ZN(n658) );
  XOR2_X1 U738 ( .A(G104), .B(n658), .Z(G6) );
  NOR2_X1 U739 ( .A1(n659), .A2(n676), .ZN(n661) );
  XNOR2_X1 U740 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n660) );
  XNOR2_X1 U741 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U742 ( .A(G107), .B(n662), .ZN(G9) );
  XNOR2_X1 U743 ( .A(n663), .B(n406), .ZN(G12) );
  XOR2_X1 U744 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n666) );
  NAND2_X1 U745 ( .A1(n671), .A2(n664), .ZN(n665) );
  XNOR2_X1 U746 ( .A(n666), .B(n665), .ZN(n668) );
  XOR2_X1 U747 ( .A(G128), .B(KEYINPUT112), .Z(n667) );
  XNOR2_X1 U748 ( .A(n668), .B(n667), .ZN(G30) );
  XNOR2_X1 U749 ( .A(G143), .B(n669), .ZN(G45) );
  NAND2_X1 U750 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U751 ( .A(n672), .B(G146), .ZN(G48) );
  NOR2_X1 U752 ( .A1(n673), .A2(n675), .ZN(n674) );
  XOR2_X1 U753 ( .A(G113), .B(n674), .Z(G15) );
  NOR2_X1 U754 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U755 ( .A(G116), .B(n677), .Z(G18) );
  XNOR2_X1 U756 ( .A(n678), .B(KEYINPUT114), .ZN(n679) );
  XNOR2_X1 U757 ( .A(n679), .B(KEYINPUT37), .ZN(n680) );
  XNOR2_X1 U758 ( .A(G125), .B(n680), .ZN(G27) );
  XNOR2_X1 U759 ( .A(G134), .B(n681), .ZN(G36) );
  XOR2_X1 U760 ( .A(G140), .B(n682), .Z(G42) );
  NOR2_X1 U761 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U762 ( .A(n685), .B(KEYINPUT49), .ZN(n686) );
  NAND2_X1 U763 ( .A1(n687), .A2(n686), .ZN(n692) );
  NAND2_X1 U764 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U765 ( .A(KEYINPUT50), .B(n690), .Z(n691) );
  NOR2_X1 U766 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U767 ( .A(KEYINPUT115), .B(n693), .ZN(n695) );
  NAND2_X1 U768 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U769 ( .A(n696), .B(KEYINPUT116), .ZN(n697) );
  XOR2_X1 U770 ( .A(KEYINPUT51), .B(n697), .Z(n698) );
  NAND2_X1 U771 ( .A1(n717), .A2(n698), .ZN(n699) );
  XNOR2_X1 U772 ( .A(n699), .B(KEYINPUT117), .ZN(n712) );
  INV_X1 U773 ( .A(n718), .ZN(n710) );
  AND2_X1 U774 ( .A1(n701), .A2(n700), .ZN(n708) );
  INV_X1 U775 ( .A(n702), .ZN(n706) );
  NOR2_X1 U776 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U777 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U778 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U779 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U781 ( .A(n713), .B(KEYINPUT118), .ZN(n714) );
  XNOR2_X1 U782 ( .A(KEYINPUT52), .B(n714), .ZN(n715) );
  NOR2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n722) );
  NAND2_X1 U784 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U786 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U787 ( .A1(n767), .A2(n723), .ZN(n724) );
  XOR2_X1 U788 ( .A(KEYINPUT53), .B(n724), .Z(G75) );
  NAND2_X1 U789 ( .A1(n741), .A2(G210), .ZN(n727) );
  XOR2_X1 U790 ( .A(KEYINPUT84), .B(KEYINPUT55), .Z(n726) );
  XOR2_X1 U791 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n729) );
  XNOR2_X1 U792 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n728) );
  XNOR2_X1 U793 ( .A(n729), .B(n728), .ZN(n730) );
  XOR2_X1 U794 ( .A(n731), .B(n730), .Z(n733) );
  NAND2_X1 U795 ( .A1(n738), .A2(G469), .ZN(n732) );
  NAND2_X1 U796 ( .A1(n741), .A2(G475), .ZN(n736) );
  XOR2_X1 U797 ( .A(KEYINPUT59), .B(KEYINPUT86), .Z(n734) );
  XOR2_X1 U798 ( .A(n737), .B(KEYINPUT121), .Z(n740) );
  NAND2_X1 U799 ( .A1(n738), .A2(G478), .ZN(n739) );
  NAND2_X1 U800 ( .A1(G953), .A2(G224), .ZN(n744) );
  XOR2_X1 U801 ( .A(KEYINPUT61), .B(n744), .Z(n745) );
  NOR2_X1 U802 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U803 ( .A(n747), .B(KEYINPUT123), .ZN(n750) );
  NAND2_X1 U804 ( .A1(n748), .A2(n767), .ZN(n749) );
  NAND2_X1 U805 ( .A1(n750), .A2(n749), .ZN(n758) );
  BUF_X1 U806 ( .A(n751), .Z(n752) );
  XOR2_X1 U807 ( .A(G101), .B(n752), .Z(n753) );
  XNOR2_X1 U808 ( .A(n408), .B(n753), .ZN(n756) );
  NAND2_X1 U809 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U810 ( .A(n758), .B(n757), .Z(n759) );
  XNOR2_X1 U811 ( .A(KEYINPUT124), .B(n759), .ZN(G69) );
  XOR2_X1 U812 ( .A(n760), .B(KEYINPUT125), .Z(n761) );
  XNOR2_X1 U813 ( .A(n762), .B(n761), .ZN(n763) );
  XOR2_X1 U814 ( .A(n764), .B(n763), .Z(n770) );
  INV_X1 U815 ( .A(n770), .ZN(n766) );
  XOR2_X1 U816 ( .A(n765), .B(n766), .Z(n768) );
  NAND2_X1 U817 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U818 ( .A(KEYINPUT126), .B(n769), .ZN(n775) );
  XOR2_X1 U819 ( .A(G227), .B(n770), .Z(n771) );
  NAND2_X1 U820 ( .A1(n771), .A2(G900), .ZN(n772) );
  NAND2_X1 U821 ( .A1(G953), .A2(n772), .ZN(n773) );
  XOR2_X1 U822 ( .A(KEYINPUT127), .B(n773), .Z(n774) );
  NAND2_X1 U823 ( .A1(n775), .A2(n774), .ZN(G72) );
  XOR2_X1 U824 ( .A(n776), .B(G137), .Z(G39) );
  INV_X1 U825 ( .A(n354), .ZN(n778) );
  XOR2_X1 U826 ( .A(G122), .B(n778), .Z(G24) );
  XNOR2_X1 U827 ( .A(n780), .B(G119), .ZN(G21) );
  XOR2_X1 U828 ( .A(n781), .B(G131), .Z(G33) );
endmodule

