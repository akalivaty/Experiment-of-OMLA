//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT66), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(G113), .A3(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT67), .B1(new_n472), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(new_n475), .A3(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G137), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n471), .A2(new_n478), .A3(new_n480), .ZN(G160));
  AND2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(new_n475), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT69), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n479), .A2(G136), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT68), .Z(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  XNOR2_X1  g069(.A(KEYINPUT3), .B(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n475), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  OAI22_X1  g074(.A1(new_n496), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(new_n475), .A3(G138), .ZN(new_n502));
  NOR3_X1   g077(.A1(new_n484), .A2(KEYINPUT70), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  AND3_X1   g079(.A1(new_n501), .A2(new_n475), .A3(G138), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n504), .B1(new_n495), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g082(.A(G138), .B(new_n475), .C1(new_n482), .C2(new_n483), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT4), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n500), .B1(new_n507), .B2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G62), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n513), .A2(new_n514), .B1(G75), .B2(G543), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n512), .A2(KEYINPUT72), .A3(G62), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n511), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT71), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(new_n521), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(G543), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n523), .A2(new_n512), .A3(new_n524), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n518), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n517), .A2(new_n528), .ZN(G166));
  INV_X1    g104(.A(new_n526), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G89), .ZN(new_n531));
  INV_X1    g106(.A(new_n525), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G51), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n535), .A2(new_n536), .B1(new_n512), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n531), .A2(new_n533), .A3(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  AOI22_X1  g115(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n511), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT73), .ZN(new_n543));
  AOI22_X1  g118(.A1(G52), .A2(new_n532), .B1(new_n530), .B2(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  AOI22_X1  g121(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n511), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n549), .A2(new_n525), .B1(new_n526), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n551), .A2(KEYINPUT74), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(KEYINPUT74), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n548), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  AOI22_X1  g135(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n511), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n563), .A2(new_n564), .B1(new_n530), .B2(G91), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n523), .A2(G53), .A3(G543), .A4(new_n524), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G299));
  OR2_X1    g143(.A1(new_n517), .A2(new_n528), .ZN(G303));
  NAND4_X1  g144(.A1(new_n523), .A2(G87), .A3(new_n512), .A4(new_n524), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n523), .A2(G49), .A3(G543), .A4(new_n524), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G288));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n575));
  AND2_X1   g150(.A1(G73), .A2(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n512), .B2(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n575), .B1(new_n577), .B2(new_n511), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OR2_X1    g154(.A1(KEYINPUT5), .A2(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(KEYINPUT5), .A2(G543), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g157(.A(KEYINPUT76), .B(G651), .C1(new_n582), .C2(new_n576), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n523), .A2(G48), .A3(G543), .A4(new_n524), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n523), .A2(G86), .A3(new_n512), .A4(new_n524), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G305));
  XOR2_X1   g164(.A(KEYINPUT78), .B(G47), .Z(new_n590));
  AOI22_X1  g165(.A1(G85), .A2(new_n530), .B1(new_n532), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n592), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n511), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT77), .Z(new_n598));
  NAND3_X1  g173(.A1(new_n594), .A2(new_n595), .A3(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n532), .A2(G54), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n512), .A2(G66), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G651), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n526), .A2(new_n607), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(KEYINPUT10), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n600), .B1(G868), .B2(new_n611), .ZN(G284));
  OAI21_X1  g187(.A(new_n600), .B1(G868), .B2(new_n611), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G299), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  INV_X1    g194(.A(new_n611), .ZN(new_n620));
  OAI21_X1  g195(.A(G868), .B1(new_n620), .B2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g197(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n623));
  XNOR2_X1  g198(.A(G323), .B(new_n623), .ZN(G282));
  NAND2_X1  g199(.A1(new_n477), .A2(new_n495), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XOR2_X1   g201(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n479), .A2(G135), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n475), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n632), .B1(new_n633), .B2(new_n634), .C1(new_n635), .C2(new_n496), .ZN(new_n636));
  INV_X1    g211(.A(G2096), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n630), .A2(new_n631), .A3(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT82), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2427), .B(G2430), .Z(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  AND3_X1   g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(G401));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(new_n629), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n637), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n672), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n670), .A2(KEYINPUT84), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  NOR3_X1   g253(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT20), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT85), .ZN(new_n682));
  XOR2_X1   g257(.A(G1981), .B(G1986), .Z(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n682), .B(new_n687), .ZN(G229));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G23), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n572), .A2(new_n573), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT33), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT86), .B(G16), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n696), .A2(G22), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G166), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1971), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n699), .A2(KEYINPUT89), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(KEYINPUT89), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n689), .A2(G6), .ZN(new_n702));
  INV_X1    g277(.A(G305), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n689), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT32), .B(G1981), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT88), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n694), .A2(new_n700), .A3(new_n701), .A4(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT87), .B(KEYINPUT34), .Z(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n479), .A2(G131), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n475), .A2(G107), .ZN(new_n713));
  OAI21_X1  g288(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n714));
  INV_X1    g289(.A(G119), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n712), .B1(new_n713), .B2(new_n714), .C1(new_n715), .C2(new_n496), .ZN(new_n716));
  MUX2_X1   g291(.A(G25), .B(new_n716), .S(G29), .Z(new_n717));
  XOR2_X1   g292(.A(KEYINPUT35), .B(G1991), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G24), .B(G290), .S(new_n696), .Z(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G1986), .Z(new_n721));
  NAND4_X1  g296(.A1(new_n710), .A2(new_n711), .A3(new_n719), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT36), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G35), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G162), .B2(new_n724), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G2090), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n695), .A2(G20), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT23), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n615), .B2(new_n689), .ZN(new_n731));
  INV_X1    g306(.A(G1956), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n728), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT96), .ZN(new_n735));
  NAND2_X1  g310(.A1(G160), .A2(G29), .ZN(new_n736));
  INV_X1    g311(.A(G34), .ZN(new_n737));
  AOI21_X1  g312(.A(G29), .B1(new_n737), .B2(KEYINPUT24), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(KEYINPUT24), .B2(new_n737), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G2084), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n689), .A2(G5), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G171), .B2(new_n689), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n742), .B1(new_n744), .B2(G1961), .ZN(new_n745));
  AOI22_X1  g320(.A1(G141), .A2(new_n479), .B1(new_n477), .B2(G105), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n485), .A2(G129), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT26), .Z(new_n749));
  NAND3_X1  g324(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT92), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  MUX2_X1   g327(.A(G32), .B(new_n752), .S(G29), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT93), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT27), .B(G1996), .Z(new_n755));
  AOI21_X1  g330(.A(new_n745), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT95), .Z(new_n757));
  OAI22_X1  g332(.A1(new_n727), .A2(G2090), .B1(new_n755), .B2(new_n754), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n724), .A2(G33), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n479), .A2(G139), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT90), .Z(new_n761));
  NAND3_X1  g336(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT25), .Z(new_n763));
  AOI22_X1  g338(.A1(new_n495), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n761), .B(new_n763), .C1(new_n475), .C2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n759), .B1(new_n765), .B2(G29), .ZN(new_n766));
  INV_X1    g341(.A(G2072), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT91), .Z(new_n769));
  NOR2_X1   g344(.A1(new_n696), .A2(G19), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n555), .B2(new_n696), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G1341), .Z(new_n772));
  NOR2_X1   g347(.A1(G4), .A2(G16), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n611), .B2(G16), .ZN(new_n774));
  INV_X1    g349(.A(G1348), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n769), .A2(new_n772), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(G168), .A2(G16), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n778), .B(KEYINPUT94), .C1(G16), .C2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(KEYINPUT94), .B2(new_n778), .ZN(new_n780));
  INV_X1    g355(.A(G1966), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G164), .A2(new_n724), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G27), .B2(new_n724), .ZN(new_n784));
  INV_X1    g359(.A(G2078), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  AOI211_X1 g362(.A(new_n786), .B(new_n787), .C1(new_n767), .C2(new_n766), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT31), .B(G11), .Z(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT30), .B(G28), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n789), .B1(new_n724), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n636), .B2(new_n724), .ZN(new_n792));
  INV_X1    g367(.A(G2067), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n724), .A2(G26), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT28), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n479), .A2(G140), .ZN(new_n796));
  OR2_X1    g371(.A1(G104), .A2(G2105), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n797), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n798));
  INV_X1    g373(.A(G128), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n796), .B(new_n798), .C1(new_n799), .C2(new_n496), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n795), .B1(new_n800), .B2(G29), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n792), .B1(new_n793), .B2(new_n801), .ZN(new_n802));
  OAI221_X1 g377(.A(new_n802), .B1(new_n793), .B2(new_n801), .C1(new_n741), .C2(new_n740), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G1961), .B2(new_n744), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n782), .A2(new_n788), .A3(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n758), .A2(new_n777), .A3(new_n805), .ZN(new_n806));
  AND3_X1   g381(.A1(new_n735), .A2(new_n757), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n723), .A2(new_n807), .ZN(G150));
  INV_X1    g383(.A(G150), .ZN(G311));
  AND2_X1   g384(.A1(new_n530), .A2(G93), .ZN(new_n810));
  INV_X1    g385(.A(G55), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n525), .A2(new_n811), .B1(new_n812), .B2(new_n511), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G860), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT37), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n611), .A2(G559), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT97), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  INV_X1    g395(.A(new_n814), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n554), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n814), .B(new_n548), .C1(new_n552), .C2(new_n553), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n820), .B(new_n824), .Z(new_n825));
  AND2_X1   g400(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n815), .B1(new_n825), .B2(KEYINPUT39), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n817), .B1(new_n826), .B2(new_n827), .ZN(G145));
  XNOR2_X1  g403(.A(new_n765), .B(new_n800), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n626), .B(new_n716), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n752), .B(G164), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n479), .A2(G142), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT98), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  INV_X1    g410(.A(G118), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n835), .A2(KEYINPUT99), .B1(new_n836), .B2(G2105), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(KEYINPUT99), .B2(new_n835), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n485), .A2(G130), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n834), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n832), .B(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n831), .B(new_n841), .Z(new_n842));
  XOR2_X1   g417(.A(G160), .B(new_n636), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n493), .B(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(G37), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n844), .B2(new_n842), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(G395));
  NOR2_X1   g423(.A1(new_n620), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n824), .B(new_n849), .ZN(new_n850));
  OR3_X1    g425(.A1(new_n611), .A2(G299), .A3(KEYINPUT101), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT101), .B1(new_n611), .B2(G299), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n611), .A2(G299), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT41), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n851), .A2(new_n856), .A3(new_n852), .A4(new_n853), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n850), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n854), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n858), .B1(new_n850), .B2(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(KEYINPUT42), .ZN(new_n861));
  NAND2_X1  g436(.A1(G290), .A2(new_n691), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n863));
  NAND2_X1  g438(.A1(G303), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(G166), .A2(KEYINPUT102), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n703), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n594), .A2(G288), .A3(new_n595), .A4(new_n598), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n864), .A2(G305), .A3(new_n865), .ZN(new_n869));
  AND4_X1   g444(.A1(new_n862), .A2(new_n867), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n867), .A2(new_n869), .B1(new_n862), .B2(new_n868), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n860), .A2(KEYINPUT42), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n861), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n872), .B1(new_n861), .B2(new_n873), .ZN(new_n875));
  OAI21_X1  g450(.A(G868), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(G868), .B2(new_n814), .ZN(G295));
  OAI21_X1  g452(.A(new_n876), .B1(G868), .B2(new_n814), .ZN(G331));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n879));
  NAND3_X1  g454(.A1(G301), .A2(new_n879), .A3(G286), .ZN(new_n880));
  NAND2_X1  g455(.A1(G286), .A2(new_n879), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n531), .A2(new_n533), .A3(KEYINPUT104), .A4(new_n538), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n881), .A2(new_n543), .A3(new_n882), .A4(new_n544), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n824), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n822), .A2(new_n880), .A3(new_n823), .A4(new_n883), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(KEYINPUT105), .A3(new_n886), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n880), .A2(new_n883), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n888), .A2(new_n889), .A3(new_n822), .A4(new_n823), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n887), .A2(new_n855), .A3(new_n890), .A4(new_n857), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n885), .A2(new_n854), .A3(new_n886), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n872), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n872), .B1(new_n891), .B2(new_n892), .ZN(new_n896));
  OR3_X1    g471(.A1(new_n895), .A2(KEYINPUT43), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n872), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n885), .A2(new_n886), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n899), .A2(new_n855), .A3(new_n857), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n859), .B1(new_n887), .B2(new_n890), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n900), .B1(new_n901), .B2(KEYINPUT106), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n903));
  AOI211_X1 g478(.A(new_n903), .B(new_n859), .C1(new_n887), .C2(new_n890), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n898), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n893), .A2(new_n894), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n908));
  OAI211_X1 g483(.A(KEYINPUT44), .B(new_n897), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT43), .B1(new_n895), .B2(new_n896), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT107), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n916));
  AOI211_X1 g491(.A(new_n916), .B(new_n913), .C1(new_n910), .C2(new_n911), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n909), .B1(new_n915), .B2(new_n917), .ZN(G397));
  OAI21_X1  g493(.A(KEYINPUT70), .B1(new_n484), .B2(new_n502), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n495), .A2(new_n505), .A3(new_n504), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n509), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n498), .A2(new_n499), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n485), .B2(G126), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G1384), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n471), .A2(G40), .A3(new_n478), .A4(new_n480), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT108), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n752), .B(G1996), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n800), .B(new_n793), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n716), .B(new_n718), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(G290), .B(G1986), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n931), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n928), .B1(new_n926), .B2(KEYINPUT50), .ZN(new_n940));
  AOI21_X1  g515(.A(G1384), .B1(new_n921), .B2(new_n923), .ZN(new_n941));
  XOR2_X1   g516(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n942));
  AND3_X1   g517(.A1(new_n941), .A2(KEYINPUT111), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT111), .B1(new_n941), .B2(new_n942), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n940), .B(new_n741), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT117), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n941), .A2(new_n946), .A3(KEYINPUT45), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n929), .B1(new_n941), .B2(KEYINPUT45), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n946), .B1(new_n941), .B2(KEYINPUT45), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OAI211_X1 g526(.A(G168), .B(new_n945), .C1(new_n951), .C2(G1966), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(G8), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n928), .B1(new_n926), .B2(new_n927), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n924), .A2(KEYINPUT45), .A3(new_n925), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT117), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n956), .A3(new_n947), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n781), .ZN(new_n958));
  AOI21_X1  g533(.A(G168), .B1(new_n958), .B2(new_n945), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT51), .B1(new_n953), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n952), .A2(new_n961), .A3(G8), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT121), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n960), .B2(new_n962), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n967));
  INV_X1    g542(.A(G1961), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n926), .A2(new_n927), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n969), .A2(new_n785), .A3(new_n929), .A4(new_n955), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n967), .A2(new_n968), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT124), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT123), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n928), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n928), .A2(new_n974), .ZN(new_n976));
  OAI22_X1  g551(.A1(new_n975), .A2(new_n976), .B1(KEYINPUT45), .B2(new_n941), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n971), .A2(G2078), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n955), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n973), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n928), .B(new_n974), .ZN(new_n981));
  INV_X1    g556(.A(new_n978), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n941), .B2(KEYINPUT45), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n981), .A2(new_n969), .A3(new_n983), .A4(KEYINPUT124), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(G301), .B1(new_n972), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT126), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT54), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI211_X1 g563(.A(KEYINPUT126), .B(G301), .C1(new_n972), .C2(new_n985), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI211_X1 g565(.A(new_n927), .B(G1384), .C1(new_n921), .C2(new_n923), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n949), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT53), .B1(new_n992), .B2(new_n785), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT122), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n924), .A2(new_n925), .A3(new_n942), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n941), .A2(KEYINPUT111), .A3(new_n942), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(G1961), .B1(new_n999), .B2(new_n940), .ZN(new_n1000));
  AND4_X1   g575(.A1(new_n954), .A2(new_n956), .A3(new_n947), .A4(new_n978), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n994), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n954), .A2(new_n956), .A3(new_n947), .A4(new_n978), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n929), .B1(new_n941), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n997), .B2(new_n998), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1003), .B(KEYINPUT122), .C1(new_n1006), .C2(G1961), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n993), .B1(new_n1002), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(G301), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n972), .A2(G301), .A3(new_n985), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n1008), .B2(G301), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n990), .A2(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1971), .B1(new_n954), .B2(new_n955), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n929), .B1(new_n941), .B2(new_n942), .ZN(new_n1016));
  AOI211_X1 g591(.A(KEYINPUT50), .B(G1384), .C1(new_n921), .C2(new_n923), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT112), .B(G2090), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(G8), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1022));
  NAND3_X1  g597(.A1(G303), .A2(G8), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G166), .A2(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1014), .B1(new_n1021), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1971), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n949), .B2(new_n991), .ZN(new_n1031));
  INV_X1    g606(.A(new_n942), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(G164), .B2(G1384), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n941), .A2(new_n1004), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1033), .A2(new_n929), .A3(new_n1034), .A4(new_n1018), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1024), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1036), .A2(KEYINPUT116), .A3(new_n1027), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1029), .A2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n940), .B(new_n1018), .C1(new_n943), .C2(new_n944), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT109), .B(new_n1030), .C1(new_n949), .C2(new_n991), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n954), .A2(new_n955), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT109), .B1(new_n1042), .B2(new_n1030), .ZN(new_n1043));
  OAI211_X1 g618(.A(G8), .B(new_n1027), .C1(new_n1041), .C2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n941), .A2(new_n929), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n573), .A2(new_n570), .A3(G1976), .A4(new_n571), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT114), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n572), .A2(new_n1048), .A3(G1976), .A4(new_n573), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1045), .A2(G8), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT52), .ZN(new_n1051));
  INV_X1    g626(.A(G1976), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(G288), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1024), .B1(new_n941), .B2(new_n929), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT49), .ZN(new_n1057));
  INV_X1    g632(.A(G1981), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n584), .A2(new_n588), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n584), .B2(new_n588), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT115), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1063), .B(new_n1057), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1054), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1066), .B1(new_n1067), .B2(KEYINPUT49), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1056), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1044), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT125), .B1(new_n1038), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1021), .A2(new_n1014), .A3(new_n1028), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n1036), .B2(new_n1027), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT125), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1044), .A4(new_n1069), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n966), .A2(new_n1013), .A3(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT56), .B(G2072), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n992), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n565), .A2(new_n1081), .A3(new_n567), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n565), .B2(new_n567), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n732), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1080), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1084), .B1(new_n1080), .B2(new_n1085), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT61), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1084), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT61), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1080), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1042), .A2(G1996), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1045), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT58), .B(G1341), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n555), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT59), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1101), .B(new_n555), .C1(new_n1095), .C2(new_n1098), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1088), .A2(new_n1094), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1096), .A2(new_n793), .ZN(new_n1104));
  OAI211_X1 g679(.A(KEYINPUT60), .B(new_n1104), .C1(new_n1006), .C2(G1348), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(KEYINPUT119), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(KEYINPUT119), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n611), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(KEYINPUT119), .A3(new_n620), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n967), .A2(new_n775), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT60), .B1(new_n1111), .B2(new_n1104), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1103), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n620), .B1(new_n1111), .B2(new_n1104), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1087), .B1(new_n1114), .B2(new_n1093), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1113), .A2(KEYINPUT120), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT120), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1078), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n964), .B2(new_n965), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n960), .A2(new_n962), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(KEYINPUT62), .A3(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1008), .A2(G301), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1071), .A2(new_n1076), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1120), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1128));
  NOR2_X1   g703(.A1(G288), .A2(G1976), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1059), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1069), .ZN(new_n1131));
  OAI22_X1  g706(.A1(new_n1130), .A2(new_n1066), .B1(new_n1131), .B2(new_n1044), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1070), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT109), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1031), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1027), .B1(new_n1137), .B2(G8), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n958), .A2(new_n945), .ZN(new_n1139));
  NOR2_X1   g714(.A1(G286), .A2(new_n1024), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(KEYINPUT63), .A3(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1133), .B1(new_n1134), .B2(new_n1142), .ZN(new_n1143));
  NOR4_X1   g718(.A1(new_n1070), .A2(new_n1138), .A3(new_n1141), .A4(KEYINPUT118), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1134), .A2(new_n1074), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1132), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1127), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n939), .B1(new_n1118), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(G1996), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n931), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT46), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n931), .B1(new_n752), .B2(new_n934), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT47), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1161));
  NOR2_X1   g736(.A1(G290), .A2(G1986), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n931), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  AOI22_X1  g739(.A1(new_n937), .A2(new_n931), .B1(new_n1164), .B2(KEYINPUT48), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1164), .A2(KEYINPUT48), .ZN(new_n1166));
  INV_X1    g741(.A(new_n718), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n716), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n935), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(G2067), .B2(new_n800), .ZN(new_n1170));
  AOI22_X1  g745(.A1(new_n1165), .A2(new_n1166), .B1(new_n1170), .B2(new_n931), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1160), .A2(new_n1161), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1152), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g748(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n912), .A2(new_n846), .A3(new_n1175), .ZN(G225));
  INV_X1    g750(.A(G225), .ZN(G308));
endmodule


