//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282, new_n1283;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n210));
  INV_X1    g0010(.A(G116), .ZN(new_n211));
  INV_X1    g0011(.A(G270), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G97), .A2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n213), .B(new_n218), .C1(G58), .C2(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G1), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT1), .Z(new_n224));
  INV_X1    g0024(.A(new_n201), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR3_X1   g0027(.A1(new_n226), .A2(new_n221), .A3(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G13), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n231), .B(G250), .C1(G257), .C2(G264), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT0), .Z(new_n233));
  NOR3_X1   g0033(.A1(new_n224), .A2(new_n228), .A3(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G264), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n212), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT65), .Z(new_n238));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT2), .ZN(new_n241));
  INV_X1    g0041(.A(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n238), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(new_n211), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n227), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(KEYINPUT7), .B1(new_n257), .B2(new_n221), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n221), .A4(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(G68), .B1(new_n258), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NOR3_X1   g0067(.A1(KEYINPUT67), .A2(G20), .A3(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G159), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G58), .A2(G68), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n221), .B1(new_n225), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n265), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT16), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n261), .A2(new_n221), .A3(new_n262), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT7), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n263), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n274), .B1(new_n281), .B2(G68), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT16), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(new_n283), .A3(new_n272), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n254), .B1(new_n277), .B2(new_n284), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n220), .A2(G20), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n220), .A2(G13), .A3(G20), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n254), .A2(KEYINPUT68), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n291), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n288), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n285), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT17), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n220), .B1(G41), .B2(G45), .ZN(new_n297));
  INV_X1    g0097(.A(G274), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n261), .A2(new_n262), .ZN(new_n300));
  INV_X1    g0100(.A(G1698), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(G223), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G87), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(G1698), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n302), .B1(new_n260), .B2(new_n303), .C1(new_n304), .C2(new_n242), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n299), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G41), .ZN(new_n308));
  OAI211_X1 g0108(.A(G1), .B(G13), .C1(new_n260), .C2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n309), .A2(new_n297), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G232), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G200), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n307), .A2(G190), .A3(new_n311), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n295), .A2(new_n296), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n283), .B1(new_n282), .B2(new_n272), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n216), .B1(new_n280), .B2(new_n263), .ZN(new_n317));
  NOR4_X1   g0117(.A1(new_n317), .A2(new_n271), .A3(KEYINPUT16), .A4(new_n274), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n253), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n292), .ZN(new_n320));
  INV_X1    g0120(.A(new_n294), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .A4(new_n314), .ZN(new_n322));
  INV_X1    g0122(.A(new_n313), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT17), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n315), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(G169), .B1(new_n307), .B2(new_n311), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n277), .A2(new_n284), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n292), .B1(new_n327), .B2(new_n253), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n326), .B1(new_n328), .B2(new_n321), .ZN(new_n329));
  INV_X1    g0129(.A(new_n312), .ZN(new_n330));
  INV_X1    g0130(.A(G179), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT18), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n334));
  INV_X1    g0134(.A(new_n326), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT18), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n325), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n216), .A2(G20), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n221), .A2(G33), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT66), .ZN(new_n342));
  INV_X1    g0142(.A(G77), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n340), .B1(new_n269), .B2(new_n202), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  XOR2_X1   g0144(.A(KEYINPUT71), .B(KEYINPUT11), .Z(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n253), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n253), .B1(new_n220), .B2(G20), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT12), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n229), .A2(G1), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(G20), .A3(new_n216), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n347), .A2(G68), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n350), .A2(new_n348), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n345), .B1(new_n344), .B2(new_n253), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT13), .ZN(new_n356));
  OAI211_X1 g0156(.A(G226), .B(new_n301), .C1(new_n255), .C2(new_n256), .ZN(new_n357));
  OAI211_X1 g0157(.A(G232), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G97), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n306), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n310), .A2(G238), .ZN(new_n362));
  INV_X1    g0162(.A(new_n299), .ZN(new_n363));
  AND4_X1   g0163(.A1(new_n356), .A2(new_n361), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n299), .B1(new_n360), .B2(new_n306), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n356), .B1(new_n365), .B2(new_n362), .ZN(new_n366));
  OAI21_X1  g0166(.A(G169), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT14), .ZN(new_n368));
  INV_X1    g0168(.A(new_n366), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n365), .A2(new_n356), .A3(new_n362), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(G179), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT14), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(G169), .C1(new_n364), .C2(new_n366), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n368), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT73), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n368), .A2(KEYINPUT73), .A3(new_n371), .A4(new_n373), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n355), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n369), .A2(G190), .A3(new_n370), .ZN(new_n379));
  OAI21_X1  g0179(.A(G200), .B1(new_n364), .B2(new_n366), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n355), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT72), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT72), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n355), .A2(new_n380), .A3(new_n383), .A4(new_n379), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n300), .A2(G222), .A3(new_n301), .ZN(new_n387));
  INV_X1    g0187(.A(G223), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n387), .B1(new_n343), .B2(new_n300), .C1(new_n304), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n306), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n310), .A2(G226), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n363), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G169), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n290), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G50), .ZN(new_n396));
  INV_X1    g0196(.A(new_n288), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n202), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n203), .A2(G20), .ZN(new_n399));
  INV_X1    g0199(.A(G150), .ZN(new_n400));
  OAI221_X1 g0200(.A(new_n399), .B1(new_n269), .B2(new_n400), .C1(new_n342), .C2(new_n291), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n253), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n396), .A2(new_n398), .A3(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n394), .B(new_n403), .C1(G179), .C2(new_n392), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n300), .A2(G232), .A3(new_n301), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n405), .B1(new_n207), .B2(new_n300), .C1(new_n304), .C2(new_n217), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n306), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n310), .A2(G244), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(new_n363), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G190), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(G200), .B2(new_n409), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G20), .A2(G77), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT15), .B(G87), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n413), .B1(new_n341), .B2(new_n414), .C1(new_n269), .C2(new_n291), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n415), .A2(new_n253), .B1(new_n343), .B2(new_n397), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n347), .A2(G77), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT69), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n418), .B(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n409), .A2(new_n393), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n407), .A2(new_n363), .A3(new_n408), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(new_n331), .B1(new_n416), .B2(new_n417), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n412), .A2(new_n420), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n392), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G190), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT9), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n403), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n396), .A2(KEYINPUT9), .A3(new_n402), .A4(new_n398), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n392), .A2(G200), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n426), .A2(new_n428), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n431), .A2(KEYINPUT10), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(KEYINPUT10), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n404), .B(new_n424), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT70), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n431), .B(KEYINPUT10), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n437), .A2(KEYINPUT70), .A3(new_n404), .A4(new_n424), .ZN(new_n438));
  AOI211_X1 g0238(.A(new_n339), .B(new_n386), .C1(new_n436), .C2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT74), .ZN(new_n440));
  NAND2_X1  g0240(.A1(KEYINPUT6), .A2(G97), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n440), .B1(new_n441), .B2(G107), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n207), .A2(KEYINPUT74), .A3(KEYINPUT6), .A4(G97), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G97), .A2(G107), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT6), .B1(new_n208), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT75), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT6), .ZN(new_n448));
  INV_X1    g0248(.A(new_n445), .ZN(new_n449));
  NOR2_X1   g0249(.A1(G97), .A2(G107), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT75), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n451), .A2(new_n452), .A3(new_n442), .A4(new_n443), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n447), .A2(G20), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n281), .A2(G107), .ZN(new_n455));
  OAI21_X1  g0255(.A(G77), .B1(new_n267), .B2(new_n268), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n253), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n220), .A2(G33), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n288), .A2(new_n459), .A3(new_n227), .A4(new_n252), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G97), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(G97), .B2(new_n397), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT76), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT76), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n461), .B(new_n464), .C1(G97), .C2(new_n397), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(G244), .B(new_n301), .C1(new_n255), .C2(new_n256), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT4), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n300), .A2(KEYINPUT4), .A3(G244), .A4(new_n301), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n300), .A2(G250), .A3(G1698), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G283), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n470), .A2(new_n471), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n306), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT5), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n308), .ZN(new_n477));
  NAND2_X1  g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n220), .A2(G45), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(G257), .A3(new_n309), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n480), .B1(new_n477), .B2(new_n478), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G274), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n475), .A2(new_n487), .A3(new_n331), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n475), .A2(new_n487), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n393), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n467), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n457), .A2(new_n253), .B1(new_n465), .B2(new_n463), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n489), .A2(G190), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n486), .B1(new_n306), .B2(new_n474), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(G200), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n492), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT77), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n491), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT19), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n221), .B1(new_n359), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n450), .A2(new_n303), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n221), .B(G68), .C1(new_n255), .C2(new_n256), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n221), .A2(G33), .A3(G97), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n499), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n253), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n460), .A2(new_n414), .ZN(new_n508));
  INV_X1    g0308(.A(new_n414), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(new_n288), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT78), .ZN(new_n513));
  OAI211_X1 g0313(.A(G238), .B(new_n301), .C1(new_n255), .C2(new_n256), .ZN(new_n514));
  OAI211_X1 g0314(.A(G244), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G116), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n306), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n306), .A2(new_n481), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(G250), .B1(G274), .B2(new_n481), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n393), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n518), .A2(new_n520), .A3(new_n331), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT78), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n507), .A2(new_n524), .A3(new_n511), .A4(new_n508), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n513), .A2(new_n522), .A3(new_n523), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n521), .A2(G200), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n500), .A2(new_n501), .B1(new_n499), .B2(new_n504), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n254), .B1(new_n528), .B2(new_n503), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n460), .A2(new_n303), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n529), .A2(new_n510), .A3(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n527), .B(new_n531), .C1(new_n410), .C2(new_n521), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT79), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n526), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n526), .A2(new_n532), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT79), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n498), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n349), .A2(G20), .A3(new_n211), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n252), .A2(new_n227), .B1(G20), .B2(new_n211), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n473), .B(new_n221), .C1(G33), .C2(new_n206), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n539), .A2(KEYINPUT20), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT20), .B1(new_n539), .B2(new_n540), .ZN(new_n542));
  OAI221_X1 g0342(.A(new_n538), .B1(new_n211), .B2(new_n460), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(G257), .B(new_n301), .C1(new_n255), .C2(new_n256), .ZN(new_n544));
  OAI211_X1 g0344(.A(G264), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n261), .A2(G303), .A3(new_n262), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n306), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n482), .A2(G270), .A3(new_n309), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n485), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n543), .A2(new_n550), .A3(G169), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT21), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(G200), .ZN(new_n554));
  INV_X1    g0354(.A(new_n543), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n554), .B(new_n555), .C1(new_n410), .C2(new_n550), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT80), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n550), .A2(KEYINPUT21), .A3(G169), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n548), .A2(G179), .A3(new_n485), .A4(new_n549), .ZN(new_n559));
  AOI211_X1 g0359(.A(new_n557), .B(new_n555), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT80), .B1(new_n561), .B2(new_n543), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n553), .B(new_n556), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n497), .B1(new_n491), .B2(new_n496), .ZN(new_n565));
  OAI211_X1 g0365(.A(G257), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n566));
  OAI211_X1 g0366(.A(G250), .B(new_n301), .C1(new_n255), .C2(new_n256), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G294), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n306), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n484), .A2(new_n306), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G264), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n572), .A3(new_n485), .ZN(new_n573));
  INV_X1    g0373(.A(G200), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT86), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT85), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n569), .A2(new_n578), .A3(new_n306), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n579), .A2(new_n485), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n570), .A2(KEYINPUT85), .B1(G264), .B2(new_n571), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n580), .A2(new_n581), .A3(new_n410), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n573), .A2(KEYINPUT86), .A3(new_n574), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n577), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n221), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  XOR2_X1   g0386(.A(KEYINPUT81), .B(KEYINPUT22), .Z(new_n587));
  INV_X1    g0387(.A(new_n341), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n586), .A2(new_n587), .B1(G116), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g0389(.A(KEYINPUT82), .B(KEYINPUT24), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n221), .A2(G107), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n592), .B(KEYINPUT23), .ZN(new_n593));
  XNOR2_X1  g0393(.A(KEYINPUT81), .B(KEYINPUT22), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n585), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n589), .A2(new_n591), .A3(new_n593), .A4(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n587), .A2(new_n221), .A3(G87), .A4(new_n300), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n588), .A2(G116), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n597), .A2(new_n593), .A3(new_n595), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n590), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(new_n600), .A3(new_n253), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n349), .A2(new_n592), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(KEYINPUT83), .A3(KEYINPUT25), .ZN(new_n603));
  OR2_X1    g0403(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n604));
  NAND2_X1  g0404(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n349), .A2(new_n592), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n603), .B(new_n606), .C1(new_n460), .C2(new_n207), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT84), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n607), .B(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n584), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n601), .A2(new_n609), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n393), .B1(new_n580), .B2(new_n581), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n573), .A2(new_n331), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n565), .A2(new_n616), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n439), .A2(new_n537), .A3(new_n564), .A4(new_n617), .ZN(G372));
  AND2_X1   g0418(.A1(new_n491), .A2(new_n496), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n531), .B1(new_n410), .B2(new_n521), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n517), .A2(KEYINPUT87), .A3(new_n306), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT87), .B1(new_n517), .B2(new_n306), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n520), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n620), .B1(G200), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n520), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT87), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n518), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n626), .B1(new_n628), .B2(new_n621), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT88), .B1(new_n629), .B2(G169), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT88), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n624), .A2(new_n631), .A3(new_n393), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n513), .A2(new_n523), .A3(new_n525), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n625), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n561), .A2(new_n543), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n613), .A2(new_n614), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n553), .B(new_n636), .C1(new_n637), .C2(new_n610), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n619), .A2(new_n635), .A3(new_n638), .A4(new_n611), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n488), .B1(G169), .B2(new_n494), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n492), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n536), .A2(new_n534), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT26), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n633), .A2(new_n634), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT89), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n640), .B2(new_n492), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n467), .A2(KEYINPUT89), .A3(new_n488), .A4(new_n490), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n635), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n639), .A2(new_n643), .A3(new_n644), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n439), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n404), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n336), .B(new_n337), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n423), .A2(new_n421), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n378), .B1(new_n381), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n325), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n653), .B1(new_n659), .B2(new_n437), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n652), .A2(new_n660), .ZN(G369));
  NAND2_X1  g0461(.A1(new_n636), .A2(new_n553), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n349), .A2(new_n221), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT90), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(KEYINPUT90), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n665), .A2(G213), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(new_n555), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n662), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n563), .B2(new_n672), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  INV_X1    g0475(.A(new_n616), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n610), .B2(new_n671), .ZN(new_n677));
  INV_X1    g0477(.A(new_n615), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n670), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g0481(.A(new_n681), .B(KEYINPUT91), .Z(new_n682));
  OAI21_X1  g0482(.A(new_n553), .B1(new_n560), .B2(new_n562), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n683), .A2(new_n671), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n684), .A2(new_n676), .B1(new_n678), .B2(new_n671), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n682), .A2(new_n685), .ZN(G399));
  INV_X1    g0486(.A(KEYINPUT29), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n619), .A2(new_n611), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n688), .B(new_n635), .C1(new_n683), .C2(new_n678), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n635), .A2(new_n648), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT26), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n642), .A2(KEYINPUT26), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n689), .A2(new_n691), .A3(new_n644), .A4(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n687), .B1(new_n693), .B2(new_n671), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n651), .A2(new_n671), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n537), .A2(new_n617), .A3(new_n564), .A4(new_n671), .ZN(new_n698));
  INV_X1    g0498(.A(new_n559), .ZN(new_n699));
  INV_X1    g0499(.A(new_n521), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n570), .A2(new_n572), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n699), .A2(new_n494), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT30), .Z(new_n703));
  AND2_X1   g0503(.A1(new_n550), .A2(new_n331), .ZN(new_n704));
  AND4_X1   g0504(.A1(new_n489), .A2(new_n704), .A3(new_n573), .A4(new_n624), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n670), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n706), .A2(KEYINPUT31), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G330), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n697), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n220), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n231), .A2(KEYINPUT92), .A3(new_n308), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT92), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n230), .B2(G41), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n501), .A2(G116), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n717), .A2(new_n220), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n226), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n717), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n722), .B(KEYINPUT28), .Z(new_n723));
  NAND2_X1  g0523(.A1(new_n712), .A2(new_n723), .ZN(G364));
  NOR2_X1   g0524(.A1(new_n229), .A2(G20), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n220), .B1(new_n725), .B2(G45), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n717), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n675), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(G330), .B2(new_n674), .ZN(new_n730));
  INV_X1    g0530(.A(new_n728), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n227), .B1(G20), .B2(new_n393), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR4_X1   g0533(.A1(new_n221), .A2(new_n331), .A3(G190), .A4(G200), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G311), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR4_X1   g0537(.A1(new_n221), .A2(new_n331), .A3(new_n574), .A4(G190), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OR2_X1    g0539(.A1(KEYINPUT33), .A2(G317), .ZN(new_n740));
  NAND2_X1  g0540(.A1(KEYINPUT33), .A2(G317), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n221), .A2(new_n410), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(G179), .A3(new_n574), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n737), .B(new_n742), .C1(G322), .C2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n221), .A2(G190), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(new_n331), .A3(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G283), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n743), .A2(new_n331), .A3(G200), .ZN(new_n751));
  INV_X1    g0551(.A(G303), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n257), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT95), .Z(new_n754));
  NAND3_X1  g0554(.A1(new_n743), .A2(G179), .A3(G200), .ZN(new_n755));
  INV_X1    g0555(.A(G326), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n747), .A2(new_n331), .A3(new_n574), .ZN(new_n757));
  INV_X1    g0557(.A(G329), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n755), .A2(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n410), .A2(G179), .A3(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n221), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n759), .B1(G294), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n746), .A2(new_n750), .A3(new_n754), .A4(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G58), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n300), .B1(new_n765), .B2(new_n744), .C1(new_n739), .C2(new_n216), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(G77), .B2(new_n734), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n761), .A2(new_n206), .B1(new_n748), .B2(new_n207), .ZN(new_n768));
  INV_X1    g0568(.A(new_n755), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n768), .B1(G50), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n751), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G87), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n757), .A2(new_n270), .ZN(new_n773));
  XOR2_X1   g0573(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n774));
  XNOR2_X1  g0574(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n767), .A2(new_n770), .A3(new_n772), .A4(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n733), .B1(new_n764), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n247), .A2(G45), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n230), .A2(new_n300), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n778), .B(new_n779), .C1(G45), .C2(new_n226), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n231), .A2(new_n300), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT93), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G355), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n780), .B(new_n783), .C1(G116), .C2(new_n231), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n732), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n777), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n787), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n789), .B1(new_n674), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n730), .B1(new_n731), .B2(new_n791), .ZN(G396));
  NAND2_X1  g0592(.A1(new_n422), .A2(new_n331), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n793), .A2(new_n421), .A3(new_n418), .A4(new_n670), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT100), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n418), .A2(new_n670), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n424), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n651), .A2(new_n671), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT101), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n710), .B(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n799), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n695), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n803), .B(new_n805), .Z(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n731), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n732), .A2(new_n785), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n257), .B1(new_n735), .B2(new_n211), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G283), .B2(new_n738), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n745), .A2(G294), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n207), .A2(new_n751), .B1(new_n755), .B2(new_n752), .ZN(new_n813));
  INV_X1    g0613(.A(new_n757), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(G311), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n748), .A2(new_n303), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G97), .B2(new_n762), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n811), .A2(new_n812), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G137), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n739), .A2(new_n400), .B1(new_n819), .B2(new_n755), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT96), .ZN(new_n821));
  INV_X1    g0621(.A(G143), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n822), .B2(new_n744), .C1(new_n270), .C2(new_n735), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT34), .Z(new_n824));
  AOI22_X1  g0624(.A1(G58), .A2(new_n762), .B1(new_n771), .B2(G50), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n748), .A2(new_n216), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(new_n257), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n825), .B(new_n827), .C1(new_n828), .C2(new_n757), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT97), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n818), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT98), .Z(new_n832));
  OAI221_X1 g0632(.A(new_n728), .B1(G77), .B2(new_n809), .C1(new_n832), .C2(new_n733), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT99), .Z(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n786), .B2(new_n799), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n807), .A2(new_n835), .ZN(G384));
  NOR2_X1   g0636(.A1(new_n655), .A2(new_n670), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n800), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n376), .A2(new_n377), .ZN(new_n840));
  INV_X1    g0640(.A(new_n355), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n670), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n842), .A2(new_n381), .A3(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n841), .B(new_n670), .C1(new_n385), .C2(new_n840), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n839), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT103), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT38), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n328), .A2(new_n321), .A3(new_n313), .A4(new_n314), .ZN(new_n851));
  INV_X1    g0651(.A(new_n668), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n334), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n336), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT37), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT104), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n336), .A2(new_n851), .A3(new_n857), .A4(new_n853), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n854), .A2(KEYINPUT104), .A3(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n853), .B1(new_n654), .B2(new_n325), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n850), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n853), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n339), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n865), .A2(KEYINPUT38), .A3(new_n859), .A4(new_n860), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n839), .A2(KEYINPUT103), .A3(new_n846), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n849), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n654), .A2(new_n852), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n869), .A2(KEYINPUT105), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT105), .B1(new_n869), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n842), .A2(new_n670), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT39), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n855), .A2(new_n858), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT106), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT106), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n855), .A2(new_n880), .A3(new_n858), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n879), .A2(new_n865), .A3(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n877), .B(new_n866), .C1(new_n882), .C2(KEYINPUT38), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n875), .B1(new_n876), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n872), .A2(new_n873), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n439), .B1(new_n694), .B2(new_n696), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n886), .A2(new_n660), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n885), .B(new_n887), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n707), .A2(new_n708), .A3(new_n799), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n878), .A2(KEYINPUT106), .B1(new_n339), .B2(new_n864), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n890), .B2(new_n881), .ZN(new_n891));
  INV_X1    g0691(.A(new_n866), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n846), .B(new_n889), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  AND4_X1   g0693(.A1(new_n707), .A2(new_n846), .A3(new_n708), .A4(new_n799), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT40), .B1(new_n863), .B2(new_n866), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n893), .A2(KEYINPUT40), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n439), .A2(new_n709), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n896), .B(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(G330), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n888), .B(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n220), .B2(new_n725), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n273), .A2(G77), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n226), .A2(new_n903), .B1(G50), .B2(new_n216), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(G1), .A3(new_n229), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n447), .A2(new_n453), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT35), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n221), .B(new_n227), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n908), .B(G116), .C1(new_n907), .C2(new_n906), .ZN(new_n909));
  XOR2_X1   g0709(.A(KEYINPUT102), .B(KEYINPUT36), .Z(new_n910));
  XNOR2_X1  g0710(.A(new_n909), .B(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n902), .A2(new_n905), .A3(new_n911), .ZN(G367));
  INV_X1    g0712(.A(KEYINPUT108), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n683), .A2(new_n671), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n491), .B(new_n496), .C1(new_n492), .C2(new_n671), .ZN(new_n915));
  OR4_X1    g0715(.A1(KEYINPUT42), .A2(new_n914), .A3(new_n616), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n684), .A2(new_n676), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT42), .B1(new_n917), .B2(new_n915), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n641), .A2(new_n670), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT107), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n915), .A2(KEYINPUT107), .A3(new_n920), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(new_n678), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n670), .B1(new_n925), .B2(new_n491), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n913), .B1(new_n919), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n916), .A2(new_n918), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n929), .A2(new_n926), .A3(KEYINPUT108), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n671), .A2(new_n531), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n644), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n635), .A2(new_n932), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT109), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n931), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT110), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT109), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n919), .A2(new_n913), .A3(new_n927), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT108), .B1(new_n929), .B2(new_n926), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n941), .B1(new_n945), .B2(new_n936), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT109), .B1(new_n928), .B2(new_n930), .ZN(new_n947));
  INV_X1    g0747(.A(new_n936), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(KEYINPUT110), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n940), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n923), .A2(new_n924), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n682), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n954));
  OR3_X1    g0754(.A1(new_n685), .A2(new_n921), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT111), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n956), .B(KEYINPUT44), .C1(new_n685), .C2(new_n921), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n685), .A2(KEYINPUT45), .A3(new_n921), .ZN(new_n958));
  AOI21_X1  g0758(.A(KEYINPUT45), .B1(new_n685), .B2(new_n921), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n955), .B(new_n957), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n682), .B(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n677), .A2(new_n679), .A3(new_n914), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT112), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n962), .A2(new_n963), .B1(new_n676), .B2(new_n684), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n917), .A2(KEYINPUT112), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n964), .A2(new_n675), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n675), .B1(new_n964), .B2(new_n965), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n711), .B1(new_n961), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n716), .B(KEYINPUT41), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n726), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n950), .A2(new_n952), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n953), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n762), .A2(G107), .B1(new_n749), .B2(G97), .ZN(new_n974));
  INV_X1    g0774(.A(G317), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n974), .B1(new_n736), .B2(new_n755), .C1(new_n975), .C2(new_n757), .ZN(new_n976));
  INV_X1    g0776(.A(G294), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n257), .B1(new_n752), .B2(new_n744), .C1(new_n739), .C2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT46), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n771), .A2(G116), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n979), .B2(new_n980), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n976), .B(new_n982), .C1(G283), .C2(new_n734), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n734), .A2(G50), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n771), .A2(G58), .B1(new_n749), .B2(G77), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n822), .B2(new_n755), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n761), .A2(new_n216), .B1(new_n757), .B2(new_n819), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n300), .B1(new_n400), .B2(new_n744), .C1(new_n739), .C2(new_n270), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n983), .B1(new_n984), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n731), .B1(new_n992), .B2(new_n732), .ZN(new_n993));
  INV_X1    g0793(.A(new_n779), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n788), .B1(new_n231), .B2(new_n414), .C1(new_n237), .C2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n933), .A2(new_n787), .A3(new_n934), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n973), .A2(new_n997), .ZN(G387));
  NOR2_X1   g0798(.A1(new_n757), .A2(new_n756), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n762), .A2(G283), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n738), .A2(G311), .B1(new_n734), .B2(G303), .ZN(new_n1001));
  INV_X1    g0801(.A(G322), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1001), .B1(new_n975), .B2(new_n744), .C1(new_n1002), .C2(new_n755), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT48), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1000), .B1(new_n977), .B2(new_n751), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1006), .A2(KEYINPUT114), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(KEYINPUT114), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1007), .A2(new_n1008), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n257), .B1(new_n211), .B2(new_n748), .C1(new_n1009), .C2(KEYINPUT49), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n999), .B(new_n1010), .C1(KEYINPUT49), .C2(new_n1009), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n762), .A2(new_n509), .B1(new_n814), .B2(G150), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n270), .B2(new_n755), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n300), .B1(new_n202), .B2(new_n744), .C1(new_n739), .C2(new_n291), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n735), .A2(new_n216), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n751), .A2(new_n343), .B1(new_n748), .B2(new_n206), .ZN(new_n1016));
  NOR4_X1   g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n732), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n677), .A2(new_n679), .A3(new_n787), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n291), .A2(G50), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT50), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n718), .B1(new_n216), .B2(new_n343), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  AOI211_X1 g0822(.A(G45), .B(new_n1022), .C1(new_n1021), .C2(new_n1020), .ZN(new_n1023));
  INV_X1    g0823(.A(G45), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n779), .B1(new_n243), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n782), .A2(new_n719), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n231), .A2(G107), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n788), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1018), .A2(new_n728), .A3(new_n1019), .A4(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT115), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n968), .A2(new_n727), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n711), .B(new_n968), .Z(new_n1033));
  OAI211_X1 g0833(.A(new_n1031), .B(new_n1032), .C1(new_n716), .C2(new_n1033), .ZN(G393));
  AOI21_X1  g0834(.A(new_n711), .B1(new_n967), .B2(new_n966), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(new_n961), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n961), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1036), .A2(new_n717), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(G283), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n751), .A2(new_n1039), .B1(new_n748), .B2(new_n207), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n257), .B1(new_n735), .B2(new_n977), .C1(new_n739), .C2(new_n752), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(G116), .C2(new_n762), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n744), .A2(new_n736), .B1(new_n755), .B2(new_n975), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT52), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(new_n1002), .C2(new_n757), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT116), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n744), .A2(new_n270), .B1(new_n755), .B2(new_n400), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT51), .Z(new_n1048));
  NOR2_X1   g0848(.A1(new_n757), .A2(new_n822), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n816), .B1(G68), .B2(new_n771), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n343), .B2(new_n761), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n300), .B1(new_n735), .B2(new_n291), .C1(new_n739), .C2(new_n202), .ZN(new_n1052));
  NOR4_X1   g0852(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1046), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n731), .B1(new_n1054), .B2(new_n732), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n788), .B1(new_n206), .B2(new_n231), .C1(new_n250), .C2(new_n994), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n951), .A2(new_n787), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n961), .B2(new_n727), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1038), .A2(new_n1059), .ZN(G390));
  NAND2_X1  g0860(.A1(new_n693), .A2(new_n671), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n838), .B1(new_n1061), .B2(new_n804), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n846), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n866), .B1(new_n882), .B2(KEYINPUT38), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1063), .A2(new_n875), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n847), .A2(new_n875), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n876), .A2(new_n883), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n889), .A2(G330), .A3(new_n846), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1065), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n439), .A2(G330), .A3(new_n709), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n886), .A2(new_n1074), .A3(new_n660), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n707), .A2(G330), .A3(new_n708), .A4(new_n799), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n846), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1069), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n839), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1062), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n1069), .A3(new_n1078), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1075), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1073), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1071), .A2(new_n1072), .A3(new_n1083), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n717), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT117), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1073), .A2(new_n726), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n876), .A2(new_n785), .A3(new_n883), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n739), .A2(new_n819), .B1(new_n270), .B2(new_n761), .ZN(new_n1092));
  XOR2_X1   g0892(.A(KEYINPUT54), .B(G143), .Z(new_n1093));
  AOI21_X1  g0893(.A(new_n1092), .B1(new_n734), .B2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT118), .Z(new_n1095));
  NAND2_X1  g0895(.A1(new_n771), .A2(G150), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT53), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n749), .A2(G50), .B1(new_n814), .B2(G125), .ZN(new_n1098));
  INV_X1    g0898(.A(G128), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1098), .B(new_n300), .C1(new_n1099), .C2(new_n755), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1095), .B(new_n1101), .C1(new_n828), .C2(new_n744), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n772), .B(new_n257), .C1(new_n211), .C2(new_n744), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n826), .B(new_n1103), .C1(G294), .C2(new_n814), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n769), .A2(G283), .B1(new_n738), .B2(G107), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n206), .B2(new_n735), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT119), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1104), .B(new_n1107), .C1(new_n343), .C2(new_n761), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n733), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n809), .A2(new_n293), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1091), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1090), .B1(new_n728), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1089), .A2(new_n1112), .ZN(G378));
  NAND2_X1  g0913(.A1(new_n403), .A2(new_n852), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n437), .A2(new_n404), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1114), .B1(new_n437), .B2(new_n404), .ZN(new_n1117));
  OAI21_X1  g0917(.A(KEYINPUT55), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1117), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT55), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n1120), .A3(new_n1115), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1118), .A2(new_n1121), .A3(KEYINPUT56), .ZN(new_n1122));
  AOI21_X1  g0922(.A(KEYINPUT56), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n896), .B2(new_n899), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n895), .A2(new_n894), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT40), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n1064), .B2(new_n894), .ZN(new_n1129));
  OAI211_X1 g0929(.A(G330), .B(new_n1124), .C1(new_n1127), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n885), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT105), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n863), .A2(new_n866), .ZN(new_n1134));
  AOI221_X4 g0934(.A(new_n848), .B1(new_n844), .B2(new_n845), .C1(new_n800), .C2(new_n838), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT103), .B1(new_n839), .B2(new_n846), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1133), .B1(new_n1137), .B2(new_n870), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n884), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n869), .A2(KEYINPUT105), .A3(new_n871), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1141), .A2(new_n1130), .A3(new_n1126), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1132), .A2(new_n1142), .A3(KEYINPUT122), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT122), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1141), .A2(new_n1144), .A3(new_n1130), .A4(new_n1126), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT57), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1075), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n1086), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1143), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n717), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT123), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1132), .A2(new_n1142), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1086), .A2(new_n1147), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n1146), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1149), .A2(KEYINPUT123), .A3(new_n717), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1152), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1124), .A2(new_n785), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n808), .A2(new_n202), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n735), .A2(new_n819), .B1(new_n1099), .B2(new_n744), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G132), .B2(new_n738), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n769), .A2(G125), .B1(new_n771), .B2(new_n1093), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n400), .C2(new_n761), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(G33), .B1(new_n749), .B2(G159), .ZN(new_n1167));
  AOI21_X1  g0967(.A(G41), .B1(new_n814), .B2(G124), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n735), .A2(new_n414), .B1(new_n207), .B2(new_n744), .ZN(new_n1170));
  AOI211_X1 g0970(.A(G41), .B(new_n1170), .C1(G97), .C2(new_n738), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n814), .A2(G283), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G116), .A2(new_n769), .B1(new_n749), .B2(G58), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n761), .A2(new_n216), .B1(new_n751), .B2(new_n343), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1174), .A2(new_n300), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT58), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n202), .B1(new_n255), .B2(G41), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1169), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT121), .Z(new_n1180));
  AOI21_X1  g0980(.A(new_n731), .B1(new_n1180), .B2(new_n732), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1159), .A2(new_n1160), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1153), .B2(new_n727), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1158), .A2(new_n1184), .ZN(G375));
  OAI22_X1  g0985(.A1(new_n755), .A2(new_n977), .B1(new_n757), .B2(new_n752), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G97), .B2(new_n771), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n257), .B1(new_n744), .B2(new_n1039), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G116), .B2(new_n738), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n734), .A2(G107), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n762), .A2(new_n509), .B1(new_n749), .B2(G77), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1187), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n751), .A2(new_n270), .B1(new_n757), .B2(new_n1099), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G50), .B2(new_n762), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n300), .B1(new_n744), .B2(new_n819), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n738), .B2(new_n1093), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G132), .A2(new_n769), .B1(new_n749), .B2(G58), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1194), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n735), .A2(new_n400), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1192), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n732), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(G68), .B2(new_n809), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n731), .B(new_n1202), .C1(new_n1077), .C2(new_n785), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1079), .A2(new_n1062), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1069), .A2(new_n1078), .B1(new_n800), .B2(new_n838), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1203), .B1(new_n1207), .B2(new_n727), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1075), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1210), .A2(new_n970), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1208), .B1(new_n1211), .B2(new_n1083), .ZN(G381));
  AND2_X1   g1012(.A1(new_n1112), .A2(new_n1087), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1158), .A2(new_n1184), .A3(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(G381), .A2(G387), .ZN(new_n1215));
  NOR4_X1   g1015(.A1(G384), .A2(G390), .A3(G393), .A4(G396), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(G407));
  INV_X1    g1017(.A(G213), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1214), .B2(new_n669), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(G407), .ZN(G409));
  INV_X1    g1020(.A(new_n997), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n952), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n950), .B(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1221), .B1(new_n1223), .B2(new_n971), .ZN(new_n1224));
  OAI21_X1  g1024(.A(KEYINPUT125), .B1(new_n1224), .B2(G390), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT124), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1226), .A3(G390), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n973), .A2(new_n997), .A3(G390), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT124), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT125), .ZN(new_n1230));
  INV_X1    g1030(.A(G390), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(G387), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1225), .A2(new_n1227), .A3(new_n1229), .A4(new_n1232), .ZN(new_n1233));
  XOR2_X1   g1033(.A(G393), .B(G396), .Z(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1224), .A2(G390), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1228), .ZN(new_n1237));
  OR3_X1    g1037(.A1(new_n1234), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1235), .A2(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1218), .A2(G343), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1158), .A2(G378), .A3(new_n1184), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1143), .A2(new_n727), .A3(new_n1145), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(new_n1182), .C1(new_n970), .C2(new_n1155), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1213), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1240), .B1(new_n1241), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT62), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1210), .A2(KEYINPUT60), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1210), .A2(KEYINPUT60), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1247), .A2(new_n1248), .A3(new_n717), .A4(new_n1084), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1249), .A2(G384), .A3(new_n1208), .ZN(new_n1250));
  AOI21_X1  g1050(.A(G384), .B1(new_n1249), .B2(new_n1208), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1245), .A2(new_n1246), .A3(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1246), .B1(new_n1245), .B2(new_n1252), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1240), .A2(G2897), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1252), .A2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G2897), .B(new_n1240), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1240), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1259), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1262), .A2(KEYINPUT61), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1239), .B1(new_n1255), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1245), .A2(new_n1252), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1265), .B1(new_n1262), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT61), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT126), .B1(new_n1239), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1252), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1240), .B(new_n1270), .C1(new_n1241), .C2(new_n1244), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1269), .B1(new_n1271), .B2(KEYINPUT63), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1239), .A2(KEYINPUT126), .A3(new_n1268), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1267), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(KEYINPUT127), .B1(new_n1264), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT127), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1267), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1277));
  NOR4_X1   g1077(.A1(new_n1253), .A2(new_n1254), .A3(KEYINPUT61), .A4(new_n1262), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1276), .B(new_n1277), .C1(new_n1278), .C2(new_n1239), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1275), .A2(new_n1279), .ZN(G405));
  NAND2_X1  g1080(.A1(G375), .A2(new_n1213), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1281), .A2(new_n1241), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(new_n1252), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(new_n1239), .ZN(G402));
endmodule


