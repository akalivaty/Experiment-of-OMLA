//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(new_n203), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n210), .A2(new_n211), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n201), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n208), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n218), .B1(new_n211), .B2(new_n210), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT65), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n216), .A2(G33), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n215), .B1(new_n208), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G13), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(G1), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n201), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n254), .B1(new_n260), .B2(G20), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n259), .B1(new_n261), .B2(new_n201), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  XOR2_X1   g0063(.A(new_n263), .B(KEYINPUT9), .Z(new_n264));
  NAND2_X1  g0064(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G33), .ZN(new_n267));
  AND3_X1   g0067(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT68), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT68), .B1(new_n265), .B2(new_n267), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G223), .A3(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(G222), .A3(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n271), .B(new_n273), .C1(new_n221), .C2(new_n270), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(new_n215), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT69), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT69), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n274), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(G274), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n280), .A2(new_n284), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n286), .B1(new_n288), .B2(G226), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT67), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n283), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n264), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  OR3_X1    g0096(.A1(new_n294), .A2(KEYINPUT10), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT10), .B1(new_n294), .B2(new_n296), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n263), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n291), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n300), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G20), .A2(G77), .ZN(new_n306));
  INV_X1    g0106(.A(new_n248), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT15), .B(G87), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n306), .B1(new_n250), .B2(new_n307), .C1(new_n251), .C2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n309), .A2(new_n254), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n261), .A2(G77), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(G77), .B2(new_n258), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT68), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n266), .A2(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT68), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n318), .A2(G238), .A3(G1698), .A4(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n318), .A2(G232), .A3(new_n272), .A4(new_n319), .ZN(new_n321));
  INV_X1    g0121(.A(G107), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n320), .B(new_n321), .C1(new_n270), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n282), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n286), .B1(new_n288), .B2(G244), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n324), .A2(G179), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n301), .B1(new_n324), .B2(new_n325), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n314), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n324), .A2(new_n295), .A3(new_n325), .ZN(new_n329));
  AOI21_X1  g0129(.A(G200), .B1(new_n324), .B2(new_n325), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n313), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n305), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n318), .A2(G226), .A3(new_n272), .A4(new_n319), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n318), .A2(G232), .A3(G1698), .A4(new_n319), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G97), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n282), .ZN(new_n338));
  INV_X1    g0138(.A(new_n286), .ZN(new_n339));
  INV_X1    g0139(.A(G238), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n287), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n333), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  AOI211_X1 g0143(.A(KEYINPUT13), .B(new_n341), .C1(new_n337), .C2(new_n282), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT14), .B1(new_n345), .B2(new_n301), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n338), .A2(new_n342), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT13), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n338), .A2(new_n333), .A3(new_n342), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT14), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(G169), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n345), .A2(G179), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n346), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n257), .A2(G20), .A3(new_n203), .ZN(new_n355));
  XOR2_X1   g0155(.A(new_n355), .B(KEYINPUT12), .Z(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(G68), .B2(new_n261), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n248), .A2(KEYINPUT71), .A3(G50), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n358), .B1(new_n216), .B2(G68), .C1(new_n221), .C2(new_n251), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT71), .B1(new_n248), .B2(G50), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n254), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT11), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n362), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n357), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n354), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT70), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n345), .B2(new_n293), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n350), .A2(KEYINPUT70), .A3(G200), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n365), .B1(new_n345), .B2(G190), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n299), .A2(new_n332), .A3(new_n366), .A4(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n339), .B1(new_n287), .B2(new_n233), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n272), .A2(G223), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n220), .B2(new_n272), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT3), .B(G33), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G87), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n378), .B1(new_n253), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n374), .B1(new_n282), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n295), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(G200), .B2(new_n381), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n258), .A2(new_n250), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n261), .B2(new_n250), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G58), .A2(G68), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n212), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G20), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT73), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT73), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n390), .A3(G20), .ZN(new_n391));
  INV_X1    g0191(.A(G159), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n389), .B(new_n391), .C1(new_n392), .C2(new_n307), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n216), .B1(new_n268), .B2(new_n269), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n267), .A2(KEYINPUT74), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT74), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(new_n266), .A3(G33), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n265), .A3(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n395), .A2(G20), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n203), .B1(new_n396), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT75), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n393), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n394), .A2(new_n395), .B1(new_n400), .B2(new_n401), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT75), .B1(new_n406), .B2(new_n203), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT16), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n265), .A2(new_n267), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(KEYINPUT7), .A3(new_n216), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT72), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT72), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n409), .A2(new_n412), .A3(KEYINPUT7), .A4(new_n216), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n395), .B1(new_n377), .B2(G20), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G68), .ZN(new_n416));
  INV_X1    g0216(.A(new_n393), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT16), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n254), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n383), .B(new_n385), .C1(new_n408), .C2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n385), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT16), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n318), .A2(new_n319), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT7), .B1(new_n425), .B2(new_n216), .ZN(new_n426));
  INV_X1    g0226(.A(new_n402), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n404), .B(G68), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n417), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n396), .A2(new_n402), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n404), .B1(new_n430), .B2(G68), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n424), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n254), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n393), .B1(G68), .B2(new_n415), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(KEYINPUT16), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n423), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(KEYINPUT17), .A3(new_n383), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n422), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n381), .A2(G169), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(new_n303), .B2(new_n381), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT18), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT76), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT18), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n407), .A2(new_n428), .A3(new_n417), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n419), .B1(new_n424), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n445), .B(new_n441), .C1(new_n447), .C2(new_n423), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n443), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n444), .B1(new_n443), .B2(new_n448), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n439), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n373), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n322), .A2(G20), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT23), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G116), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n454), .B1(new_n216), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n377), .A2(new_n216), .A3(G87), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT86), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT22), .ZN(new_n460));
  OR3_X1    g0260(.A1(new_n379), .A2(KEYINPUT22), .A3(G20), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n425), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n459), .B1(new_n458), .B2(KEYINPUT22), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n457), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT24), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(KEYINPUT24), .B(new_n457), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n466), .A2(new_n254), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n257), .A2(G20), .A3(new_n322), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n469), .B(KEYINPUT25), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n260), .A2(G33), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n433), .A2(new_n258), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(G107), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G257), .A2(G1698), .ZN(new_n474));
  INV_X1    g0274(.A(G250), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(G1698), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n377), .A2(new_n476), .B1(G33), .B2(G294), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n260), .A2(G45), .ZN(new_n479));
  OR2_X1    g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  NAND2_X1  g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(new_n277), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n282), .A2(new_n478), .B1(new_n483), .B2(G264), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(G274), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(G179), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(G264), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n279), .A2(new_n281), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n485), .C1(new_n488), .C2(new_n477), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G169), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n468), .A2(new_n473), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT87), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n293), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(G190), .B2(new_n489), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n468), .A2(new_n473), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n492), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n496), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT87), .B1(new_n498), .B2(new_n491), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n253), .A2(G97), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G283), .ZN(new_n502));
  AOI21_X1  g0302(.A(G20), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G116), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n216), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n254), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT20), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(KEYINPUT20), .B(new_n254), .C1(new_n503), .C2(new_n505), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n258), .A2(new_n504), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n472), .B2(new_n504), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G169), .ZN(new_n514));
  AND2_X1   g0314(.A1(G264), .A2(G1698), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n265), .A2(new_n267), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT84), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n377), .A2(KEYINPUT84), .A3(new_n515), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n377), .A2(G257), .A3(new_n272), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G303), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n318), .B2(new_n319), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n282), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n483), .A2(G270), .B1(G274), .B2(new_n482), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT85), .B1(new_n514), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT21), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT21), .ZN(new_n530));
  OAI211_X1 g0330(.A(KEYINPUT85), .B(new_n530), .C1(new_n514), .C2(new_n527), .ZN(new_n531));
  INV_X1    g0331(.A(new_n513), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n526), .A2(G190), .ZN(new_n533));
  AOI21_X1  g0333(.A(G200), .B1(new_n524), .B2(new_n525), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n524), .A2(G179), .A3(new_n525), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n513), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n529), .A2(new_n531), .A3(new_n535), .A4(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n308), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n472), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n540), .A2(new_n258), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G87), .A2(G97), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n543), .A2(new_n322), .B1(new_n336), .B2(new_n216), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n216), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n544), .A2(new_n545), .B1(new_n336), .B2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n377), .A2(KEYINPUT81), .A3(new_n216), .A4(G68), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n265), .A2(new_n267), .A3(new_n216), .A4(G68), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT81), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n542), .B1(new_n552), .B2(new_n254), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT82), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI211_X1 g0355(.A(KEYINPUT82), .B(new_n542), .C1(new_n552), .C2(new_n254), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n541), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n479), .A2(G250), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n260), .A2(G45), .A3(G274), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n277), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n377), .A2(G238), .A3(new_n272), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n377), .A2(G244), .A3(G1698), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(new_n455), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n560), .B1(new_n282), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G179), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n301), .B2(new_n564), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n557), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n282), .A2(new_n563), .ZN(new_n568));
  INV_X1    g0368(.A(new_n560), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n295), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(G200), .B2(new_n564), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n472), .A2(G87), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n556), .C2(new_n555), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT83), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n567), .A2(KEYINPUT83), .A3(new_n573), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n539), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g0378(.A(KEYINPUT77), .B(KEYINPUT6), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n322), .A2(G97), .ZN(new_n580));
  INV_X1    g0380(.A(G97), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G107), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  OR2_X1    g0383(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n584));
  NAND2_X1  g0384(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n584), .A2(G97), .A3(new_n322), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT78), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT78), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n583), .A2(new_n589), .A3(new_n586), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(G20), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n248), .A2(G77), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n591), .B(new_n592), .C1(new_n322), .C2(new_n406), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n258), .A2(new_n581), .ZN(new_n594));
  OR2_X1    g0394(.A1(new_n472), .A2(new_n581), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n593), .A2(new_n254), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n483), .A2(G257), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n485), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT4), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(new_n222), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n318), .A2(new_n272), .A3(new_n319), .A4(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n318), .A2(G250), .A3(G1698), .A4(new_n319), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n377), .A2(G244), .A3(new_n272), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n599), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n601), .A2(new_n602), .A3(new_n604), .A4(new_n502), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n598), .B1(new_n605), .B2(new_n282), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G190), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(KEYINPUT79), .A3(new_n282), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT79), .B1(new_n605), .B2(new_n282), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n609), .A2(new_n610), .A3(new_n598), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n596), .B(new_n607), .C1(new_n611), .C2(new_n293), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT80), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n591), .A2(new_n592), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n406), .A2(new_n322), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n254), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n595), .A2(new_n594), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n610), .ZN(new_n619));
  INV_X1    g0419(.A(new_n598), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n619), .A2(new_n303), .A3(new_n608), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n605), .A2(new_n282), .ZN(new_n622));
  AOI21_X1  g0422(.A(G169), .B1(new_n622), .B2(new_n620), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n618), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n612), .A2(new_n613), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n613), .B1(new_n612), .B2(new_n625), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n452), .A2(new_n500), .A3(new_n578), .A4(new_n628), .ZN(G372));
  INV_X1    g0429(.A(new_n305), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n385), .B1(new_n408), .B2(new_n419), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n445), .B1(new_n631), .B2(new_n441), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n436), .A2(KEYINPUT18), .A3(new_n442), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n366), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n328), .A2(KEYINPUT90), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT90), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n637), .B(new_n314), .C1(new_n326), .C2(new_n327), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n635), .B1(new_n372), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n634), .B1(new_n640), .B2(new_n438), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n299), .A2(KEYINPUT91), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT91), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n297), .A2(new_n643), .A3(new_n298), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n630), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n452), .ZN(new_n647));
  INV_X1    g0447(.A(new_n612), .ZN(new_n648));
  INV_X1    g0448(.A(new_n625), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n498), .A2(new_n574), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n529), .A2(new_n538), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n531), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n650), .B(new_n651), .C1(new_n653), .C2(new_n491), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  INV_X1    g0456(.A(new_n574), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT88), .ZN(new_n658));
  AND4_X1   g0458(.A1(new_n658), .A2(new_n618), .A3(new_n621), .A4(new_n624), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n623), .B1(new_n616), .B2(new_n617), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n658), .B1(new_n660), .B2(new_n621), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n656), .B(new_n657), .C1(new_n659), .C2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n625), .B1(new_n576), .B2(new_n577), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n662), .B(new_n567), .C1(new_n663), .C2(new_n656), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT89), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n567), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n567), .A2(KEYINPUT83), .A3(new_n573), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT83), .B1(new_n567), .B2(new_n573), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n649), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n667), .B1(new_n670), .B2(KEYINPUT26), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(KEYINPUT89), .A3(new_n662), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n655), .B1(new_n666), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n646), .B1(new_n647), .B2(new_n673), .ZN(G369));
  NOR2_X1   g0474(.A1(new_n256), .A2(G20), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n260), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT92), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT27), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G213), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n677), .B2(new_n678), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT93), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(G343), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(G343), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(KEYINPUT94), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT94), .ZN(new_n689));
  INV_X1    g0489(.A(new_n687), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(new_n682), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n652), .A2(new_n513), .A3(new_n531), .A4(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n692), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n539), .B1(new_n532), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n468), .A2(new_n473), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n692), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT95), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n701), .A2(new_n500), .B1(new_n491), .B2(new_n692), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n500), .A2(new_n701), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n653), .A2(new_n694), .ZN(new_n705));
  OAI22_X1  g0505(.A1(new_n704), .A2(new_n705), .B1(new_n492), .B2(new_n692), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n703), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n209), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G1), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n543), .A2(new_n322), .A3(new_n504), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n711), .A2(new_n712), .B1(new_n213), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  INV_X1    g0514(.A(G330), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n622), .A2(new_n620), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n484), .A2(new_n564), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n716), .A2(new_n536), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n619), .A2(new_n608), .A3(new_n620), .ZN(new_n719));
  INV_X1    g0519(.A(new_n564), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n526), .A2(new_n720), .A3(new_n303), .A4(new_n489), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI22_X1  g0522(.A1(KEYINPUT30), .A2(new_n718), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n484), .A2(new_n564), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n537), .A2(new_n724), .A3(new_n606), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g0528(.A(KEYINPUT96), .B(KEYINPUT31), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(new_n692), .A3(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT97), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n725), .A2(new_n732), .A3(new_n726), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n732), .B1(new_n725), .B2(new_n726), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n723), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT31), .B1(new_n736), .B2(new_n692), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT98), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n731), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n611), .A2(new_n721), .B1(new_n725), .B2(new_n726), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n727), .A2(KEYINPUT97), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n740), .B1(new_n741), .B2(new_n733), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n694), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n743), .A2(KEYINPUT98), .A3(KEYINPUT31), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n628), .A2(new_n500), .A3(new_n578), .A4(new_n694), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n715), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n666), .A2(new_n672), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n692), .B1(new_n748), .B2(new_n654), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT29), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n663), .A2(new_n656), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n567), .B(KEYINPUT99), .Z(new_n752));
  NAND3_X1  g0552(.A1(new_n654), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n659), .A2(new_n661), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n656), .B1(new_n754), .B2(new_n657), .ZN(new_n755));
  OAI211_X1 g0555(.A(KEYINPUT29), .B(new_n694), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n747), .B1(new_n750), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n714), .B1(new_n757), .B2(G1), .ZN(G364));
  NOR2_X1   g0558(.A1(G13), .A2(G33), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n696), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n711), .B1(G45), .B2(new_n675), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n215), .B1(G20), .B2(new_n301), .ZN(new_n764));
  NAND2_X1  g0564(.A1(G20), .A2(G179), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT101), .Z(new_n766));
  NOR2_X1   g0566(.A1(new_n295), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n293), .A2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G20), .A3(G190), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT102), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G322), .A2(new_n769), .B1(new_n772), .B2(G303), .ZN(new_n773));
  INV_X1    g0573(.A(G326), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n295), .A2(new_n293), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n766), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n773), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n216), .A2(G190), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n770), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G283), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G179), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G329), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n779), .A2(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n781), .A2(G190), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n784), .B(new_n270), .C1(G294), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n766), .A2(new_n295), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n293), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(KEYINPUT33), .B(G317), .Z(new_n791));
  OAI21_X1  g0591(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n788), .A2(G200), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n777), .B(new_n792), .C1(G311), .C2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n786), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n581), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n771), .A2(new_n379), .B1(new_n779), .B2(new_n322), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n796), .A2(new_n797), .A3(new_n425), .ZN(new_n798));
  INV_X1    g0598(.A(new_n793), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n798), .B1(new_n799), .B2(new_n221), .C1(new_n203), .C2(new_n790), .ZN(new_n800));
  INV_X1    g0600(.A(new_n782), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G159), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT32), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n201), .A2(new_n776), .B1(new_n768), .B2(new_n202), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n800), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n764), .B1(new_n794), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n761), .A2(new_n764), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n708), .A2(new_n377), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n242), .A2(G45), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n214), .A2(G45), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n425), .A2(new_n708), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G355), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(G116), .B2(new_n209), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n807), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n762), .A2(new_n763), .A3(new_n806), .A4(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n697), .A2(G330), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(KEYINPUT100), .ZN(new_n819));
  INV_X1    g0619(.A(new_n763), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n818), .B1(new_n698), .B2(KEYINPUT100), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n817), .B1(new_n821), .B2(new_n822), .ZN(G396));
  AOI21_X1  g0623(.A(new_n313), .B1(new_n688), .B2(new_n691), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n636), .A2(new_n638), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT106), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n636), .A2(KEYINPUT106), .A3(new_n638), .A4(new_n824), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT105), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n328), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(KEYINPUT105), .B(new_n314), .C1(new_n326), .C2(new_n327), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n692), .A2(new_n314), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n834), .A2(new_n331), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n827), .A2(new_n828), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n749), .A2(new_n837), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n673), .A2(new_n692), .A3(new_n836), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n763), .B1(new_n840), .B2(new_n747), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n747), .B2(new_n840), .ZN(new_n842));
  INV_X1    g0642(.A(G311), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n425), .B1(new_n379), .B2(new_n779), .C1(new_n843), .C2(new_n782), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n796), .B(new_n844), .C1(G283), .C2(new_n789), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n504), .B2(new_n799), .ZN(new_n846));
  INV_X1    g0646(.A(new_n776), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G303), .A2(new_n847), .B1(new_n772), .B2(G107), .ZN(new_n848));
  INV_X1    g0648(.A(G294), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(new_n768), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT104), .Z(new_n852));
  AOI22_X1  g0652(.A1(G137), .A2(new_n847), .B1(new_n769), .B2(G143), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n392), .B2(new_n799), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(G150), .B2(new_n789), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n855), .A2(KEYINPUT34), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(KEYINPUT34), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n409), .B1(new_n801), .B2(G132), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n858), .B1(new_n202), .B2(new_n795), .C1(new_n203), .C2(new_n779), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(G50), .B2(new_n772), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n856), .A2(new_n857), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n764), .B1(new_n852), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n764), .A2(new_n759), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT103), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n820), .B1(new_n865), .B2(new_n221), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n862), .B(new_n866), .C1(new_n837), .C2(new_n760), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n842), .A2(new_n867), .ZN(G384));
  NAND2_X1  g0668(.A1(new_n386), .A2(G77), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n213), .A2(new_n869), .B1(G50), .B2(new_n203), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(G1), .A3(new_n256), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT107), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n217), .A2(G116), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n588), .A2(new_n590), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT35), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n875), .B2(new_n874), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT36), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n878), .B2(new_n877), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT110), .B1(new_n742), .B2(new_n694), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT110), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n736), .A2(new_n882), .A3(new_n692), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n729), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n743), .A2(KEYINPUT31), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n746), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n366), .A2(KEYINPUT108), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n370), .A2(new_n371), .B1(new_n365), .B2(new_n692), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT108), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n354), .A2(new_n889), .A3(new_n365), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n888), .A2(new_n366), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n836), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n886), .A2(new_n893), .A3(KEYINPUT40), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT111), .ZN(new_n895));
  INV_X1    g0695(.A(new_n420), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n435), .B1(KEYINPUT16), .B2(new_n434), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n897), .A2(new_n385), .B1(new_n442), .B2(new_n682), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT37), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n631), .A2(new_n441), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n683), .B1(new_n447), .B2(new_n423), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT37), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n900), .A2(new_n901), .A3(new_n902), .A4(new_n420), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT76), .B1(new_n632), .B2(new_n633), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n443), .A2(new_n444), .A3(new_n448), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n438), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n897), .A2(new_n385), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n683), .ZN(new_n909));
  OAI211_X1 g0709(.A(KEYINPUT38), .B(new_n904), .C1(new_n907), .C2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n900), .A2(new_n901), .A3(new_n420), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n903), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n443), .A2(new_n422), .A3(new_n437), .A4(new_n448), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n631), .A3(new_n683), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT38), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n910), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n894), .A2(new_n895), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n913), .B2(new_n915), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n899), .A2(new_n903), .ZN(new_n922));
  INV_X1    g0722(.A(new_n909), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n922), .B1(new_n451), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n921), .B1(new_n924), .B2(KEYINPUT38), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n886), .A2(new_n893), .A3(KEYINPUT40), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT111), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n886), .A2(new_n893), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n924), .A2(KEYINPUT38), .ZN(new_n929));
  INV_X1    g0729(.A(new_n910), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n920), .A2(new_n927), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT112), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n452), .A2(new_n886), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(G330), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n891), .A2(new_n892), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n664), .A2(new_n665), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT89), .B1(new_n671), .B2(new_n662), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n654), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(new_n694), .A3(new_n837), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n833), .A2(new_n692), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n940), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n904), .B1(new_n907), .B2(new_n909), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n917), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n910), .ZN(new_n950));
  INV_X1    g0750(.A(new_n634), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n947), .A2(new_n950), .B1(new_n951), .B2(new_n682), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n887), .A2(new_n890), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(new_n692), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT39), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n910), .A2(new_n918), .A3(new_n955), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n950), .A2(KEYINPUT39), .B1(new_n956), .B2(KEYINPUT109), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT109), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n958), .B(new_n955), .C1(new_n949), .C2(new_n910), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n954), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n952), .A2(new_n960), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n452), .B(new_n756), .C1(new_n749), .C2(KEYINPUT29), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n646), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n961), .B(new_n963), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n938), .A2(new_n964), .B1(new_n260), .B2(new_n675), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT113), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n938), .A2(new_n964), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n965), .A2(KEYINPUT113), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n880), .B1(new_n968), .B2(new_n969), .ZN(G367));
  NOR2_X1   g0770(.A1(new_n237), .A2(new_n809), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n807), .B1(new_n209), .B2(new_n308), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n763), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n771), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n974), .A2(G58), .B1(new_n801), .B2(G137), .ZN(new_n975));
  INV_X1    g0775(.A(G150), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n975), .B1(new_n203), .B2(new_n795), .C1(new_n768), .C2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G143), .B2(new_n847), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G50), .A2(new_n793), .B1(new_n789), .B2(G159), .ZN(new_n979));
  INV_X1    g0779(.A(new_n779), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n425), .B1(G77), .B2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT114), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(KEYINPUT114), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n978), .A2(new_n979), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT46), .B1(new_n974), .B2(G116), .ZN(new_n985));
  INV_X1    g0785(.A(G317), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n409), .B1(new_n782), .B2(new_n986), .C1(new_n581), .C2(new_n779), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n985), .B(new_n987), .C1(G107), .C2(new_n786), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n780), .B2(new_n799), .C1(new_n849), .C2(new_n790), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n772), .A2(KEYINPUT46), .A3(G116), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n522), .B2(new_n768), .C1(new_n843), .C2(new_n776), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n984), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT47), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n994), .A2(new_n764), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(new_n993), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n973), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n761), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n572), .B1(new_n555), .B2(new_n556), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n692), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n667), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n574), .B2(new_n1000), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n997), .B1(new_n998), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n260), .B1(new_n675), .B2(G45), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n650), .B1(new_n596), .B2(new_n694), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n649), .A2(new_n692), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n706), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT45), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n706), .A2(new_n1009), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT44), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n703), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n698), .B(new_n702), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(new_n705), .Z(new_n1019));
  AND2_X1   g0819(.A1(new_n757), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n757), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n709), .B(KEYINPUT41), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1005), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n1009), .A2(new_n702), .A3(new_n705), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT42), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n649), .B1(new_n491), .B2(new_n612), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n692), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1025), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n703), .A2(new_n1008), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1003), .B1(new_n1024), .B2(new_n1036), .ZN(G387));
  INV_X1    g0837(.A(new_n250), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G68), .A2(new_n793), .B1(new_n789), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n795), .A2(new_n308), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n377), .B1(new_n779), .B2(new_n581), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n771), .A2(new_n221), .B1(new_n782), .B2(new_n976), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G50), .A2(new_n769), .B1(new_n847), .B2(G159), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1039), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n377), .B1(new_n980), .B2(G116), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n795), .A2(new_n780), .B1(new_n771), .B2(new_n849), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G317), .A2(new_n769), .B1(new_n847), .B2(G322), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n522), .B2(new_n799), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G311), .B2(new_n789), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1047), .B1(new_n1050), .B2(KEYINPUT48), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(KEYINPUT48), .B2(new_n1050), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1046), .B1(new_n774), .B2(new_n782), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1045), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n764), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n702), .A2(new_n761), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n809), .B1(new_n234), .B2(G45), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n712), .B2(new_n813), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1038), .A2(new_n201), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT50), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n203), .A2(new_n221), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1062), .A2(G45), .A3(new_n1063), .A4(new_n712), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n1060), .A2(new_n1064), .B1(G107), .B2(new_n209), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n820), .B1(new_n1065), .B2(new_n807), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1057), .A2(new_n1058), .A3(new_n1066), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT115), .Z(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1019), .B2(new_n1005), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1020), .A2(new_n710), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n757), .A2(new_n1019), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(G393));
  NAND2_X1  g0872(.A1(new_n1017), .A2(new_n1005), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1009), .A2(new_n761), .ZN(new_n1074));
  INV_X1    g0874(.A(G322), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n779), .A2(new_n322), .B1(new_n782), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n425), .B1(new_n504), .B2(new_n795), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(G283), .C2(new_n974), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(new_n849), .B2(new_n799), .C1(new_n522), .C2(new_n790), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n843), .A2(new_n768), .B1(new_n776), .B2(new_n986), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT52), .Z(new_n1081));
  OAI22_X1  g0881(.A1(new_n976), .A2(new_n776), .B1(new_n768), .B2(new_n392), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT51), .Z(new_n1083));
  OAI21_X1  g0883(.A(new_n377), .B1(new_n779), .B2(new_n379), .ZN(new_n1084));
  INV_X1    g0884(.A(G143), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n771), .A2(new_n203), .B1(new_n782), .B2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1084), .B(new_n1086), .C1(G77), .C2(new_n786), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n799), .B2(new_n250), .C1(new_n201), .C2(new_n790), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1079), .A2(new_n1081), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n764), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n807), .B1(new_n581), .B2(new_n209), .C1(new_n246), .C2(new_n809), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1074), .A2(new_n763), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1021), .A2(new_n709), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1073), .B(new_n1092), .C1(new_n1093), .C2(new_n1094), .ZN(G390));
  OAI211_X1 g0895(.A(new_n694), .B(new_n837), .C1(new_n753), .C2(new_n755), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n946), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n939), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n954), .B(KEYINPUT116), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1098), .A2(new_n1099), .A3(new_n919), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n747), .A2(new_n893), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n944), .A2(new_n946), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n954), .B1(new_n1102), .B2(new_n939), .ZN(new_n1103));
  OAI211_X1 g0903(.A(KEYINPUT109), .B(KEYINPUT39), .C1(new_n929), .C2(new_n930), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n958), .B1(new_n925), .B2(new_n955), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n955), .B1(new_n949), .B2(new_n910), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1100), .B(new_n1101), .C1(new_n1103), .C2(new_n1107), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1098), .A2(new_n1099), .A3(new_n919), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n957), .A2(new_n959), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n954), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n945), .B1(new_n749), .B2(new_n837), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1111), .B1(new_n1112), .B2(new_n940), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1109), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n886), .A2(G330), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n893), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1108), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(new_n1004), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1110), .A2(new_n759), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n763), .B1(new_n864), .B2(new_n1038), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n974), .A2(G150), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT53), .ZN(new_n1124));
  INV_X1    g0924(.A(G128), .ZN(new_n1125));
  INV_X1    g0925(.A(G132), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1125), .A2(new_n776), .B1(new_n768), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n793), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n789), .A2(G137), .ZN(new_n1132));
  INV_X1    g0932(.A(G125), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n779), .A2(new_n201), .B1(new_n782), .B2(new_n1133), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n425), .B(new_n1134), .C1(G159), .C2(new_n786), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1128), .A2(new_n1131), .A3(new_n1132), .A4(new_n1135), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n790), .A2(new_n322), .B1(new_n776), .B2(new_n780), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G97), .B2(new_n793), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT118), .Z(new_n1139));
  AOI22_X1  g0939(.A1(G116), .A2(new_n769), .B1(new_n772), .B2(G87), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n786), .A2(G77), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n779), .A2(new_n203), .B1(new_n782), .B2(new_n849), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n270), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1136), .B1(new_n1139), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1122), .B1(new_n1145), .B2(new_n764), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1120), .B1(new_n1121), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n452), .A2(new_n886), .A3(G330), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n962), .A2(new_n646), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1097), .B1(new_n747), .B2(new_n893), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT117), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1115), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n886), .A2(KEYINPUT117), .A3(G330), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n836), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1150), .B1(new_n1154), .B2(new_n939), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n939), .B1(new_n747), .B2(new_n837), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1102), .B1(new_n1156), .B2(new_n1117), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1149), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1119), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1108), .B(new_n1158), .C1(new_n1114), .C2(new_n1118), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n709), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1147), .A2(new_n1162), .ZN(G378));
  NOR2_X1   g0963(.A1(new_n682), .A2(new_n263), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n642), .A2(new_n305), .A3(new_n644), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(KEYINPUT119), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1165), .A2(KEYINPUT119), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1164), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1168), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1164), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n1166), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g0973(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1174), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1169), .A2(new_n1172), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT120), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1175), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n927), .A2(new_n920), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n931), .A2(new_n932), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(G330), .A3(new_n1181), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n952), .A2(new_n1182), .A3(new_n960), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(new_n960), .B2(new_n952), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1179), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT39), .B1(new_n929), .B2(new_n930), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n956), .A2(KEYINPUT109), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1111), .B1(new_n1188), .B2(new_n1104), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n950), .B(new_n939), .C1(new_n839), .C2(new_n945), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n951), .A2(new_n682), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(G330), .B(new_n933), .C1(new_n1189), .C2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n952), .A2(new_n1182), .A3(new_n960), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1179), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1149), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1185), .A2(new_n1196), .B1(new_n1197), .B2(new_n1161), .ZN(new_n1198));
  OAI21_X1  g0998(.A(KEYINPUT122), .B1(new_n1198), .B2(KEYINPUT57), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1161), .A2(new_n1197), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1195), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1200), .B(KEYINPUT57), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT121), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1198), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1199), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT122), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1200), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1208), .B(new_n1209), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n709), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1207), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1185), .A2(new_n1196), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1175), .A2(new_n1177), .A3(new_n759), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n763), .B1(new_n864), .B2(G50), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G97), .A2(new_n789), .B1(new_n793), .B2(new_n540), .ZN(new_n1218));
  INV_X1    g1018(.A(G41), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n409), .C1(new_n782), .C2(new_n780), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n771), .A2(new_n221), .B1(new_n779), .B2(new_n202), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(G68), .C2(new_n786), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G107), .A2(new_n769), .B1(new_n847), .B2(G116), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1218), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n409), .A2(new_n1219), .ZN(new_n1226));
  AOI21_X1  g1026(.A(G50), .B1(new_n253), .B2(new_n1219), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1225), .A2(KEYINPUT58), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n790), .A2(new_n1126), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n974), .A2(new_n1130), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n786), .A2(G150), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n776), .B2(new_n1133), .C1(new_n1125), .C2(new_n768), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1229), .B(new_n1233), .C1(G137), .C2(new_n793), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n253), .B(new_n1219), .C1(new_n779), .C2(new_n392), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G124), .B2(new_n801), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT59), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1238), .B1(new_n1234), .B2(new_n1239), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1228), .B1(KEYINPUT58), .B2(new_n1225), .C1(new_n1236), .C2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1217), .B1(new_n1241), .B2(new_n764), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1215), .A2(new_n1005), .B1(new_n1216), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1214), .A2(new_n1243), .ZN(G375));
  NAND2_X1  g1044(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1005), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n779), .A2(new_n221), .B1(new_n782), .B2(new_n522), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1040), .A2(new_n270), .A3(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n790), .B2(new_n504), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G283), .A2(new_n769), .B1(new_n772), .B2(G97), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n849), .B2(new_n776), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1249), .B(new_n1251), .C1(G107), .C2(new_n793), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n847), .A2(G132), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(KEYINPUT124), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n377), .B1(new_n782), .B2(new_n1125), .C1(new_n202), .C2(new_n779), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G50), .B2(new_n786), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(G137), .A2(new_n769), .B1(new_n772), .B2(G159), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G150), .A2(new_n793), .B1(new_n789), .B2(new_n1130), .ZN(new_n1258));
  AND4_X1   g1058(.A1(new_n1254), .A2(new_n1256), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n764), .B1(new_n1252), .B2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n820), .B1(new_n865), .B2(new_n203), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(new_n939), .C2(new_n760), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1246), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1155), .A2(new_n1149), .A3(new_n1157), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1023), .B(KEYINPUT123), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1159), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1268), .B(KEYINPUT125), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(G381));
  INV_X1    g1070(.A(G375), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G378), .A2(KEYINPUT126), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT126), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1147), .A2(new_n1273), .A3(new_n1162), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(G387), .A2(G390), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1276), .A2(new_n1269), .A3(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1271), .A2(new_n1275), .A3(new_n1278), .ZN(G407));
  NOR2_X1   g1079(.A1(new_n687), .A2(new_n680), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1271), .A2(new_n1275), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(G407), .A2(new_n1281), .A3(G213), .ZN(G409));
  OAI211_X1 g1082(.A(G378), .B(new_n1243), .C1(new_n1207), .C2(new_n1213), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1198), .A2(new_n1266), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1243), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1272), .A2(new_n1274), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1280), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1265), .A2(KEYINPUT60), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1265), .A2(KEYINPUT60), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n709), .B(new_n1159), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1264), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n842), .A2(new_n867), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1291), .A2(G384), .A3(new_n1264), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT127), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1294), .A2(KEYINPUT127), .A3(new_n1295), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1297), .A2(G2897), .A3(new_n1280), .A4(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1280), .A2(G2897), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1298), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1300), .B1(new_n1301), .B2(new_n1296), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(KEYINPUT63), .B1(new_n1287), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1287), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1276), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(G387), .A2(G390), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  XOR2_X1   g1111(.A(G393), .B(G396), .Z(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1312), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1309), .A2(new_n1315), .A3(new_n1310), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1313), .A2(new_n1314), .A3(new_n1316), .ZN(new_n1317));
  AOI211_X1 g1117(.A(new_n1280), .B(new_n1305), .C1(new_n1283), .C2(new_n1286), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1317), .B1(new_n1318), .B2(KEYINPUT63), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1308), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1287), .A2(new_n1321), .A3(new_n1306), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1314), .B1(new_n1287), .B2(new_n1303), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1321), .B1(new_n1287), .B2(new_n1306), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1322), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1316), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1315), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1320), .B1(new_n1325), .B2(new_n1328), .ZN(G405));
  OAI21_X1  g1129(.A(new_n1305), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1313), .A2(new_n1306), .A3(new_n1316), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G375), .A2(new_n1275), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1283), .ZN(new_n1334));
  XOR2_X1   g1134(.A(new_n1332), .B(new_n1334), .Z(G402));
endmodule


