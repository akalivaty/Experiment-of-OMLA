

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593;

  XOR2_X1 U325 ( .A(n376), .B(n375), .Z(n293) );
  NAND2_X1 U326 ( .A1(n532), .A2(n562), .ZN(n294) );
  XNOR2_X1 U327 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n424) );
  XNOR2_X1 U328 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U329 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n433) );
  XNOR2_X1 U330 ( .A(n434), .B(n433), .ZN(n541) );
  INV_X1 U331 ( .A(G190GAT), .ZN(n461) );
  XNOR2_X1 U332 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U333 ( .A(n464), .B(n463), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(G120GAT), .B(G71GAT), .Z(n366) );
  XOR2_X1 U335 ( .A(KEYINPUT85), .B(KEYINPUT0), .Z(n296) );
  XNOR2_X1 U336 ( .A(G113GAT), .B(KEYINPUT84), .ZN(n295) );
  XNOR2_X1 U337 ( .A(n296), .B(n295), .ZN(n449) );
  XNOR2_X1 U338 ( .A(n366), .B(n449), .ZN(n297) );
  XOR2_X1 U339 ( .A(G15GAT), .B(G127GAT), .Z(n386) );
  XNOR2_X1 U340 ( .A(n297), .B(n386), .ZN(n303) );
  XOR2_X1 U341 ( .A(G183GAT), .B(KEYINPUT17), .Z(n299) );
  XNOR2_X1 U342 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n299), .B(n298), .ZN(n351) );
  XOR2_X1 U344 ( .A(KEYINPUT86), .B(n351), .Z(n301) );
  NAND2_X1 U345 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U347 ( .A(n303), .B(n302), .Z(n311) );
  XOR2_X1 U348 ( .A(G99GAT), .B(G134GAT), .Z(n305) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(G190GAT), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U351 ( .A(G176GAT), .B(KEYINPUT20), .Z(n307) );
  XNOR2_X1 U352 ( .A(G169GAT), .B(KEYINPUT87), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U355 ( .A(n311), .B(n310), .Z(n532) );
  XOR2_X1 U356 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n313) );
  XOR2_X1 U357 ( .A(G134GAT), .B(KEYINPUT80), .Z(n448) );
  XOR2_X1 U358 ( .A(G99GAT), .B(G85GAT), .Z(n374) );
  XNOR2_X1 U359 ( .A(n448), .B(n374), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U361 ( .A(n314), .B(KEYINPUT10), .ZN(n319) );
  XOR2_X1 U362 ( .A(KEYINPUT78), .B(KEYINPUT67), .Z(n316) );
  XNOR2_X1 U363 ( .A(G106GAT), .B(KEYINPUT79), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U365 ( .A(G218GAT), .B(n317), .Z(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U367 ( .A(G36GAT), .B(G190GAT), .Z(n358) );
  XOR2_X1 U368 ( .A(n358), .B(G92GAT), .Z(n321) );
  NAND2_X1 U369 ( .A1(G232GAT), .A2(G233GAT), .ZN(n320) );
  XOR2_X1 U370 ( .A(n321), .B(n320), .Z(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n328) );
  XOR2_X1 U372 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n325) );
  XNOR2_X1 U373 ( .A(G43GAT), .B(G29GAT), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U375 ( .A(KEYINPUT70), .B(n326), .Z(n416) );
  XOR2_X1 U376 ( .A(G50GAT), .B(G162GAT), .Z(n332) );
  XNOR2_X1 U377 ( .A(n416), .B(n332), .ZN(n327) );
  XOR2_X1 U378 ( .A(n328), .B(n327), .Z(n562) );
  XOR2_X1 U379 ( .A(KEYINPUT92), .B(G218GAT), .Z(n330) );
  XNOR2_X1 U380 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U382 ( .A(G197GAT), .B(n331), .ZN(n361) );
  XOR2_X1 U383 ( .A(KEYINPUT94), .B(KEYINPUT24), .Z(n334) );
  XOR2_X1 U384 ( .A(G22GAT), .B(G155GAT), .Z(n384) );
  XNOR2_X1 U385 ( .A(n332), .B(n384), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n334), .B(n333), .ZN(n347) );
  XOR2_X1 U387 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n336) );
  XNOR2_X1 U388 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U390 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n338) );
  XNOR2_X1 U391 ( .A(G204GAT), .B(KEYINPUT95), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U393 ( .A(n340), .B(n339), .Z(n345) );
  XNOR2_X1 U394 ( .A(G106GAT), .B(G78GAT), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n341), .B(G148GAT), .ZN(n369) );
  XOR2_X1 U396 ( .A(KEYINPUT93), .B(KEYINPUT3), .Z(n343) );
  XNOR2_X1 U397 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n445) );
  XNOR2_X1 U399 ( .A(n369), .B(n445), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U401 ( .A(n347), .B(n346), .Z(n349) );
  NAND2_X1 U402 ( .A1(G228GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U404 ( .A(n361), .B(n350), .Z(n475) );
  XOR2_X1 U405 ( .A(KEYINPUT81), .B(n351), .Z(n353) );
  NAND2_X1 U406 ( .A1(G226GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U408 ( .A(KEYINPUT75), .B(G64GAT), .Z(n355) );
  XNOR2_X1 U409 ( .A(G204GAT), .B(G92GAT), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U411 ( .A(G176GAT), .B(n356), .Z(n365) );
  XOR2_X1 U412 ( .A(n357), .B(n365), .Z(n360) );
  XOR2_X1 U413 ( .A(G169GAT), .B(G8GAT), .Z(n408) );
  XNOR2_X1 U414 ( .A(n408), .B(n358), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n362) );
  XOR2_X1 U416 ( .A(n362), .B(n361), .Z(n505) );
  INV_X1 U417 ( .A(n505), .ZN(n528) );
  XOR2_X1 U418 ( .A(KEYINPUT73), .B(KEYINPUT33), .Z(n364) );
  XNOR2_X1 U419 ( .A(KEYINPUT31), .B(KEYINPUT74), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n381) );
  XNOR2_X1 U421 ( .A(n366), .B(n365), .ZN(n379) );
  INV_X1 U422 ( .A(n369), .ZN(n368) );
  INV_X1 U423 ( .A(KEYINPUT32), .ZN(n367) );
  NAND2_X1 U424 ( .A1(n368), .A2(n367), .ZN(n371) );
  NAND2_X1 U425 ( .A1(n369), .A2(KEYINPUT32), .ZN(n370) );
  NAND2_X1 U426 ( .A1(n371), .A2(n370), .ZN(n373) );
  AND2_X1 U427 ( .A1(G230GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U429 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n376) );
  XOR2_X1 U430 ( .A(G57GAT), .B(KEYINPUT13), .Z(n385) );
  XNOR2_X1 U431 ( .A(n374), .B(n385), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n377), .B(n293), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n381), .B(n380), .ZN(n423) );
  XOR2_X1 U435 ( .A(G78GAT), .B(G211GAT), .Z(n383) );
  XNOR2_X1 U436 ( .A(G183GAT), .B(G71GAT), .ZN(n382) );
  XNOR2_X1 U437 ( .A(n383), .B(n382), .ZN(n399) );
  XOR2_X1 U438 ( .A(n385), .B(n384), .Z(n388) );
  XOR2_X1 U439 ( .A(G1GAT), .B(KEYINPUT71), .Z(n415) );
  XNOR2_X1 U440 ( .A(n415), .B(n386), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U442 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n390) );
  NAND2_X1 U443 ( .A1(G231GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U445 ( .A(n392), .B(n391), .Z(n397) );
  XOR2_X1 U446 ( .A(G64GAT), .B(KEYINPUT82), .Z(n394) );
  XNOR2_X1 U447 ( .A(G8GAT), .B(KEYINPUT81), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n395), .B(KEYINPUT12), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U451 ( .A(n399), .B(n398), .Z(n494) );
  INV_X1 U452 ( .A(n494), .ZN(n588) );
  XNOR2_X1 U453 ( .A(KEYINPUT36), .B(n562), .ZN(n590) );
  NAND2_X1 U454 ( .A1(n588), .A2(n590), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n400), .B(KEYINPUT66), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n401), .B(KEYINPUT45), .ZN(n402) );
  NOR2_X1 U457 ( .A1(n423), .A2(n402), .ZN(n421) );
  XOR2_X1 U458 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n404) );
  XNOR2_X1 U459 ( .A(G15GAT), .B(KEYINPUT72), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n420) );
  XOR2_X1 U461 ( .A(G113GAT), .B(G141GAT), .Z(n406) );
  XNOR2_X1 U462 ( .A(G197GAT), .B(G22GAT), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U464 ( .A(n407), .B(G50GAT), .Z(n410) );
  XNOR2_X1 U465 ( .A(n408), .B(G36GAT), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U467 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n412) );
  NAND2_X1 U468 ( .A1(G229GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U470 ( .A(n414), .B(n413), .Z(n418) );
  XNOR2_X1 U471 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n420), .B(n419), .ZN(n581) );
  INV_X1 U474 ( .A(n581), .ZN(n538) );
  NAND2_X1 U475 ( .A1(n421), .A2(n538), .ZN(n432) );
  INV_X1 U476 ( .A(KEYINPUT41), .ZN(n422) );
  XNOR2_X1 U477 ( .A(n423), .B(n422), .ZN(n573) );
  NAND2_X1 U478 ( .A1(n581), .A2(n573), .ZN(n425) );
  NAND2_X1 U479 ( .A1(n426), .A2(n494), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n427), .B(KEYINPUT115), .ZN(n428) );
  INV_X1 U481 ( .A(n562), .ZN(n466) );
  NAND2_X1 U482 ( .A1(n428), .A2(n466), .ZN(n430) );
  XOR2_X1 U483 ( .A(KEYINPUT47), .B(KEYINPUT116), .Z(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  NAND2_X1 U485 ( .A1(n432), .A2(n431), .ZN(n434) );
  NAND2_X1 U486 ( .A1(n528), .A2(n541), .ZN(n436) );
  XOR2_X1 U487 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n458) );
  XOR2_X1 U489 ( .A(KEYINPUT97), .B(G57GAT), .Z(n438) );
  XNOR2_X1 U490 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n457) );
  XOR2_X1 U492 ( .A(G85GAT), .B(G155GAT), .Z(n440) );
  XNOR2_X1 U493 ( .A(G120GAT), .B(G148GAT), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U495 ( .A(KEYINPUT96), .B(KEYINPUT6), .Z(n442) );
  XNOR2_X1 U496 ( .A(G1GAT), .B(G127GAT), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U498 ( .A(n444), .B(n443), .Z(n455) );
  XOR2_X1 U499 ( .A(n445), .B(KEYINPUT5), .Z(n447) );
  NAND2_X1 U500 ( .A1(G225GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n453) );
  XOR2_X1 U502 ( .A(n448), .B(G162GAT), .Z(n451) );
  XNOR2_X1 U503 ( .A(G29GAT), .B(n449), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U506 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U507 ( .A(n457), .B(n456), .ZN(n526) );
  INV_X1 U508 ( .A(n526), .ZN(n540) );
  NAND2_X1 U509 ( .A1(n458), .A2(n540), .ZN(n459) );
  XOR2_X1 U510 ( .A(KEYINPUT65), .B(n459), .Z(n579) );
  NOR2_X1 U511 ( .A1(n475), .A2(n579), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT55), .ZN(n567) );
  OR2_X1 U513 ( .A1(n294), .A2(n567), .ZN(n464) );
  XOR2_X1 U514 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n462) );
  XNOR2_X1 U515 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n485) );
  INV_X1 U516 ( .A(n423), .ZN(n465) );
  NAND2_X1 U517 ( .A1(n465), .A2(n581), .ZN(n499) );
  XOR2_X1 U518 ( .A(KEYINPUT16), .B(KEYINPUT83), .Z(n468) );
  NAND2_X1 U519 ( .A1(n466), .A2(n588), .ZN(n467) );
  XNOR2_X1 U520 ( .A(n468), .B(n467), .ZN(n482) );
  XOR2_X1 U521 ( .A(KEYINPUT28), .B(n475), .Z(n511) );
  INV_X1 U522 ( .A(n511), .ZN(n545) );
  XNOR2_X1 U523 ( .A(n505), .B(KEYINPUT27), .ZN(n539) );
  NOR2_X1 U524 ( .A1(n545), .A2(n539), .ZN(n469) );
  INV_X1 U525 ( .A(n532), .ZN(n568) );
  NAND2_X1 U526 ( .A1(n469), .A2(n568), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n526), .A2(n470), .ZN(n481) );
  NAND2_X1 U528 ( .A1(n528), .A2(n532), .ZN(n471) );
  XOR2_X1 U529 ( .A(KEYINPUT98), .B(n471), .Z(n472) );
  NOR2_X1 U530 ( .A1(n475), .A2(n472), .ZN(n474) );
  XNOR2_X1 U531 ( .A(KEYINPUT99), .B(KEYINPUT25), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n474), .B(n473), .ZN(n478) );
  NAND2_X1 U533 ( .A1(n475), .A2(n568), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n476), .B(KEYINPUT26), .ZN(n580) );
  NOR2_X1 U535 ( .A1(n580), .A2(n539), .ZN(n477) );
  NOR2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n479) );
  NAND2_X1 U537 ( .A1(n540), .A2(n479), .ZN(n480) );
  NAND2_X1 U538 ( .A1(n481), .A2(n480), .ZN(n496) );
  OR2_X1 U539 ( .A1(n482), .A2(n496), .ZN(n515) );
  NOR2_X1 U540 ( .A1(n499), .A2(n515), .ZN(n483) );
  XNOR2_X1 U541 ( .A(KEYINPUT100), .B(n483), .ZN(n491) );
  NAND2_X1 U542 ( .A1(n526), .A2(n491), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1324GAT) );
  XOR2_X1 U544 ( .A(G8GAT), .B(KEYINPUT101), .Z(n487) );
  NAND2_X1 U545 ( .A1(n528), .A2(n491), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(G1325GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n489) );
  NAND2_X1 U548 ( .A1(n491), .A2(n532), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(n490), .ZN(G1326GAT) );
  NAND2_X1 U551 ( .A1(n491), .A2(n545), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U553 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n503) );
  XOR2_X1 U554 ( .A(KEYINPUT104), .B(KEYINPUT37), .Z(n493) );
  XNOR2_X1 U555 ( .A(KEYINPUT103), .B(n493), .ZN(n498) );
  NAND2_X1 U556 ( .A1(n494), .A2(n590), .ZN(n495) );
  NOR2_X1 U557 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(n525) );
  NOR2_X1 U559 ( .A1(n525), .A2(n499), .ZN(n501) );
  XNOR2_X1 U560 ( .A(KEYINPUT105), .B(KEYINPUT38), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(n512) );
  NOR2_X1 U562 ( .A1(n540), .A2(n512), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(n504), .ZN(G1328GAT) );
  NOR2_X1 U565 ( .A1(n512), .A2(n505), .ZN(n507) );
  XNOR2_X1 U566 ( .A(G36GAT), .B(KEYINPUT107), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n507), .B(n506), .ZN(G1329GAT) );
  XNOR2_X1 U568 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n509) );
  NOR2_X1 U569 ( .A1(n568), .A2(n512), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U571 ( .A(G43GAT), .B(n510), .Z(G1330GAT) );
  NOR2_X1 U572 ( .A1(n512), .A2(n511), .ZN(n513) );
  XOR2_X1 U573 ( .A(G50GAT), .B(n513), .Z(G1331GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n517) );
  NAND2_X1 U575 ( .A1(n573), .A2(n538), .ZN(n514) );
  XOR2_X1 U576 ( .A(KEYINPUT109), .B(n514), .Z(n524) );
  NOR2_X1 U577 ( .A1(n515), .A2(n524), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n521), .A2(n526), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U580 ( .A(G57GAT), .B(n518), .Z(G1332GAT) );
  NAND2_X1 U581 ( .A1(n521), .A2(n528), .ZN(n519) );
  XNOR2_X1 U582 ( .A(n519), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U583 ( .A1(n532), .A2(n521), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .Z(n523) );
  NAND2_X1 U586 ( .A1(n521), .A2(n545), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  NOR2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n535), .A2(n526), .ZN(n527) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(n527), .ZN(G1336GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n530) );
  NAND2_X1 U592 ( .A1(n535), .A2(n528), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U594 ( .A(G92GAT), .B(n531), .ZN(G1337GAT) );
  XOR2_X1 U595 ( .A(G99GAT), .B(KEYINPUT113), .Z(n534) );
  NAND2_X1 U596 ( .A1(n535), .A2(n532), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n534), .B(n533), .ZN(G1338GAT) );
  NAND2_X1 U598 ( .A1(n535), .A2(n545), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n536), .B(KEYINPUT44), .ZN(n537) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n537), .ZN(G1339GAT) );
  NOR2_X1 U601 ( .A1(n540), .A2(n539), .ZN(n542) );
  NAND2_X1 U602 ( .A1(n542), .A2(n541), .ZN(n555) );
  NOR2_X1 U603 ( .A1(n568), .A2(n555), .ZN(n543) );
  XNOR2_X1 U604 ( .A(n543), .B(KEYINPUT117), .ZN(n544) );
  NOR2_X1 U605 ( .A1(n545), .A2(n544), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n581), .A2(n552), .ZN(n546) );
  XNOR2_X1 U607 ( .A(n546), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n548) );
  NAND2_X1 U609 ( .A1(n552), .A2(n573), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U611 ( .A(G120GAT), .B(n549), .ZN(G1341GAT) );
  NAND2_X1 U612 ( .A1(n588), .A2(n552), .ZN(n550) );
  XNOR2_X1 U613 ( .A(n550), .B(KEYINPUT50), .ZN(n551) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT51), .Z(n554) );
  NAND2_X1 U616 ( .A1(n552), .A2(n562), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n554), .B(n553), .ZN(G1343GAT) );
  NOR2_X1 U618 ( .A1(n580), .A2(n555), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n563), .A2(n581), .ZN(n556) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n558) );
  NAND2_X1 U622 ( .A1(n563), .A2(n573), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(n560) );
  XOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT119), .Z(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  NAND2_X1 U626 ( .A1(n588), .A2(n563), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n565) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G162GAT), .B(n566), .ZN(G1347GAT) );
  NOR2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n576) );
  NAND2_X1 U633 ( .A1(n581), .A2(n576), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n571) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT56), .B(n572), .Z(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1349GAT) );
  XOR2_X1 U641 ( .A(G183GAT), .B(KEYINPUT125), .Z(n578) );
  NAND2_X1 U642 ( .A1(n576), .A2(n588), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1350GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n583) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n591) );
  NAND2_X1 U646 ( .A1(n591), .A2(n581), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U650 ( .A1(n591), .A2(n423), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U652 ( .A(G204GAT), .B(n587), .Z(G1353GAT) );
  NAND2_X1 U653 ( .A1(n588), .A2(n591), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(n592), .B(KEYINPUT62), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

