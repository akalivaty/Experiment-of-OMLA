//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(new_n203), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n213), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT64), .Z(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n210), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n219), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n201), .A2(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n203), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n242), .B(new_n247), .ZN(G351));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  AOI22_X1  g0049(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT8), .A2(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT68), .B(G58), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n251), .B1(new_n252), .B2(KEYINPUT8), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n208), .A2(G33), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n250), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n214), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT67), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT67), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(new_n260), .A3(new_n214), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n264));
  AND3_X1   g0064(.A1(new_n259), .A2(new_n264), .A3(new_n261), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n207), .A2(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G50), .A3(new_n266), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n263), .B(new_n267), .C1(G50), .C2(new_n264), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT9), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT10), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G223), .A3(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G77), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT66), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT66), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n271), .ZN(new_n279));
  INV_X1    g0079(.A(G222), .ZN(new_n280));
  OAI221_X1 g0080(.A(new_n272), .B1(new_n273), .B2(new_n271), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  OAI211_X1 g0085(.A(G1), .B(G13), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n282), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G45), .ZN(new_n292));
  AOI21_X1  g0092(.A(G1), .B1(new_n285), .B2(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(G226), .A2(new_n289), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n283), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(G200), .B2(new_n295), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n269), .A2(new_n270), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n270), .B1(new_n269), .B2(new_n298), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n268), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(new_n295), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(G179), .B2(new_n295), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n278), .A2(new_n271), .A3(G223), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G33), .A2(G87), .ZN(new_n308));
  INV_X1    g0108(.A(G226), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n271), .A2(G1698), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n307), .B(new_n308), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n282), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n286), .A2(G274), .A3(new_n293), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n286), .A2(G232), .A3(new_n287), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(G179), .B1(new_n311), .B2(new_n282), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT73), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n313), .A2(new_n314), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n319), .B1(new_n313), .B2(new_n314), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n317), .A2(new_n303), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n284), .A2(KEYINPUT3), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT3), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G33), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OR2_X1    g0127(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n328));
  NAND2_X1  g0128(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n327), .A2(new_n208), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT7), .B1(new_n271), .B2(G20), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(new_n331), .A3(G68), .ZN(new_n332));
  INV_X1    g0132(.A(G159), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n333), .A2(G20), .A3(G33), .ZN(new_n334));
  AND2_X1   g0134(.A1(KEYINPUT68), .A2(G58), .ZN(new_n335));
  NOR2_X1   g0135(.A1(KEYINPUT68), .A2(G58), .ZN(new_n336));
  OAI21_X1  g0136(.A(G68), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n216), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n334), .B1(new_n338), .B2(G20), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n332), .A2(new_n339), .A3(KEYINPUT16), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n258), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT69), .B(KEYINPUT7), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n208), .B2(new_n327), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT71), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT70), .ZN(new_n345));
  OAI211_X1 g0145(.A(KEYINPUT7), .B(new_n208), .C1(new_n324), .C2(KEYINPUT70), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n208), .A2(KEYINPUT7), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n325), .A2(G33), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT70), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT70), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(KEYINPUT71), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n343), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n339), .B1(new_n354), .B2(new_n203), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n341), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n259), .A2(new_n264), .A3(new_n261), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n252), .A2(KEYINPUT8), .ZN(new_n359));
  INV_X1    g0159(.A(new_n251), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n360), .A3(new_n266), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n358), .B1(new_n361), .B2(KEYINPUT72), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT72), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n253), .A2(new_n363), .A3(new_n266), .ZN(new_n364));
  INV_X1    g0164(.A(new_n264), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n362), .A2(new_n364), .B1(new_n365), .B2(new_n254), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(KEYINPUT18), .B(new_n323), .C1(new_n357), .C2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT74), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n323), .B1(new_n357), .B2(new_n367), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT18), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(new_n369), .A3(new_n372), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n355), .A2(new_n356), .ZN(new_n377));
  INV_X1    g0177(.A(new_n341), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n367), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n312), .A2(new_n296), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n320), .A2(new_n321), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n315), .B1(new_n311), .B2(new_n282), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n380), .A2(new_n381), .B1(new_n382), .B2(G200), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT17), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  AOI21_X1  g0185(.A(G190), .B1(new_n311), .B2(new_n282), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n317), .A2(new_n385), .B1(new_n386), .B2(new_n322), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT17), .ZN(new_n388));
  NOR4_X1   g0188(.A1(new_n357), .A2(new_n387), .A3(new_n388), .A4(new_n367), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n376), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n365), .A2(new_n203), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT12), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n249), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n273), .B2(new_n255), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n262), .A2(new_n395), .A3(KEYINPUT11), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n365), .A2(new_n258), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(G68), .A3(new_n266), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT11), .B1(new_n262), .B2(new_n395), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n309), .B1(new_n275), .B2(new_n277), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n232), .A2(new_n274), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n271), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n286), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G238), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n313), .B1(new_n288), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT13), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n409), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT13), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT66), .B(G1698), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n413), .A2(new_n309), .B1(new_n232), .B2(new_n274), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n271), .B1(G33), .B2(G97), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n411), .B(new_n412), .C1(new_n415), .C2(new_n286), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n410), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT14), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(G169), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n410), .A2(new_n416), .A3(G179), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n418), .B1(new_n417), .B2(G169), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n402), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n417), .A2(G200), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n410), .A2(new_n416), .A3(G190), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(new_n401), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  XOR2_X1   g0227(.A(KEYINPUT8), .B(G58), .Z(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(new_n249), .B1(G20), .B2(G77), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT15), .B(G87), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n429), .B1(new_n255), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n258), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n397), .A2(G77), .A3(new_n266), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n432), .B(new_n433), .C1(G77), .C2(new_n264), .ZN(new_n434));
  INV_X1    g0234(.A(G244), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n313), .B1(new_n288), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n327), .A2(G107), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n437), .B1(new_n310), .B2(new_n408), .C1(new_n279), .C2(new_n232), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n436), .B1(new_n438), .B2(new_n282), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n434), .B1(G190), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n439), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G200), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n441), .A2(G179), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n434), .B1(new_n439), .B2(G169), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR4_X1   g0246(.A1(new_n306), .A2(new_n391), .A3(new_n427), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT21), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n292), .A2(G1), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT76), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n449), .B(new_n450), .C1(KEYINPUT5), .C2(new_n285), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n207), .B(G45), .C1(new_n285), .C2(KEYINPUT5), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT76), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n285), .A2(KEYINPUT5), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n451), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(G270), .A3(new_n286), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT77), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n454), .B(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n458), .A2(new_n291), .A3(new_n451), .A4(new_n453), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n278), .A2(new_n271), .A3(G257), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT82), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n278), .A2(new_n271), .A3(KEYINPUT82), .A4(G257), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n327), .A2(G303), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n271), .A2(G264), .A3(G1698), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n463), .A2(new_n464), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n460), .B1(new_n282), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G116), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n207), .B2(G33), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n397), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G283), .ZN(new_n472));
  INV_X1    g0272(.A(G97), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n472), .B(new_n208), .C1(G33), .C2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT20), .ZN(new_n475));
  AOI22_X1  g0275(.A1(KEYINPUT83), .A2(new_n475), .B1(new_n469), .B2(G20), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT83), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT20), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n474), .A2(new_n476), .A3(new_n478), .A4(new_n258), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n365), .A2(new_n469), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n471), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n474), .A2(new_n476), .A3(new_n258), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(new_n477), .A3(KEYINPUT20), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G169), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n448), .B1(new_n468), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n468), .A2(G179), .A3(new_n484), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n456), .A2(new_n459), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n467), .A2(new_n282), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n490), .A2(KEYINPUT21), .A3(G169), .A4(new_n484), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n486), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT84), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n385), .B1(new_n488), .B2(new_n489), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(new_n484), .ZN(new_n495));
  INV_X1    g0295(.A(new_n484), .ZN(new_n496));
  OAI211_X1 g0296(.A(KEYINPUT84), .B(new_n496), .C1(new_n468), .C2(new_n385), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n468), .A2(G190), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT85), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT85), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n495), .A2(new_n497), .A3(new_n501), .A4(new_n498), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n492), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT80), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n208), .A2(G68), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n327), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n271), .A2(KEYINPUT80), .A3(new_n208), .A4(G68), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT19), .ZN(new_n508));
  NOR2_X1   g0308(.A1(G97), .A2(G107), .ZN(new_n509));
  INV_X1    g0309(.A(G87), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n406), .A2(new_n208), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n255), .A2(KEYINPUT19), .A3(new_n473), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n506), .B(new_n507), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n258), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT81), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n430), .B(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n518), .B(new_n265), .C1(G1), .C2(new_n284), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n430), .A2(new_n365), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n516), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n278), .A2(new_n271), .A3(G238), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n324), .A2(new_n326), .A3(G244), .A4(G1698), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G116), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n282), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G179), .ZN(new_n528));
  NAND2_X1  g0328(.A1(KEYINPUT79), .A2(G250), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n449), .A2(new_n290), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(G250), .ZN(new_n531));
  OAI22_X1  g0331(.A1(KEYINPUT79), .A2(new_n531), .B1(new_n292), .B2(G1), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n286), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n527), .A2(new_n528), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n526), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n286), .B1(new_n535), .B2(new_n522), .ZN(new_n536));
  INV_X1    g0336(.A(new_n533), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n303), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n521), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(G200), .B1(new_n536), .B2(new_n537), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n527), .A2(G190), .A3(new_n533), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n515), .A2(new_n258), .B1(new_n365), .B2(new_n430), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n265), .B(G87), .C1(G1), .C2(new_n284), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n540), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n324), .A2(new_n326), .A3(G250), .A4(G1698), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n472), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT4), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n278), .A2(new_n271), .A3(G244), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n278), .A2(new_n271), .A3(KEYINPUT4), .A4(G244), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n286), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n455), .A2(G257), .A3(new_n286), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n459), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n303), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n553), .A2(new_n459), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n549), .A2(new_n548), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n557), .A2(new_n472), .A3(new_n551), .A4(new_n546), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n282), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n556), .A2(new_n559), .A3(new_n528), .ZN(new_n560));
  INV_X1    g0360(.A(new_n343), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n351), .A2(KEYINPUT71), .A3(new_n352), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT71), .B1(new_n351), .B2(new_n352), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G107), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n249), .A2(G77), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n566), .B(KEYINPUT75), .ZN(new_n567));
  INV_X1    g0367(.A(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(KEYINPUT6), .A3(G97), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n473), .A2(new_n568), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(new_n509), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n571), .B2(KEYINPUT6), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n567), .B1(G20), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n565), .A2(new_n573), .B1(new_n214), .B2(new_n257), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n365), .A2(new_n473), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n265), .B1(G1), .B2(new_n284), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n575), .B1(new_n576), .B2(new_n473), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n555), .B(new_n560), .C1(new_n574), .C2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(G200), .B1(new_n552), .B2(new_n554), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n552), .A2(new_n554), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n579), .A2(KEYINPUT78), .B1(new_n580), .B2(G190), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n573), .B1(new_n354), .B2(new_n568), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n577), .B1(new_n582), .B2(new_n258), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n556), .A2(new_n559), .A3(KEYINPUT78), .A4(G190), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n545), .B(new_n578), .C1(new_n581), .C2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n279), .A2(new_n531), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n271), .A2(G257), .A3(G1698), .ZN(new_n588));
  INV_X1    g0388(.A(G294), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n589), .A2(KEYINPUT88), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(KEYINPUT88), .ZN(new_n591));
  OAI21_X1  g0391(.A(G33), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n282), .B1(new_n587), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n455), .A2(G264), .A3(new_n286), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n459), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(G190), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n595), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT89), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT89), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n594), .A2(new_n600), .A3(new_n595), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n459), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n597), .B1(new_n602), .B2(new_n385), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n264), .A2(G107), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n604), .B(KEYINPUT25), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n576), .B2(new_n568), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n208), .A2(KEYINPUT86), .A3(G87), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n271), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT22), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n271), .A2(new_n607), .A3(KEYINPUT22), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT23), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(new_n568), .A3(G20), .ZN(new_n615));
  NAND2_X1  g0415(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n612), .A2(new_n613), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n610), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  OR2_X1    g0418(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n618), .B(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n606), .B1(new_n620), .B2(new_n258), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n603), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n599), .A2(G179), .A3(new_n459), .A4(new_n601), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n596), .A2(G169), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n586), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n447), .A2(new_n503), .A3(new_n627), .ZN(G372));
  NOR2_X1   g0428(.A1(new_n626), .A2(new_n492), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n629), .A2(new_n586), .A3(new_n623), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n552), .A2(G179), .A3(new_n554), .ZN(new_n631));
  AOI21_X1  g0431(.A(G169), .B1(new_n556), .B2(new_n559), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n583), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(KEYINPUT26), .A3(new_n545), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n539), .A2(new_n544), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n635), .B1(new_n578), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n539), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n447), .B1(new_n630), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n305), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n373), .A2(new_n368), .ZN(new_n642));
  INV_X1    g0442(.A(new_n423), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n445), .A2(new_n444), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n426), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n564), .A2(G68), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT16), .B1(new_n646), .B2(new_n339), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n383), .B(new_n366), .C1(new_n647), .C2(new_n341), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n388), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n379), .A2(KEYINPUT17), .A3(new_n383), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n642), .B1(new_n645), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n641), .B1(new_n652), .B2(new_n301), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n640), .A2(new_n653), .ZN(G369));
  XNOR2_X1  g0454(.A(KEYINPUT93), .B(G330), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT90), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT90), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n657), .A2(new_n661), .A3(new_n658), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n660), .A2(new_n662), .A3(G213), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT91), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n660), .A2(new_n662), .A3(new_n665), .A4(G213), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n484), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT92), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT92), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n503), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n492), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n655), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n602), .A2(new_n385), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n621), .B1(new_n677), .B2(new_n597), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n624), .A2(new_n625), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n622), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n622), .A2(new_n669), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n678), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n626), .A2(new_n669), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n676), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n623), .A2(new_n626), .ZN(new_n686));
  INV_X1    g0486(.A(new_n669), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n492), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n686), .A2(new_n689), .B1(new_n626), .B2(new_n687), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n685), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n211), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n511), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n217), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT94), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n536), .A2(new_n537), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n580), .A2(new_n599), .A3(new_n601), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n468), .A2(G179), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n599), .A2(new_n601), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n490), .A2(new_n528), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n701), .A2(new_n556), .A3(new_n559), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n705), .A2(new_n706), .A3(KEYINPUT30), .A4(new_n707), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n580), .A2(G179), .A3(new_n701), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(new_n490), .A3(new_n602), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n704), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT31), .B1(new_n711), .B2(new_n669), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT95), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n669), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT31), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT95), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(new_n719), .A3(new_n712), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n627), .A2(new_n503), .A3(new_n687), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n715), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n655), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n486), .A2(new_n487), .A3(new_n491), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n680), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n582), .A2(new_n258), .ZN(new_n727));
  INV_X1    g0527(.A(new_n577), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n584), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n579), .A2(KEYINPUT78), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n580), .A2(G190), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n631), .A2(new_n632), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n727), .A2(new_n728), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n729), .A2(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n726), .A2(new_n678), .A3(new_n735), .A4(new_n545), .ZN(new_n736));
  INV_X1    g0536(.A(new_n539), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(new_n634), .B2(new_n637), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n669), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT29), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n724), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n699), .B1(new_n742), .B2(G1), .ZN(G364));
  AND2_X1   g0543(.A1(new_n208), .A2(G13), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G45), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT96), .Z(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n747), .A2(new_n207), .A3(new_n693), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n676), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n673), .A2(new_n675), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n749), .B1(new_n723), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G13), .A2(G33), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n214), .B1(G20), .B2(new_n303), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n247), .A2(new_n292), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n692), .A2(new_n271), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n758), .B(new_n760), .C1(new_n292), .C2(new_n218), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT97), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n211), .A2(new_n271), .ZN(new_n763));
  INV_X1    g0563(.A(G355), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n763), .A2(new_n764), .B1(G116), .B2(new_n211), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n761), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n765), .A2(new_n762), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n757), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n748), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n208), .A2(new_n528), .A3(new_n296), .A4(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G322), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n208), .A2(new_n528), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G190), .A2(G200), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n327), .B1(new_n771), .B2(new_n772), .C1(new_n773), .C2(new_n777), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n590), .A2(new_n591), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n296), .A2(G179), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n208), .ZN(new_n782));
  INV_X1    g0582(.A(G326), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n774), .A2(G190), .A3(G200), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n780), .A2(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n208), .A2(new_n385), .A3(G179), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G190), .ZN(new_n787));
  INV_X1    g0587(.A(G303), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n774), .A2(new_n296), .A3(G200), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT33), .B(G317), .Z(new_n790));
  OAI22_X1  g0590(.A1(new_n787), .A2(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n778), .A2(new_n785), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n775), .A2(G20), .A3(new_n528), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT98), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(KEYINPUT98), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n786), .A2(new_n296), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n797), .A2(G329), .B1(G283), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n800), .A2(KEYINPUT99), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(KEYINPUT99), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n792), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT100), .ZN(new_n804));
  INV_X1    g0604(.A(new_n793), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G159), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n806), .A2(KEYINPUT32), .B1(new_n787), .B2(new_n510), .ZN(new_n807));
  INV_X1    g0607(.A(new_n789), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(G68), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n271), .B1(new_n777), .B2(new_n273), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(new_n252), .B2(new_n770), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G107), .A2(new_n799), .B1(new_n806), .B2(KEYINPUT32), .ZN(new_n812));
  INV_X1    g0612(.A(new_n782), .ZN(new_n813));
  INV_X1    g0613(.A(new_n784), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G97), .A2(new_n813), .B1(new_n814), .B2(G50), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n809), .A2(new_n811), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n803), .A2(KEYINPUT100), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n804), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n768), .B(new_n769), .C1(new_n818), .C2(new_n755), .ZN(new_n819));
  INV_X1    g0619(.A(new_n754), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n750), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n751), .A2(new_n821), .ZN(G396));
  NAND2_X1  g0622(.A1(new_n644), .A2(new_n687), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n440), .A2(new_n442), .B1(new_n669), .B2(new_n434), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n644), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n739), .B(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n748), .B1(new_n724), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n724), .B2(new_n827), .ZN(new_n829));
  INV_X1    g0629(.A(new_n755), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G159), .A2(new_n776), .B1(new_n770), .B2(G143), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  INV_X1    g0632(.A(G150), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n831), .B1(new_n832), .B2(new_n784), .C1(new_n833), .C2(new_n789), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT34), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n797), .A2(G132), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n201), .A2(new_n787), .B1(new_n798), .B2(new_n203), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n327), .B(new_n839), .C1(new_n252), .C2(new_n813), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n327), .B1(new_n771), .B2(new_n589), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G116), .B2(new_n776), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n510), .A2(new_n798), .B1(new_n787), .B2(new_n568), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G283), .B2(new_n808), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n797), .A2(G311), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G97), .A2(new_n813), .B1(new_n814), .B2(G303), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n843), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n830), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n755), .A2(new_n752), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT101), .Z(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n769), .B(new_n849), .C1(new_n273), .C2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n826), .B2(new_n753), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n829), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G384));
  OR2_X1    g0656(.A1(new_n572), .A2(KEYINPUT35), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n572), .A2(KEYINPUT35), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n857), .A2(G116), .A3(new_n215), .A4(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT36), .Z(new_n860));
  NAND3_X1  g0660(.A1(new_n218), .A2(G77), .A3(new_n337), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n207), .B(G13), .C1(new_n861), .C2(new_n243), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT29), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n739), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n447), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n653), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT105), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n340), .A2(new_n262), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT16), .B1(new_n332), .B2(new_n339), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n366), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT104), .ZN(new_n872));
  INV_X1    g0672(.A(new_n667), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT104), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n366), .B(new_n874), .C1(new_n869), .C2(new_n870), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n872), .A2(new_n323), .A3(new_n875), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n648), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n873), .B1(new_n357), .B2(new_n367), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n371), .A2(new_n880), .A3(new_n648), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n651), .B1(new_n374), .B2(new_n375), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n883), .B(KEYINPUT38), .C1(new_n884), .C2(new_n876), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n371), .A2(new_n880), .A3(new_n648), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(new_n881), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n880), .B1(new_n390), .B2(new_n642), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT39), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n876), .B1(new_n376), .B2(new_n390), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n879), .A2(new_n882), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n886), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n643), .A2(new_n687), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n893), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n642), .A2(new_n873), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n896), .A2(new_n885), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n669), .A2(new_n402), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n423), .A2(new_n426), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n417), .A2(G169), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT14), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n426), .A2(new_n906), .A3(new_n420), .A4(new_n419), .ZN(new_n907));
  INV_X1    g0707(.A(new_n903), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(KEYINPUT103), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT103), .B1(new_n907), .B2(new_n908), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n687), .B(new_n826), .C1(new_n630), .C2(new_n639), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n823), .B(KEYINPUT102), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n912), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n901), .B1(new_n902), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n900), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n868), .B(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n826), .B1(new_n910), .B2(new_n911), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n713), .A2(new_n714), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(new_n721), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT106), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n923), .A2(KEYINPUT40), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n922), .A2(new_n924), .B1(new_n885), .B2(new_n896), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n921), .A2(new_n721), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT106), .B1(new_n926), .B2(new_n920), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n922), .A2(new_n891), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n925), .A2(new_n927), .B1(KEYINPUT40), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n921), .A2(new_n721), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n447), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n932), .A2(new_n655), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n919), .A2(new_n933), .B1(new_n207), .B2(new_n744), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n919), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n863), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT107), .Z(G367));
  OAI221_X1 g0737(.A(new_n756), .B1(new_n211), .B2(new_n430), .C1(new_n760), .C2(new_n238), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT112), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n769), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n939), .B2(new_n938), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n789), .A2(new_n333), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n798), .A2(new_n273), .ZN(new_n943));
  INV_X1    g0743(.A(new_n787), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n942), .B(new_n943), .C1(new_n252), .C2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n327), .B1(new_n805), .B2(G137), .ZN(new_n946));
  AOI22_X1  g0746(.A1(G50), .A2(new_n776), .B1(new_n770), .B2(G150), .ZN(new_n947));
  AOI22_X1  g0747(.A1(G68), .A2(new_n813), .B1(new_n814), .B2(G143), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n945), .A2(new_n946), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n798), .A2(new_n473), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n271), .B(new_n950), .C1(G317), .C2(new_n805), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT113), .ZN(new_n952));
  INV_X1    g0752(.A(G283), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n953), .A2(new_n777), .B1(new_n771), .B2(new_n788), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(G107), .B2(new_n813), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n779), .A2(new_n808), .B1(new_n814), .B2(G311), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT46), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n787), .B2(new_n469), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n944), .A2(KEYINPUT46), .A3(G116), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n955), .A2(new_n956), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n949), .B1(new_n952), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT47), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n941), .B1(new_n962), .B2(new_n755), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n542), .A2(new_n543), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n669), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n545), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n539), .B2(new_n965), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n963), .B1(new_n967), .B2(new_n820), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n747), .A2(new_n207), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT44), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n669), .A2(new_n734), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n735), .A2(KEYINPUT108), .A3(new_n972), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n972), .B(new_n578), .C1(new_n581), .C2(new_n585), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT108), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n633), .A2(new_n669), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n973), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n971), .B1(new_n690), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n690), .A2(new_n978), .A3(new_n971), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n690), .A2(new_n978), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT45), .B1(new_n690), .B2(new_n978), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n980), .A2(new_n981), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n685), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n982), .B(new_n983), .ZN(new_n989));
  OR3_X1    g0789(.A1(new_n690), .A2(new_n978), .A3(new_n971), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n979), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(new_n991), .A3(new_n685), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n676), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n682), .A2(new_n683), .A3(new_n688), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT110), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n686), .A2(new_n689), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n682), .A2(new_n683), .A3(KEYINPUT110), .A4(new_n688), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n994), .A2(new_n1000), .A3(KEYINPUT111), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n999), .A2(new_n998), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT111), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1002), .B(new_n997), .C1(new_n676), .C2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n742), .B1(new_n993), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n693), .B(KEYINPUT41), .Z(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n970), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n978), .A2(new_n686), .A3(new_n689), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1010), .A2(KEYINPUT42), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n973), .A2(new_n976), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n578), .B1(new_n1012), .B2(new_n680), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n687), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1010), .A2(KEYINPUT42), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1011), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n750), .A2(new_n723), .A3(new_n684), .A4(new_n978), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT109), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT109), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n676), .A2(new_n1023), .A3(new_n684), .A4(new_n978), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1020), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1022), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1018), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n1021), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1030), .A2(new_n1017), .A3(new_n1016), .A4(new_n1025), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n968), .B1(new_n1009), .B2(new_n1032), .ZN(G387));
  NAND2_X1  g0833(.A1(new_n1005), .A2(new_n741), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1001), .A2(new_n1004), .A3(new_n724), .A4(new_n740), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1034), .A2(new_n693), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1001), .A2(new_n1004), .A3(new_n970), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n763), .A2(new_n695), .B1(G107), .B2(new_n211), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n235), .A2(new_n292), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n428), .A2(new_n201), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT50), .Z(new_n1041));
  INV_X1    g0841(.A(new_n695), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n1042), .C1(G68), .C2(G77), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n760), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1038), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n748), .B1(new_n1045), .B2(new_n757), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G303), .A2(new_n776), .B1(new_n770), .B2(G317), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n773), .B2(new_n789), .C1(new_n772), .C2(new_n784), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n944), .A2(new_n779), .B1(new_n813), .B2(G283), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT114), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT49), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n327), .B1(new_n783), .B2(new_n793), .C1(new_n798), .C2(new_n469), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT115), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n950), .B1(G77), .B2(new_n944), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n333), .B2(new_n784), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n771), .A2(new_n201), .B1(new_n793), .B2(new_n833), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n327), .B(new_n1062), .C1(G68), .C2(new_n776), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n518), .A2(new_n813), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n253), .A2(new_n808), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1056), .A2(new_n1059), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1046), .B1(new_n1067), .B2(new_n755), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n684), .B2(new_n820), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1037), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1036), .A2(new_n1070), .ZN(G393));
  OAI221_X1 g0871(.A(new_n756), .B1(new_n473), .B2(new_n211), .C1(new_n760), .C2(new_n242), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n748), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n327), .B1(new_n772), .B2(new_n793), .C1(new_n798), .C2(new_n568), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G283), .B2(new_n944), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT116), .Z(new_n1076));
  AOI22_X1  g0876(.A1(new_n814), .A2(G317), .B1(new_n770), .B2(G311), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT52), .Z(new_n1078));
  NAND2_X1  g0878(.A1(new_n808), .A2(G303), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n813), .A2(G116), .B1(G294), .B2(new_n776), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT117), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n771), .A2(new_n333), .B1(new_n784), .B2(new_n833), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT51), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n805), .A2(G143), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n327), .B(new_n1086), .C1(new_n428), .C2(new_n776), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n782), .A2(new_n273), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n798), .A2(new_n510), .B1(new_n789), .B2(new_n201), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(G68), .C2(new_n944), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1085), .A2(new_n1087), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1083), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1073), .B1(new_n1093), .B2(new_n755), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n820), .B2(new_n978), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n993), .B2(new_n969), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1035), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(new_n992), .A3(new_n988), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1098), .A2(new_n693), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n993), .A2(new_n1035), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(G390));
  NAND2_X1  g0902(.A1(new_n893), .A2(new_n897), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n914), .B1(new_n739), .B2(new_n826), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n898), .B1(new_n1104), .B2(new_n912), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n913), .A2(new_n915), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT118), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n910), .B2(new_n911), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n911), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1109), .A2(KEYINPUT118), .A3(new_n904), .A4(new_n909), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n899), .B1(new_n885), .B2(new_n890), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1103), .A2(new_n1105), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n912), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n722), .A2(new_n723), .A3(new_n826), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(KEYINPUT119), .ZN(new_n1118));
  INV_X1    g0918(.A(G330), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n926), .A2(new_n1119), .A3(new_n920), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1106), .A2(new_n1115), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n893), .A2(new_n897), .B1(new_n1121), .B2(new_n898), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1120), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT119), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1126), .A2(new_n1127), .A3(new_n1123), .A4(new_n1116), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1118), .A2(new_n1125), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n912), .B1(new_n724), .B2(new_n825), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n926), .A2(new_n1119), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n920), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n1106), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n930), .A2(G330), .A3(new_n826), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1111), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1106), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n1116), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1131), .A2(new_n447), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1141), .A2(new_n866), .A3(new_n653), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1129), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1142), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1146), .A2(new_n1118), .A3(new_n1125), .A4(new_n1128), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1145), .A2(new_n693), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1128), .A2(new_n1125), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1127), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n970), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1103), .A2(new_n752), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n769), .B1(new_n852), .B2(new_n254), .ZN(new_n1154));
  INV_X1    g0954(.A(G128), .ZN(new_n1155));
  INV_X1    g0955(.A(G132), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n271), .B1(new_n1155), .B2(new_n784), .C1(new_n771), .C2(new_n1156), .ZN(new_n1157));
  OR3_X1    g0957(.A1(new_n787), .A2(KEYINPUT53), .A3(new_n833), .ZN(new_n1158));
  OAI21_X1  g0958(.A(KEYINPUT53), .B1(new_n787), .B2(new_n833), .ZN(new_n1159));
  INV_X1    g0959(.A(G125), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1158), .B(new_n1159), .C1(new_n1160), .C2(new_n796), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1157), .B(new_n1161), .C1(G50), .C2(new_n799), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT54), .B(G143), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n813), .A2(G159), .B1(new_n776), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n832), .B2(new_n789), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT120), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n203), .A2(new_n798), .B1(new_n787), .B2(new_n510), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n327), .B1(new_n771), .B2(new_n469), .C1(new_n473), .C2(new_n777), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(G294), .C2(new_n797), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n789), .A2(new_n568), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1171), .B(new_n1088), .C1(G283), .C2(new_n814), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1162), .A2(new_n1167), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1153), .B(new_n1154), .C1(new_n830), .C2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1148), .A2(new_n1152), .A3(new_n1174), .ZN(G378));
  NAND2_X1  g0975(.A1(new_n873), .A2(new_n268), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n306), .B(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n930), .A2(new_n1132), .A3(new_n924), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1180), .B(new_n902), .C1(new_n922), .C2(new_n923), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n928), .A2(KEYINPUT40), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n900), .A2(new_n917), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1183), .A2(new_n1184), .A3(G330), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1184), .B1(new_n1183), .B2(G330), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1179), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n918), .B1(new_n929), .B2(new_n1119), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1179), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1183), .A2(new_n1184), .A3(G330), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n970), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n769), .B1(new_n201), .B2(new_n850), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT121), .Z(new_n1195));
  OAI22_X1  g0995(.A1(new_n1160), .A2(new_n784), .B1(new_n789), .B2(new_n1156), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G137), .A2(new_n776), .B1(new_n770), .B2(G128), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n787), .B2(new_n1163), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(G150), .C2(new_n813), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n799), .A2(G159), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G33), .B(G41), .C1(new_n805), .C2(G124), .ZN(new_n1204));
  AND4_X1   g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n271), .A2(G41), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n203), .B2(new_n782), .C1(new_n771), .C2(new_n568), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G283), .B2(new_n797), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n784), .A2(new_n469), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n787), .A2(new_n273), .B1(new_n789), .B2(new_n473), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(new_n252), .C2(new_n799), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n518), .A2(new_n776), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1208), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT58), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AOI211_X1 g1015(.A(G50), .B(new_n1206), .C1(new_n284), .C2(new_n285), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(new_n1205), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1195), .B1(new_n830), .B2(new_n1218), .C1(new_n1179), .C2(new_n753), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT122), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1193), .A2(new_n1220), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1189), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1223));
  OAI21_X1  g1023(.A(KEYINPUT57), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT123), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1142), .B(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1151), .B2(new_n1146), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT124), .B1(new_n1224), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1226), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1129), .B2(new_n1144), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT124), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1230), .A2(new_n1231), .A3(KEYINPUT57), .A4(new_n1192), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1228), .A2(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1147), .A2(new_n1229), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n693), .B1(new_n1234), .B2(KEYINPUT57), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1221), .B1(new_n1233), .B2(new_n1235), .ZN(G375));
  AOI22_X1  g1036(.A1(new_n1134), .A2(new_n1106), .B1(new_n1116), .B2(new_n1138), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1142), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1144), .A2(new_n1008), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1137), .A2(new_n752), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n787), .A2(new_n473), .B1(new_n784), .B2(new_n589), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n943), .B(new_n1241), .C1(G116), .C2(new_n808), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n797), .A2(G303), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n327), .B1(new_n771), .B2(new_n953), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G107), .B2(new_n776), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1242), .A2(new_n1064), .A3(new_n1243), .A4(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n271), .B1(new_n771), .B2(new_n832), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G150), .B2(new_n776), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n787), .A2(new_n333), .B1(new_n784), .B2(new_n1156), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n808), .B2(new_n1164), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n797), .A2(G128), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n799), .A2(new_n252), .B1(new_n813), .B2(G50), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1248), .A2(new_n1250), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n830), .B1(new_n1246), .B2(new_n1253), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n769), .B(new_n1254), .C1(new_n203), .C2(new_n852), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1140), .A2(new_n970), .B1(new_n1240), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1239), .A2(new_n1256), .ZN(G381));
  OR2_X1    g1057(.A1(G375), .A2(KEYINPUT125), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G375), .A2(KEYINPUT125), .ZN(new_n1259));
  INV_X1    g1059(.A(G396), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1036), .A2(new_n1260), .A3(new_n1070), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1101), .A2(new_n855), .A3(new_n1262), .ZN(new_n1263));
  NOR4_X1   g1063(.A1(G378), .A2(G387), .A3(G381), .A4(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1258), .A2(new_n1259), .A3(new_n1264), .ZN(G407));
  INV_X1    g1065(.A(G378), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n668), .A2(G213), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1258), .A2(new_n1266), .A3(new_n1259), .A4(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1269), .A2(G213), .A3(G407), .ZN(G409));
  OAI211_X1 g1070(.A(G378), .B(new_n1221), .C1(new_n1233), .C2(new_n1235), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1234), .A2(new_n1008), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1193), .A2(new_n1219), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1266), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1267), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1238), .B1(new_n1146), .B2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1237), .A2(KEYINPUT60), .A3(new_n1142), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n693), .A3(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(G384), .A3(new_n1256), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(G384), .B1(new_n1280), .B2(new_n1256), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1268), .A2(G2897), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G2897), .B(new_n1268), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT61), .B1(new_n1276), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1280), .A2(new_n1256), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n855), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1281), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1290), .B1(new_n1276), .B2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1260), .B1(new_n1036), .B2(new_n1070), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1262), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(G387), .B2(KEYINPUT126), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G393), .A2(G396), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1261), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1007), .B1(new_n1098), .B2(new_n742), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1300), .B1(new_n1301), .B2(new_n970), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1299), .B1(new_n1302), .B2(new_n968), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1101), .B1(new_n1297), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(G387), .A2(new_n1296), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT126), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(new_n1302), .B2(new_n968), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G390), .B(new_n1305), .C1(new_n1307), .C2(new_n1296), .ZN(new_n1308));
  AND2_X1   g1108(.A1(new_n1304), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1268), .B1(new_n1271), .B2(new_n1274), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1311), .A2(KEYINPUT63), .A3(new_n1284), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1289), .A2(new_n1294), .A3(new_n1310), .A4(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1311), .A2(new_n1314), .A3(new_n1284), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1316), .B1(new_n1311), .B2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1314), .B1(new_n1311), .B2(new_n1284), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1315), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1313), .B1(new_n1320), .B2(new_n1310), .ZN(G405));
  INV_X1    g1121(.A(KEYINPUT127), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1309), .A2(new_n1271), .A3(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1309), .B1(new_n1322), .B2(new_n1271), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1284), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  AND2_X1   g1125(.A1(G375), .A2(new_n1266), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1271), .A2(new_n1322), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1310), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1309), .A2(new_n1271), .A3(new_n1322), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1328), .A2(new_n1293), .A3(new_n1329), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1325), .A2(new_n1326), .A3(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1326), .B1(new_n1325), .B2(new_n1330), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1332), .ZN(G402));
endmodule


