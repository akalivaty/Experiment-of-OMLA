//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  NAND3_X1  g001(.A1(new_n202), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT14), .B(G29gat), .Z(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(G43gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G50gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT89), .B(G50gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(new_n206), .ZN(new_n209));
  XOR2_X1   g008(.A(KEYINPUT88), .B(KEYINPUT15), .Z(new_n210));
  OAI21_X1  g009(.A(new_n205), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n206), .A2(G50gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(KEYINPUT15), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n205), .A2(KEYINPUT15), .A3(new_n213), .A4(new_n212), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT17), .ZN(new_n218));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n220), .B2(G1gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G1gat), .B2(new_n219), .ZN(new_n222));
  INV_X1    g021(.A(G8gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT90), .B(KEYINPUT17), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n215), .A2(new_n216), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n218), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n217), .ZN(new_n229));
  INV_X1    g028(.A(new_n224), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT18), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n227), .A2(KEYINPUT18), .A3(new_n228), .A4(new_n231), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n217), .B(new_n224), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n228), .B(KEYINPUT13), .Z(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n234), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G113gat), .B(G141gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(G197gat), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT11), .B(G169gat), .Z(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT12), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n232), .A2(new_n233), .B1(new_n236), .B2(new_n237), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(new_n244), .A3(new_n235), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AND2_X1   g049(.A1(G232gat), .A2(G233gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(KEYINPUT41), .ZN(new_n252));
  XNOR2_X1  g051(.A(G134gat), .B(G162gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G85gat), .A2(G92gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT7), .ZN(new_n257));
  XNOR2_X1  g056(.A(G99gat), .B(G106gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(G85gat), .A2(G92gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(G99gat), .A2(G106gat), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n259), .B1(KEYINPUT8), .B2(new_n260), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n257), .A2(new_n258), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n258), .B1(new_n257), .B2(new_n261), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT93), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n263), .A2(KEYINPUT93), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n229), .A2(new_n267), .B1(KEYINPUT41), .B2(new_n251), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n218), .A2(new_n226), .A3(new_n266), .ZN(new_n269));
  XOR2_X1   g068(.A(G190gat), .B(G218gat), .Z(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n268), .B2(new_n269), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n255), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n274), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(new_n254), .A3(new_n272), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  OR2_X1    g077(.A1(G57gat), .A2(G64gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(G57gat), .A2(G64gat), .ZN(new_n280));
  AND2_X1   g079(.A1(G71gat), .A2(G78gat), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n279), .B(new_n280), .C1(new_n281), .C2(KEYINPUT9), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(KEYINPUT91), .B2(new_n281), .ZN(new_n283));
  NOR2_X1   g082(.A1(G71gat), .A2(G78gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n283), .B(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n230), .B1(KEYINPUT21), .B2(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n283), .B(new_n285), .Z(new_n288));
  INV_X1    g087(.A(G231gat), .ZN(new_n289));
  INV_X1    g088(.A(G233gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n288), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n292), .B1(new_n288), .B2(new_n293), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n295), .A2(G127gat), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G127gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n288), .A2(new_n293), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(new_n291), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n298), .B1(new_n300), .B2(new_n294), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n287), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(G127gat), .B1(new_n295), .B2(new_n296), .ZN(new_n303));
  INV_X1    g102(.A(new_n287), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(new_n298), .A3(new_n294), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n307));
  INV_X1    g106(.A(G155gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G183gat), .B(G211gat), .ZN(new_n310));
  XOR2_X1   g109(.A(new_n309), .B(new_n310), .Z(new_n311));
  NAND3_X1  g110(.A1(new_n302), .A2(new_n306), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n302), .B2(new_n306), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n278), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT94), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n302), .A2(new_n306), .ZN(new_n317));
  INV_X1    g116(.A(new_n311), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n312), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT94), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(new_n278), .ZN(new_n322));
  INV_X1    g121(.A(G230gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(new_n290), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT10), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n262), .A2(new_n263), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n286), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n325), .B(new_n327), .C1(new_n267), .C2(new_n286), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n267), .A2(KEYINPUT10), .A3(new_n286), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n286), .B1(new_n264), .B2(new_n265), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n286), .A2(new_n326), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n324), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G120gat), .B(G148gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(KEYINPUT95), .ZN(new_n337));
  XNOR2_X1  g136(.A(G176gat), .B(G204gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  NOR3_X1   g138(.A1(new_n330), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n330), .B2(new_n335), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n316), .A2(new_n322), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G148gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT74), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G148gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n349), .A3(G141gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n346), .A2(G141gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT2), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G162gat), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n356), .B1(new_n308), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G141gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(G148gat), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n355), .B1(new_n351), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(new_n354), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n353), .A2(new_n358), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(G211gat), .A2(G218gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(G211gat), .A2(G218gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G197gat), .ZN(new_n372));
  INV_X1    g171(.A(G204gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(G197gat), .A2(G204gat), .ZN(new_n375));
  OAI22_X1  g174(.A1(new_n374), .A2(new_n375), .B1(KEYINPUT22), .B2(new_n369), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n371), .B1(new_n377), .B2(KEYINPUT70), .ZN(new_n378));
  INV_X1    g177(.A(new_n371), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT70), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n376), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n368), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G228gat), .A2(G233gat), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G141gat), .B(G148gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n363), .B1(new_n386), .B2(KEYINPUT2), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT74), .B(G148gat), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n351), .B1(new_n388), .B2(G141gat), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n362), .B1(new_n355), .B2(new_n354), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n387), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n377), .A2(new_n371), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT29), .B1(new_n376), .B2(new_n379), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(KEYINPUT82), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n365), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT82), .B1(new_n392), .B2(new_n393), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n385), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n378), .A2(new_n367), .A3(new_n381), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT83), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n378), .A2(KEYINPUT83), .A3(new_n367), .A4(new_n381), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n365), .A3(new_n402), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n403), .A2(new_n391), .B1(new_n382), .B2(new_n368), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n398), .B1(new_n404), .B2(new_n384), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT31), .B(G50gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(G78gat), .B(G106gat), .Z(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(KEYINPUT81), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(G22gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n406), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n398), .B(new_n411), .C1(new_n404), .C2(new_n384), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n407), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n410), .B1(new_n407), .B2(new_n412), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n416));
  INV_X1    g215(.A(G120gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G113gat), .ZN(new_n418));
  INV_X1    g217(.A(G113gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G120gat), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT1), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n298), .A2(G134gat), .ZN(new_n422));
  INV_X1    g221(.A(G134gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(G127gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT69), .B1(new_n298), .B2(G134gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n422), .A2(new_n424), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n426), .B1(new_n427), .B2(KEYINPUT69), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n425), .B1(new_n428), .B2(new_n421), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT75), .B1(new_n429), .B2(new_n391), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT75), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT69), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n432), .B1(new_n422), .B2(new_n424), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n418), .A2(new_n420), .ZN(new_n434));
  OAI22_X1  g233(.A1(new_n426), .A2(new_n433), .B1(new_n434), .B2(KEYINPUT1), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n364), .A2(new_n431), .A3(new_n435), .A4(new_n425), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT76), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT4), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n391), .A2(KEYINPUT3), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n366), .A2(new_n441), .A3(new_n429), .ZN(new_n442));
  NAND2_X1  g241(.A1(G225gat), .A2(G233gat), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT4), .B1(new_n430), .B2(new_n436), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n391), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT76), .B1(new_n446), .B2(new_n439), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n440), .B(new_n444), .C1(new_n445), .C2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT77), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n429), .A2(new_n391), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n430), .A2(new_n436), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n443), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n449), .B1(new_n453), .B2(KEYINPUT5), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT5), .ZN(new_n455));
  AOI211_X1 g254(.A(KEYINPUT77), .B(new_n455), .C1(new_n451), .C2(new_n452), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n448), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G1gat), .B(G29gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT0), .ZN(new_n459));
  XNOR2_X1  g258(.A(G57gat), .B(G85gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n446), .A2(KEYINPUT4), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n462), .B1(KEYINPUT4), .B2(new_n437), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n442), .A2(new_n455), .A3(new_n443), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n457), .A2(KEYINPUT78), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n461), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n463), .A2(new_n464), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(new_n457), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n416), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT78), .B1(new_n457), .B2(new_n465), .ZN(new_n471));
  INV_X1    g270(.A(new_n416), .ZN(new_n472));
  INV_X1    g271(.A(new_n468), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n453), .A2(KEYINPUT5), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT77), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n453), .A2(new_n449), .A3(KEYINPUT5), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n473), .B1(new_n477), .B2(new_n448), .ZN(new_n478));
  OAI22_X1  g277(.A1(new_n471), .A2(new_n472), .B1(new_n478), .B2(new_n467), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n470), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G183gat), .A2(G190gat), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n482));
  AND2_X1   g281(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(G190gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G169gat), .A2(G176gat), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT25), .B1(new_n486), .B2(KEYINPUT65), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n487), .B1(KEYINPUT65), .B2(new_n486), .ZN(new_n488));
  INV_X1    g287(.A(G169gat), .ZN(new_n489));
  INV_X1    g288(.A(G176gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT23), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT23), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(G169gat), .B2(G176gat), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n485), .A2(new_n488), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(new_n493), .A3(new_n486), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n496), .B1(new_n484), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT64), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT64), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n500), .B(new_n496), .C1(new_n484), .C2(new_n497), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n495), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G183gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT27), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT27), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G183gat), .ZN(new_n506));
  INV_X1    g305(.A(G190gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT66), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT28), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT28), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT67), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT26), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT26), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n517), .A2(new_n489), .A3(new_n490), .A4(KEYINPUT67), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n486), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n481), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT68), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(KEYINPUT68), .A3(new_n481), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n514), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G226gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(new_n290), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n502), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(KEYINPUT29), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n499), .A2(new_n501), .ZN(new_n529));
  INV_X1    g328(.A(new_n495), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n512), .A2(new_n513), .ZN(new_n532));
  INV_X1    g331(.A(new_n523), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT68), .B1(new_n519), .B2(new_n481), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n528), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n382), .B1(new_n527), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n531), .B(new_n535), .C1(new_n525), .C2(new_n290), .ZN(new_n538));
  OAI22_X1  g337(.A1(new_n502), .A2(new_n524), .B1(KEYINPUT29), .B2(new_n526), .ZN(new_n539));
  INV_X1    g338(.A(new_n382), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G8gat), .B(G36gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(G64gat), .B(G92gat), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n542), .B(new_n543), .Z(new_n544));
  NAND3_X1  g343(.A1(new_n537), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT72), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n537), .A2(KEYINPUT72), .A3(new_n541), .A4(new_n544), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n537), .A2(new_n541), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT86), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n551), .B(KEYINPUT37), .C1(KEYINPUT86), .C2(new_n537), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553));
  AOI211_X1 g352(.A(KEYINPUT38), .B(new_n544), .C1(new_n550), .C2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n549), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n544), .ZN(new_n556));
  OAI211_X1 g355(.A(KEYINPUT87), .B(new_n556), .C1(new_n550), .C2(new_n553), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT87), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n553), .B1(new_n537), .B2(new_n541), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n558), .B1(new_n559), .B2(new_n544), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n550), .A2(new_n553), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n557), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT38), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n480), .A2(new_n555), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n443), .B1(new_n463), .B2(new_n442), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT39), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n461), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT84), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n568), .B(KEYINPUT39), .C1(new_n451), .C2(new_n452), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT39), .B1(new_n451), .B2(new_n452), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT84), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n437), .A2(KEYINPUT4), .ZN(new_n572));
  INV_X1    g371(.A(new_n462), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n572), .A2(new_n573), .A3(new_n442), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n569), .B(new_n571), .C1(new_n574), .C2(new_n443), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n567), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT40), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n457), .A2(new_n468), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n461), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n567), .A2(new_n575), .A3(KEYINPUT40), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT73), .B(KEYINPUT30), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n547), .A2(new_n548), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT30), .ZN(new_n585));
  OR3_X1    g384(.A1(new_n545), .A2(KEYINPUT71), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n544), .B1(new_n537), .B2(new_n541), .ZN(new_n587));
  OAI22_X1  g386(.A1(new_n587), .A2(KEYINPUT71), .B1(new_n545), .B2(new_n585), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n584), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n582), .A2(KEYINPUT85), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT85), .B1(new_n582), .B2(new_n589), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n415), .B(new_n564), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT80), .B1(new_n480), .B2(new_n589), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n413), .A2(new_n414), .ZN(new_n594));
  INV_X1    g393(.A(new_n589), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT80), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n595), .A2(new_n596), .A3(new_n479), .A4(new_n470), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n593), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n599));
  INV_X1    g398(.A(new_n429), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(new_n502), .B2(new_n524), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n531), .A2(new_n535), .A3(new_n429), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(G227gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(new_n290), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT34), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT34), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n603), .A2(new_n609), .A3(new_n606), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT33), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G15gat), .B(G43gat), .Z(new_n614));
  XNOR2_X1  g413(.A(G71gat), .B(G99gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n608), .B(new_n610), .C1(new_n613), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n611), .A2(KEYINPUT32), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n617), .B1(new_n611), .B2(new_n612), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n609), .B1(new_n603), .B2(new_n606), .ZN(new_n622));
  AOI211_X1 g421(.A(KEYINPUT34), .B(new_n605), .C1(new_n601), .C2(new_n602), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n618), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n620), .B1(new_n618), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n599), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n624), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n619), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n618), .A2(new_n620), .A3(new_n624), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(KEYINPUT36), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n592), .A2(new_n598), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n631), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(new_n594), .ZN(new_n636));
  INV_X1    g435(.A(new_n480), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT35), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n636), .A2(new_n637), .A3(new_n638), .A4(new_n595), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n415), .A2(new_n631), .A3(new_n630), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n593), .B2(new_n597), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n639), .B1(new_n641), .B2(new_n638), .ZN(new_n642));
  AOI211_X1 g441(.A(new_n250), .B(new_n345), .C1(new_n634), .C2(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n637), .A2(KEYINPUT96), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n637), .A2(KEYINPUT96), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g447(.A(KEYINPUT16), .B(G8gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT97), .ZN(new_n650));
  NOR2_X1   g449(.A1(KEYINPUT98), .A2(KEYINPUT42), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n223), .A2(KEYINPUT42), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n643), .A2(new_n589), .ZN(new_n654));
  MUX2_X1   g453(.A(new_n652), .B(new_n653), .S(new_n654), .Z(G1325gat));
  INV_X1    g454(.A(G15gat), .ZN(new_n656));
  INV_X1    g455(.A(new_n635), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n643), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n627), .A2(new_n659), .A3(new_n632), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n627), .B2(new_n632), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n643), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n658), .B1(new_n664), .B2(new_n656), .ZN(G1326gat));
  NAND2_X1  g464(.A1(new_n643), .A2(new_n594), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT43), .B(G22gat), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n668), .B(new_n669), .Z(G1327gat));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n662), .A2(new_n592), .A3(new_n598), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n642), .A2(KEYINPUT103), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n674), .B(new_n639), .C1(new_n641), .C2(new_n638), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n672), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n671), .B1(new_n676), .B2(new_n278), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n634), .A2(new_n642), .ZN(new_n678));
  INV_X1    g477(.A(new_n278), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(KEYINPUT44), .A3(new_n679), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n320), .A2(new_n343), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n239), .A2(new_n245), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n244), .B1(new_n247), .B2(new_n235), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n246), .A2(KEYINPUT102), .A3(new_n248), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n681), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n646), .ZN(new_n692));
  OAI21_X1  g491(.A(G29gat), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n250), .B1(new_n634), .B2(new_n642), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n683), .A2(new_n278), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(new_n202), .A3(new_n646), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT45), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n693), .A2(new_n699), .ZN(G1328gat));
  OAI21_X1  g499(.A(G36gat), .B1(new_n691), .B2(new_n595), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n696), .A2(G36gat), .A3(new_n595), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT46), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(G1329gat));
  NAND3_X1  g503(.A1(new_n681), .A2(new_n663), .A3(new_n690), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G43gat), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n697), .A2(new_n206), .A3(new_n657), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n706), .A2(KEYINPUT47), .A3(new_n707), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1330gat));
  NAND2_X1  g511(.A1(new_n594), .A2(new_n208), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n696), .A2(new_n415), .ZN(new_n714));
  OAI22_X1  g513(.A1(new_n691), .A2(new_n713), .B1(new_n208), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g515(.A(new_n689), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n316), .A2(new_n322), .A3(new_n343), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n676), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n646), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n589), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n723));
  XOR2_X1   g522(.A(KEYINPUT49), .B(G64gat), .Z(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n722), .B2(new_n724), .ZN(G1333gat));
  INV_X1    g524(.A(G71gat), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n719), .A2(new_n726), .A3(new_n657), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n719), .A2(new_n663), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(new_n726), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n729), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g529(.A1(new_n719), .A2(new_n594), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G78gat), .ZN(G1335gat));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n320), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n344), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n681), .A2(new_n646), .A3(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n737), .A2(G85gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n673), .A2(new_n675), .ZN(new_n739));
  INV_X1    g538(.A(new_n672), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(new_n679), .A3(new_n734), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT51), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n676), .A2(new_n278), .A3(new_n735), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(G85gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n646), .A2(new_n748), .A3(new_n343), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n733), .B1(new_n738), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n737), .A2(G85gat), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n752), .B(KEYINPUT104), .C1(new_n747), .C2(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1336gat));
  NOR2_X1   g553(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n742), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n755), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n744), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n595), .A2(new_n344), .A3(G92gat), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n677), .A2(new_n589), .A3(new_n680), .A4(new_n736), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G92gat), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT52), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n278), .B1(new_n739), .B2(new_n740), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n745), .B1(new_n766), .B2(new_n734), .ZN(new_n767));
  NOR4_X1   g566(.A1(new_n676), .A2(KEYINPUT51), .A3(new_n278), .A4(new_n735), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT52), .B1(new_n769), .B2(new_n760), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT106), .B1(new_n770), .B2(new_n763), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n743), .A2(new_n746), .A3(new_n760), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  AND4_X1   g572(.A1(KEYINPUT106), .A2(new_n772), .A3(new_n763), .A4(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n765), .B1(new_n771), .B2(new_n774), .ZN(G1337gat));
  NAND3_X1  g574(.A1(new_n681), .A2(new_n663), .A3(new_n736), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G99gat), .ZN(new_n777));
  OR3_X1    g576(.A1(new_n635), .A2(G99gat), .A3(new_n344), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n747), .B2(new_n778), .ZN(G1338gat));
  NOR3_X1   g578(.A1(new_n415), .A2(G106gat), .A3(new_n344), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n743), .A2(new_n746), .A3(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n677), .A2(new_n594), .A3(new_n680), .A4(new_n736), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G106gat), .ZN(new_n783));
  XNOR2_X1  g582(.A(KEYINPUT107), .B(KEYINPUT53), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n757), .B1(new_n766), .B2(new_n734), .ZN(new_n787));
  NOR4_X1   g586(.A1(new_n676), .A2(new_n278), .A3(new_n735), .A4(new_n755), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n780), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n786), .B1(new_n789), .B2(new_n783), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT108), .B1(new_n785), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n759), .A2(new_n780), .B1(G106gat), .B2(new_n782), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n792), .B(new_n793), .C1(new_n794), .C2(new_n786), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n791), .A2(new_n795), .ZN(G1339gat));
  NAND2_X1  g595(.A1(new_n328), .A2(new_n329), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n334), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n328), .A2(new_n324), .A3(new_n329), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(KEYINPUT54), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n339), .ZN(new_n801));
  XOR2_X1   g600(.A(KEYINPUT109), .B(KEYINPUT54), .Z(new_n802));
  AOI21_X1  g601(.A(new_n801), .B1(new_n330), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n340), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n800), .A2(new_n803), .A3(KEYINPUT55), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n687), .A2(new_n806), .A3(new_n688), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n236), .A2(new_n237), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n228), .B1(new_n227), .B2(new_n231), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n243), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n248), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n343), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n278), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT110), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n806), .A2(new_n807), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n812), .A2(new_n679), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(new_n816), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n320), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n679), .B1(new_n808), .B2(new_n813), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT110), .B1(new_n823), .B2(new_n819), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n345), .A2(new_n717), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n692), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n636), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n829), .A2(KEYINPUT113), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(KEYINPUT113), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n595), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(new_n419), .A3(new_n717), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n594), .B1(new_n825), .B2(new_n827), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n646), .A2(new_n595), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n635), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT111), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT111), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n835), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n249), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n844), .A2(KEYINPUT112), .A3(G113gat), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT112), .B1(new_n844), .B2(G113gat), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n834), .B1(new_n845), .B2(new_n846), .ZN(G1340gat));
  NOR3_X1   g646(.A1(new_n842), .A2(new_n417), .A3(new_n344), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n343), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(new_n417), .ZN(G1341gat));
  OAI21_X1  g649(.A(G127gat), .B1(new_n842), .B2(new_n822), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n320), .A2(new_n298), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n832), .B2(new_n852), .ZN(G1342gat));
  NOR2_X1   g652(.A1(new_n278), .A2(G134gat), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  OAI22_X1  g654(.A1(new_n832), .A2(new_n855), .B1(KEYINPUT115), .B2(KEYINPUT56), .ZN(new_n856));
  NAND2_X1  g655(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT115), .B(KEYINPUT56), .C1(new_n832), .C2(new_n855), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n679), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(G134gat), .ZN(new_n862));
  AOI211_X1 g661(.A(KEYINPUT114), .B(new_n423), .C1(new_n843), .C2(new_n679), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n858), .B(new_n859), .C1(new_n862), .C2(new_n863), .ZN(G1343gat));
  NAND2_X1  g663(.A1(new_n825), .A2(new_n827), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n594), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n415), .A2(new_n868), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n806), .A2(new_n249), .A3(new_n807), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n679), .B1(new_n873), .B2(new_n813), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n822), .B1(new_n874), .B2(new_n819), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n826), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n822), .B(KEYINPUT117), .C1(new_n874), .C2(new_n819), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n870), .B(new_n872), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n876), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n827), .A3(new_n878), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT118), .B1(new_n881), .B2(new_n871), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n415), .B1(new_n825), .B2(new_n827), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT116), .B1(new_n884), .B2(KEYINPUT57), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n836), .A2(new_n663), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n359), .B1(new_n888), .B2(new_n249), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n663), .A2(new_n415), .A3(new_n589), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n828), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(G141gat), .A3(new_n250), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n892), .A2(KEYINPUT58), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n886), .A2(new_n717), .A3(new_n887), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n892), .B1(new_n894), .B2(G141gat), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n889), .A2(new_n893), .B1(new_n895), .B2(new_n896), .ZN(G1344gat));
  NAND3_X1  g696(.A1(new_n886), .A2(new_n343), .A3(new_n887), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n388), .A2(KEYINPUT59), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n345), .A2(new_n249), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT119), .B1(new_n901), .B2(new_n875), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(new_n415), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(KEYINPUT119), .A3(new_n875), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT57), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n872), .B1(new_n825), .B2(new_n827), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n343), .B(new_n887), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G148gat), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT59), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n900), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n891), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n388), .A3(new_n343), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n910), .A2(KEYINPUT120), .A3(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n898), .A2(new_n899), .B1(KEYINPUT59), .B2(new_n908), .ZN(new_n915));
  INV_X1    g714(.A(new_n912), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n913), .A2(new_n917), .ZN(G1345gat));
  AOI21_X1  g717(.A(G155gat), .B1(new_n911), .B2(new_n320), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n320), .A2(G155gat), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT121), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n919), .B1(new_n888), .B2(new_n921), .ZN(G1346gat));
  AOI21_X1  g721(.A(G162gat), .B1(new_n911), .B2(new_n679), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n278), .A2(new_n357), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n888), .B2(new_n924), .ZN(G1347gat));
  AOI21_X1  g724(.A(new_n646), .B1(new_n825), .B2(new_n827), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n640), .A2(new_n595), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT122), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n717), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n835), .A2(new_n657), .A3(new_n589), .A4(new_n692), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n932), .A2(new_n489), .A3(new_n250), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n931), .A2(new_n933), .ZN(G1348gat));
  NAND3_X1  g733(.A1(new_n930), .A2(new_n490), .A3(new_n343), .ZN(new_n935));
  OAI21_X1  g734(.A(G176gat), .B1(new_n932), .B2(new_n344), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1349gat));
  OAI21_X1  g736(.A(G183gat), .B1(new_n932), .B2(new_n822), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n320), .A2(new_n504), .A3(new_n506), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n930), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT124), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n938), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g744(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n945), .B(new_n946), .ZN(G1350gat));
  OAI21_X1  g746(.A(G190gat), .B1(new_n932), .B2(new_n278), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT61), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n930), .A2(new_n507), .A3(new_n679), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1351gat));
  OR2_X1    g750(.A1(new_n905), .A2(new_n906), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n663), .A2(new_n595), .A3(new_n646), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT126), .B1(new_n954), .B2(new_n250), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G197gat), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n954), .A2(KEYINPUT126), .A3(new_n250), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n663), .A2(new_n415), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(new_n589), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n926), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n717), .A2(new_n372), .ZN(new_n963));
  OAI22_X1  g762(.A1(new_n956), .A2(new_n957), .B1(new_n962), .B2(new_n963), .ZN(G1352gat));
  NOR3_X1   g763(.A1(new_n962), .A2(G204gat), .A3(new_n344), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT62), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n952), .A2(new_n953), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n967), .A2(KEYINPUT127), .A3(new_n343), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n969), .B1(new_n954), .B2(new_n344), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n968), .A2(G204gat), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n966), .A2(new_n971), .ZN(G1353gat));
  OR3_X1    g771(.A1(new_n962), .A2(G211gat), .A3(new_n822), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n967), .A2(new_n320), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n974), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G1354gat));
  OAI21_X1  g776(.A(G218gat), .B1(new_n954), .B2(new_n278), .ZN(new_n978));
  OR2_X1    g777(.A1(new_n278), .A2(G218gat), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n978), .B1(new_n962), .B2(new_n979), .ZN(G1355gat));
endmodule


