//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n582, new_n583, new_n584, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XOR2_X1   g032(.A(KEYINPUT66), .B(G2105), .Z(new_n458));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(KEYINPUT67), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(G125), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n458), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n458), .A2(G137), .A3(new_n459), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  XNOR2_X1  g048(.A(KEYINPUT66), .B(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n459), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n459), .A2(new_n474), .A3(KEYINPUT69), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n459), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT68), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n459), .A2(new_n484), .A3(new_n481), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n469), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI221_X1 g065(.A(new_n490), .B1(new_n489), .B2(new_n488), .C1(new_n458), .C2(G112), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n480), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT71), .ZN(G162));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT72), .B(G114), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n461), .A2(G138), .A3(new_n464), .A4(new_n458), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n474), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n459), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n499), .A2(KEYINPUT73), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(KEYINPUT73), .B1(new_n499), .B2(new_n503), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT74), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT74), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT75), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT6), .B1(new_n513), .B2(new_n514), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n508), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n517), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n527), .B1(new_n519), .B2(new_n521), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G88), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n529), .B1(new_n516), .B2(KEYINPUT75), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n524), .A2(new_n530), .ZN(G166));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT76), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n522), .A2(G51), .ZN(new_n537));
  INV_X1    g112(.A(G89), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT6), .ZN(new_n539));
  OR2_X1    g114(.A1(KEYINPUT74), .A2(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(KEYINPUT74), .A2(G651), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n511), .B1(new_n542), .B2(new_n520), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n537), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n536), .A2(new_n544), .ZN(G168));
  OAI211_X1 g120(.A(G90), .B(new_n511), .C1(new_n542), .C2(new_n520), .ZN(new_n546));
  XOR2_X1   g121(.A(KEYINPUT77), .B(G52), .Z(new_n547));
  OAI211_X1 g122(.A(G543), .B(new_n547), .C1(new_n542), .C2(new_n520), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT78), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n546), .A2(new_n548), .A3(KEYINPUT78), .ZN(new_n552));
  XNOR2_X1  g127(.A(KEYINPUT74), .B(G651), .ZN(new_n553));
  NAND2_X1  g128(.A1(G77), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G64), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n527), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n551), .A2(new_n552), .B1(new_n553), .B2(new_n556), .ZN(G171));
  NAND2_X1  g132(.A1(G68), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(new_n511), .B2(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT79), .B1(new_n560), .B2(new_n515), .ZN(new_n561));
  OAI21_X1  g136(.A(G56), .B1(new_n525), .B2(new_n526), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(new_n558), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(new_n564), .A3(new_n553), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(G43), .A2(new_n522), .B1(new_n528), .B2(G81), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n566), .A2(new_n567), .A3(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(new_n522), .A2(G53), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  XOR2_X1   g152(.A(KEYINPUT80), .B(G65), .Z(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n527), .ZN(new_n579));
  AOI22_X1  g154(.A1(G651), .A2(new_n579), .B1(new_n528), .B2(G91), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G299));
  NAND2_X1  g156(.A1(new_n556), .A2(new_n553), .ZN(new_n582));
  INV_X1    g157(.A(new_n552), .ZN(new_n583));
  AOI21_X1  g158(.A(KEYINPUT78), .B1(new_n546), .B2(new_n548), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(G301));
  INV_X1    g160(.A(G168), .ZN(G286));
  XNOR2_X1  g161(.A(G166), .B(KEYINPUT81), .ZN(G303));
  NAND2_X1  g162(.A1(new_n522), .A2(G49), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n528), .A2(G87), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n527), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(new_n553), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT83), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(G48), .A2(new_n522), .B1(new_n528), .B2(G86), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(new_n528), .A2(G85), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n522), .A2(G47), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n602), .B(new_n603), .C1(new_n515), .C2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(new_n528), .A2(G92), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT10), .Z(new_n607));
  AOI22_X1  g182(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G651), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n611));
  OAI21_X1  g186(.A(G54), .B1(new_n522), .B2(KEYINPUT84), .ZN(new_n612));
  OAI211_X1 g187(.A(KEYINPUT84), .B(G543), .C1(new_n542), .C2(new_n520), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n610), .B(new_n611), .C1(new_n612), .C2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n520), .B1(new_n553), .B2(KEYINPUT6), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n508), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n619), .A2(G54), .A3(new_n613), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n611), .B1(new_n620), .B2(new_n610), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n607), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n622), .A2(KEYINPUT86), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n622), .A2(KEYINPUT86), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  MUX2_X1   g201(.A(G301), .B(new_n625), .S(new_n626), .Z(G321));
  XNOR2_X1  g202(.A(G321), .B(KEYINPUT87), .ZN(G284));
  NAND2_X1  g203(.A1(G286), .A2(G868), .ZN(new_n629));
  AOI22_X1  g204(.A1(new_n629), .A2(KEYINPUT88), .B1(new_n626), .B2(G299), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(KEYINPUT88), .B2(new_n629), .ZN(G297));
  OAI21_X1  g206(.A(new_n630), .B1(KEYINPUT88), .B2(new_n629), .ZN(G280));
  INV_X1    g207(.A(new_n625), .ZN(new_n633));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND2_X1  g210(.A1(new_n566), .A2(new_n567), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(new_n626), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n625), .A2(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(new_n626), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n461), .A2(new_n464), .ZN(new_n641));
  INV_X1    g216(.A(new_n470), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT12), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  INV_X1    g220(.A(G2100), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n479), .A2(G123), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n486), .A2(G135), .ZN(new_n650));
  OAI221_X1 g225(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n458), .C2(G111), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n647), .A2(new_n648), .A3(new_n654), .ZN(G156));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2443), .B(G2446), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT89), .B(KEYINPUT14), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT15), .B(G2435), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2438), .ZN(new_n664));
  XOR2_X1   g239(.A(G2427), .B(G2430), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT90), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n662), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n664), .B2(new_n666), .ZN(new_n668));
  OAI21_X1  g243(.A(G14), .B1(new_n661), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n668), .B2(new_n661), .ZN(G401));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT17), .Z(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  INV_X1    g251(.A(new_n673), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(new_n671), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n675), .B(new_n676), .C1(new_n674), .C2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n676), .A2(new_n671), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT18), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(new_n653), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G2100), .ZN(G227));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT19), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n688), .A2(new_n689), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n687), .A2(new_n692), .A3(new_n690), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n687), .A2(new_n692), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT91), .B(KEYINPUT20), .ZN(new_n695));
  AOI211_X1 g270(.A(new_n691), .B(new_n693), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n694), .B2(new_n695), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT92), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n697), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OR3_X1    g280(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n702), .B2(new_n703), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(G229));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n709), .A2(G33), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n486), .A2(G139), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT95), .Z(new_n712));
  NAND3_X1  g287(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT25), .Z(new_n714));
  AND2_X1   g289(.A1(new_n461), .A2(new_n464), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n715), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n712), .B(new_n714), .C1(new_n458), .C2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n710), .B1(new_n717), .B2(G29), .ZN(new_n718));
  INV_X1    g293(.A(G2072), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT98), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n479), .A2(G129), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n486), .A2(G141), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT26), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n470), .A2(G105), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n722), .A2(new_n723), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  MUX2_X1   g302(.A(G32), .B(new_n727), .S(G29), .Z(new_n728));
  XOR2_X1   g303(.A(KEYINPUT27), .B(G1996), .Z(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n718), .B2(new_n719), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  AND2_X1   g307(.A1(KEYINPUT24), .A2(G34), .ZN(new_n733));
  NOR2_X1   g308(.A1(KEYINPUT24), .A2(G34), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n709), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT96), .Z(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G160), .B2(G29), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT97), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n721), .B(new_n731), .C1(new_n732), .C2(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT99), .ZN(new_n740));
  INV_X1    g315(.A(G16), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G6), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n599), .A2(new_n600), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(new_n741), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT32), .B(G1981), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n741), .A2(G22), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G166), .B2(new_n741), .ZN(new_n748));
  INV_X1    g323(.A(G1971), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n741), .A2(G23), .ZN(new_n751));
  INV_X1    g326(.A(new_n591), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(new_n741), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT33), .B(G1976), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n746), .A2(new_n750), .A3(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(KEYINPUT34), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(KEYINPUT34), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n479), .A2(G119), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n486), .A2(G131), .ZN(new_n760));
  OAI221_X1 g335(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n458), .C2(G107), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT93), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G29), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G25), .B2(G29), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT35), .B(G1991), .Z(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  MUX2_X1   g343(.A(G24), .B(G290), .S(G16), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1986), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n766), .B2(new_n767), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n757), .A2(new_n758), .A3(new_n768), .A4(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT36), .ZN(new_n773));
  OR3_X1    g348(.A1(new_n772), .A2(KEYINPUT94), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G29), .A2(G35), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G162), .B2(G29), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT29), .B(G2090), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT31), .B(G11), .ZN(new_n779));
  INV_X1    g354(.A(G28), .ZN(new_n780));
  AOI21_X1  g355(.A(G29), .B1(new_n780), .B2(KEYINPUT30), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(KEYINPUT101), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  OAI22_X1  g358(.A1(new_n781), .A2(KEYINPUT101), .B1(KEYINPUT30), .B2(new_n780), .ZN(new_n784));
  OAI221_X1 g359(.A(new_n779), .B1(new_n783), .B2(new_n784), .C1(new_n652), .C2(new_n709), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n741), .A2(G21), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G168), .B2(new_n741), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(G1966), .ZN(new_n788));
  AOI211_X1 g363(.A(new_n785), .B(new_n788), .C1(new_n728), .C2(new_n729), .ZN(new_n789));
  MUX2_X1   g364(.A(G19), .B(new_n636), .S(G16), .Z(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G1341), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n709), .A2(G26), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT28), .Z(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n794));
  INV_X1    g369(.A(G116), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n794), .B1(new_n474), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n479), .B2(G128), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n486), .A2(G140), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n793), .B1(new_n799), .B2(G29), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2067), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n778), .A2(new_n789), .A3(new_n791), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n787), .A2(G1966), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT100), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n741), .A2(G5), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G171), .B2(new_n741), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G1961), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n741), .A2(G20), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT23), .Z(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G299), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1956), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n738), .A2(new_n732), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n804), .A2(new_n807), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n709), .A2(G27), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G164), .B2(new_n709), .ZN(new_n815));
  INV_X1    g390(.A(G2078), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G1961), .B2(new_n806), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n802), .A2(new_n813), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n740), .A2(new_n774), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT94), .B(KEYINPUT36), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n772), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(G4), .A2(G16), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n633), .B2(G16), .ZN(new_n824));
  INV_X1    g399(.A(G1348), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n820), .A2(new_n827), .ZN(G311));
  INV_X1    g403(.A(G311), .ZN(G150));
  NAND2_X1  g404(.A1(new_n633), .A2(G559), .ZN(new_n830));
  AOI211_X1 g405(.A(KEYINPUT79), .B(new_n515), .C1(new_n562), .C2(new_n558), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n564), .B1(new_n563), .B2(new_n553), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g408(.A(G43), .B(G543), .C1(new_n542), .C2(new_n520), .ZN(new_n834));
  INV_X1    g409(.A(G81), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n543), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g411(.A(G93), .B(new_n511), .C1(new_n542), .C2(new_n520), .ZN(new_n837));
  OAI211_X1 g412(.A(G55), .B(G543), .C1(new_n542), .C2(new_n520), .ZN(new_n838));
  INV_X1    g413(.A(G67), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n509), .B2(new_n510), .ZN(new_n840));
  NAND2_X1  g415(.A1(G80), .A2(G543), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n553), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n837), .A2(new_n838), .A3(new_n843), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n833), .A2(new_n836), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n841), .B1(new_n527), .B2(new_n839), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n522), .A2(G55), .B1(new_n846), .B2(new_n553), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n566), .A2(new_n567), .B1(new_n847), .B2(new_n837), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT38), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n830), .B(new_n850), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n852), .A2(new_n853), .A3(G860), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n844), .A2(G860), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT37), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  INV_X1    g432(.A(G37), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n497), .A2(new_n498), .ZN(new_n859));
  INV_X1    g434(.A(new_n496), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n860), .A3(new_n503), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n799), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n727), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n717), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n865));
  INV_X1    g440(.A(G118), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n865), .B1(new_n474), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n479), .B2(G130), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n486), .A2(KEYINPUT102), .A3(G142), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT102), .B1(new_n486), .B2(G142), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n644), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n763), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n864), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n652), .B(G160), .ZN(new_n876));
  XNOR2_X1  g451(.A(G162), .B(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n864), .B2(new_n874), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n858), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n864), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n864), .A2(new_n882), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n877), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g463(.A1(new_n743), .A2(KEYINPUT104), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n890));
  NAND2_X1  g465(.A1(G305), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(G166), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n894));
  XNOR2_X1  g469(.A(G290), .B(new_n591), .ZN(new_n895));
  INV_X1    g470(.A(G166), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n889), .A2(new_n896), .A3(new_n891), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n889), .A2(new_n896), .A3(new_n891), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n896), .B1(new_n889), .B2(new_n891), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n895), .B(new_n894), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n849), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n638), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n849), .B1(new_n625), .B2(G559), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT41), .ZN(new_n908));
  INV_X1    g483(.A(new_n580), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n909), .B1(new_n574), .B2(new_n575), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n622), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n610), .B1(new_n612), .B2(new_n614), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT85), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n615), .ZN(new_n914));
  AOI21_X1  g489(.A(G299), .B1(new_n914), .B2(new_n607), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n908), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n622), .A2(new_n910), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(G299), .A3(new_n607), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(KEYINPUT41), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n907), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n911), .A2(new_n915), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n905), .A2(new_n924), .A3(new_n906), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n922), .B1(new_n921), .B2(new_n925), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n903), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n928), .ZN(new_n930));
  INV_X1    g505(.A(new_n903), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n931), .A3(new_n926), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(G868), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n844), .A2(new_n626), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n626), .B1(new_n929), .B2(new_n932), .ZN(new_n938));
  INV_X1    g513(.A(new_n936), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT106), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(G295));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n934), .A2(new_n942), .A3(new_n936), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT107), .B1(new_n938), .B2(new_n939), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(G331));
  OAI21_X1  g520(.A(G171), .B1(new_n845), .B2(new_n848), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n844), .B1(new_n833), .B2(new_n836), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n566), .A2(new_n567), .A3(new_n837), .A4(new_n847), .ZN(new_n948));
  NAND3_X1  g523(.A1(G301), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n946), .A2(G168), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(G168), .B1(new_n946), .B2(new_n949), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n952), .A2(new_n923), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n917), .A2(KEYINPUT41), .A3(new_n918), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT41), .B1(new_n917), .B2(new_n918), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT108), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n920), .A2(new_n958), .A3(new_n952), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n953), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n858), .B1(new_n960), .B2(new_n931), .ZN(new_n961));
  AOI211_X1 g536(.A(new_n953), .B(new_n903), .C1(new_n957), .C2(new_n959), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT43), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT109), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n965), .B(KEYINPUT43), .C1(new_n961), .C2(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n931), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  INV_X1    g543(.A(new_n953), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n956), .ZN(new_n970));
  AOI21_X1  g545(.A(G37), .B1(new_n970), .B2(new_n903), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n964), .A2(new_n966), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n968), .B1(new_n967), .B2(new_n971), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n920), .A2(new_n958), .A3(new_n952), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n958), .B1(new_n920), .B2(new_n952), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n969), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(G37), .B1(new_n977), .B2(new_n903), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n974), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  MUX2_X1   g555(.A(new_n973), .B(new_n980), .S(KEYINPUT44), .Z(G397));
  INV_X1    g556(.A(G1961), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT120), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n504), .B2(new_n505), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT50), .ZN(new_n986));
  INV_X1    g561(.A(new_n472), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n465), .A2(new_n466), .ZN(new_n988));
  OAI211_X1 g563(.A(G40), .B(new_n987), .C1(new_n988), .C2(new_n458), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n990));
  AOI21_X1  g565(.A(G1384), .B1(new_n499), .B2(new_n503), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n983), .B1(new_n986), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT73), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n861), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n499), .A2(KEYINPUT73), .A3(new_n503), .ZN(new_n996));
  AOI21_X1  g571(.A(G1384), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n992), .B(new_n983), .C1(new_n997), .C2(new_n990), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n982), .B1(new_n993), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G40), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n467), .A2(new_n472), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(new_n991), .B2(KEYINPUT45), .ZN(new_n1003));
  OAI211_X1 g578(.A(KEYINPUT45), .B(new_n984), .C1(new_n504), .C2(new_n505), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n1004), .B2(KEYINPUT118), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n997), .A2(new_n1006), .A3(KEYINPUT45), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(G2078), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1005), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n989), .B1(KEYINPUT45), .B2(new_n991), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n997), .B2(KEYINPUT45), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1011), .B(KEYINPUT111), .C1(new_n997), .C2(KEYINPUT45), .ZN(new_n1015));
  AOI21_X1  g590(.A(G2078), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1000), .B(new_n1010), .C1(new_n1016), .C2(KEYINPUT53), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT54), .B1(new_n1017), .B2(G171), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n985), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT111), .B1(new_n1020), .B2(new_n1011), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1015), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n816), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n992), .B1(new_n997), .B2(new_n990), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT120), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n998), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1023), .A2(new_n1008), .B1(new_n982), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n991), .A2(KEYINPUT45), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n1009), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n1029), .A2(new_n1003), .ZN(new_n1030));
  AOI21_X1  g605(.A(G301), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1018), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT125), .B(KEYINPUT54), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1017), .A2(G171), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1023), .A2(new_n1008), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1035), .A2(G301), .A3(new_n1000), .A4(new_n1030), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1033), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1966), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n986), .A2(new_n732), .A3(new_n992), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(G8), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G8), .ZN(new_n1042));
  NOR2_X1   g617(.A1(G168), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1043), .B(KEYINPUT124), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1041), .A2(KEYINPUT51), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT51), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(new_n1044), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1032), .A2(new_n1037), .A3(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT113), .B(G1976), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n861), .A2(new_n984), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(new_n989), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(new_n1042), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n752), .A2(G1976), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1052), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1057), .B1(KEYINPUT52), .B2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT114), .B(G1981), .Z(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT115), .B1(G305), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1060), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n599), .A2(new_n1062), .A3(new_n600), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n600), .A2(new_n597), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G1981), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT49), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1065), .A2(KEYINPUT49), .A3(new_n1067), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1055), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1059), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(G303), .A2(G8), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1075));
  XOR2_X1   g650(.A(new_n1074), .B(new_n1075), .Z(new_n1076));
  NAND3_X1  g651(.A1(new_n1014), .A2(new_n749), .A3(new_n1015), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1024), .A2(G2090), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1042), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1073), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1002), .B(KEYINPUT116), .C1(new_n991), .C2(new_n990), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1053), .A2(KEYINPUT50), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT116), .B1(new_n1083), .B2(new_n1002), .ZN(new_n1084));
  OR3_X1    g659(.A1(new_n1082), .A2(new_n1084), .A3(G2090), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1085), .A2(new_n1077), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1085), .B2(new_n1077), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1087), .A2(new_n1088), .A3(new_n1042), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1080), .B1(new_n1089), .B2(new_n1076), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT126), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT126), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1080), .B(new_n1092), .C1(new_n1089), .C2(new_n1076), .ZN(new_n1093));
  NAND2_X1  g668(.A1(G299), .A2(KEYINPUT119), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n910), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1094), .A2(new_n1096), .A3(KEYINPUT57), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G1956), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1028), .A2(new_n1002), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n985), .B2(new_n1019), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT56), .B(G2072), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1101), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1054), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(G2067), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n1026), .B2(new_n825), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(new_n625), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1101), .A2(new_n1103), .A3(new_n1107), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1108), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1117), .B(KEYINPUT122), .Z(new_n1118));
  INV_X1    g693(.A(G1996), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT58), .B(G1341), .Z(new_n1120));
  AOI22_X1  g695(.A1(new_n1105), .A2(new_n1119), .B1(new_n1109), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1116), .B(new_n1118), .C1(new_n1121), .C2(new_n636), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1118), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1020), .A2(new_n1119), .A3(new_n1011), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1109), .A2(new_n1120), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n636), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1123), .B1(new_n1126), .B2(new_n1115), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1113), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1130), .B2(new_n1108), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1134), .A2(new_n1113), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1128), .B(new_n1131), .C1(new_n1135), .C2(new_n1129), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n633), .B1(new_n1111), .B2(KEYINPUT60), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1111), .A2(KEYINPUT60), .ZN(new_n1138));
  AOI21_X1  g713(.A(G1348), .B1(new_n1025), .B2(new_n998), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n1140));
  NOR4_X1   g715(.A1(new_n1139), .A2(new_n1140), .A3(new_n625), .A4(new_n1110), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1137), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1114), .B1(new_n1136), .B2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1050), .A2(new_n1091), .A3(new_n1093), .A4(new_n1143), .ZN(new_n1144));
  AOI211_X1 g719(.A(G1976), .B(G288), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1065), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1055), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1147), .B1(new_n1148), .B2(new_n1073), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1041), .A2(G286), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1080), .B(new_n1151), .C1(new_n1089), .C2(new_n1076), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT63), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1155), .B(new_n1080), .C1(new_n1079), .C2(new_n1076), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1149), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1045), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n1160), .A2(KEYINPUT62), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1034), .B1(new_n1160), .B2(KEYINPUT62), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1161), .A2(new_n1162), .A3(new_n1091), .A4(new_n1093), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1144), .A2(new_n1157), .A3(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n989), .A2(new_n991), .A3(KEYINPUT45), .ZN(new_n1165));
  NAND2_X1  g740(.A1(G290), .A2(G1986), .ZN(new_n1166));
  NOR2_X1   g741(.A1(G290), .A2(G1986), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1167), .A2(KEYINPUT110), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1165), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1169), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n764), .A2(new_n767), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n799), .A2(G2067), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n799), .A2(G2067), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n727), .B(new_n1119), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n764), .A2(new_n767), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1171), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1170), .B1(new_n1177), .B2(new_n1165), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1164), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1174), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1165), .B1(new_n1180), .B2(new_n727), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1165), .A2(new_n1119), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(KEYINPUT46), .ZN(new_n1183));
  OR2_X1    g758(.A1(new_n1182), .A2(KEYINPUT46), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1181), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT47), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1177), .A2(new_n1165), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT48), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1172), .B1(new_n1193), .B2(new_n1176), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1165), .ZN(new_n1195));
  AND4_X1   g770(.A1(new_n1187), .A2(new_n1191), .A3(new_n1192), .A4(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1179), .A2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g772(.A(G319), .ZN(new_n1199));
  NOR3_X1   g773(.A1(G227), .A2(new_n1199), .A3(G401), .ZN(new_n1200));
  NAND3_X1  g774(.A1(new_n706), .A2(new_n707), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g775(.A(new_n1201), .ZN(new_n1202));
  OAI21_X1  g776(.A(new_n1202), .B1(new_n879), .B2(new_n885), .ZN(new_n1203));
  AND3_X1   g777(.A1(new_n967), .A2(new_n968), .A3(new_n971), .ZN(new_n1204));
  AOI21_X1  g778(.A(new_n1204), .B1(new_n963), .B2(KEYINPUT109), .ZN(new_n1205));
  AOI211_X1 g779(.A(KEYINPUT127), .B(new_n1203), .C1(new_n1205), .C2(new_n966), .ZN(new_n1206));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n1207));
  INV_X1    g781(.A(new_n1203), .ZN(new_n1208));
  AOI21_X1  g782(.A(new_n1207), .B1(new_n973), .B2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g783(.A1(new_n1206), .A2(new_n1209), .ZN(G308));
  AOI21_X1  g784(.A(new_n968), .B1(new_n978), .B2(new_n967), .ZN(new_n1211));
  OAI21_X1  g785(.A(new_n972), .B1(new_n1211), .B2(new_n965), .ZN(new_n1212));
  INV_X1    g786(.A(new_n966), .ZN(new_n1213));
  OAI21_X1  g787(.A(new_n1208), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n1214), .A2(KEYINPUT127), .ZN(new_n1215));
  NAND3_X1  g789(.A1(new_n973), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n1215), .A2(new_n1216), .ZN(G225));
endmodule


