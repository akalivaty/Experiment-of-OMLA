

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790;

  INV_X1 U375 ( .A(n696), .ZN(n358) );
  INV_X1 U376 ( .A(n696), .ZN(n362) );
  INV_X1 U377 ( .A(n681), .ZN(n360) );
  INV_X1 U378 ( .A(n694), .ZN(n364) );
  AND2_X1 U379 ( .A1(n377), .A2(n376), .ZN(n381) );
  INV_X1 U380 ( .A(n618), .ZN(n355) );
  XNOR2_X1 U381 ( .A(n423), .B(KEYINPUT32), .ZN(n409) );
  XNOR2_X1 U382 ( .A(n582), .B(KEYINPUT6), .ZN(n609) );
  XNOR2_X1 U383 ( .A(KEYINPUT90), .B(G113), .ZN(n531) );
  INV_X2 U384 ( .A(G953), .ZN(n771) );
  XNOR2_X1 U385 ( .A(n354), .B(n533), .ZN(n538) );
  XNOR2_X1 U386 ( .A(n535), .B(n532), .ZN(n354) );
  XNOR2_X2 U387 ( .A(n356), .B(n355), .ZN(n787) );
  NAND2_X1 U388 ( .A1(n617), .A2(n717), .ZN(n356) );
  INV_X1 U389 ( .A(n357), .ZN(n684) );
  NAND2_X1 U390 ( .A1(n359), .A2(n358), .ZN(n357) );
  XNOR2_X1 U391 ( .A(n682), .B(n360), .ZN(n359) );
  NAND2_X1 U392 ( .A1(n394), .A2(n540), .ZN(n542) );
  XNOR2_X2 U393 ( .A(n539), .B(n370), .ZN(n394) );
  INV_X1 U394 ( .A(n361), .ZN(n698) );
  NAND2_X1 U395 ( .A1(n363), .A2(n362), .ZN(n361) );
  XNOR2_X1 U396 ( .A(n695), .B(n364), .ZN(n363) );
  NOR2_X1 U397 ( .A1(G237), .A2(KEYINPUT75), .ZN(n396) );
  BUF_X1 U398 ( .A(G107), .Z(n373) );
  XNOR2_X2 U399 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n422) );
  INV_X2 U400 ( .A(G107), .ZN(n393) );
  NOR2_X2 U401 ( .A1(n372), .A2(n496), .ZN(n498) );
  AND2_X1 U402 ( .A1(n662), .A2(n661), .ZN(n664) );
  AND2_X1 U403 ( .A1(n689), .A2(n661), .ZN(n690) );
  XNOR2_X1 U404 ( .A(n385), .B(n384), .ZN(n416) );
  NAND2_X1 U405 ( .A1(n543), .A2(n424), .ZN(n423) );
  NOR2_X1 U406 ( .A1(n564), .A2(n573), .ZN(n417) );
  XNOR2_X1 U407 ( .A(n648), .B(n585), .ZN(n595) );
  XNOR2_X1 U408 ( .A(n680), .B(KEYINPUT59), .ZN(n681) );
  XNOR2_X1 U409 ( .A(n512), .B(n418), .ZN(n599) );
  NAND2_X1 U410 ( .A1(n436), .A2(n433), .ZN(n432) );
  NOR2_X2 U411 ( .A1(n787), .A2(n641), .ZN(n445) );
  XNOR2_X1 U412 ( .A(n550), .B(KEYINPUT33), .ZN(n702) );
  XNOR2_X1 U413 ( .A(n417), .B(n565), .ZN(n724) );
  INV_X1 U414 ( .A(KEYINPUT66), .ZN(n457) );
  XNOR2_X1 U415 ( .A(G902), .B(KEYINPUT15), .ZN(n656) );
  XNOR2_X1 U416 ( .A(n410), .B(G125), .ZN(n499) );
  XNOR2_X1 U417 ( .A(KEYINPUT10), .B(G146), .ZN(n410) );
  OR2_X2 U418 ( .A1(n388), .A2(n386), .ZN(n558) );
  NAND2_X1 U419 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U420 ( .A1(n420), .A2(G902), .ZN(n389) );
  XNOR2_X1 U421 ( .A(n487), .B(n486), .ZN(n569) );
  XNOR2_X1 U422 ( .A(n403), .B(n463), .ZN(n537) );
  XOR2_X1 U423 ( .A(KEYINPUT72), .B(KEYINPUT3), .Z(n463) );
  XNOR2_X1 U424 ( .A(n462), .B(KEYINPUT81), .ZN(n403) );
  XNOR2_X1 U425 ( .A(G119), .B(G101), .ZN(n462) );
  XNOR2_X1 U426 ( .A(n426), .B(G122), .ZN(n478) );
  XNOR2_X1 U427 ( .A(G113), .B(G104), .ZN(n426) );
  INV_X1 U428 ( .A(G110), .ZN(n392) );
  XNOR2_X1 U429 ( .A(n448), .B(n447), .ZN(n506) );
  INV_X1 U430 ( .A(KEYINPUT8), .ZN(n447) );
  NAND2_X1 U431 ( .A1(n771), .A2(G234), .ZN(n448) );
  XNOR2_X1 U432 ( .A(G143), .B(G140), .ZN(n479) );
  XNOR2_X1 U433 ( .A(n478), .B(KEYINPUT11), .ZN(n411) );
  NAND2_X1 U434 ( .A1(n653), .A2(n652), .ZN(n439) );
  XNOR2_X1 U435 ( .A(n429), .B(n593), .ZN(n642) );
  NAND2_X1 U436 ( .A1(n431), .A2(n430), .ZN(n429) );
  XNOR2_X1 U437 ( .A(n511), .B(n515), .ZN(n418) );
  XNOR2_X1 U438 ( .A(n492), .B(G478), .ZN(n567) );
  INV_X1 U439 ( .A(n717), .ZN(n573) );
  NAND2_X1 U440 ( .A1(n457), .A2(KEYINPUT44), .ZN(n456) );
  INV_X1 U441 ( .A(G237), .ZN(n399) );
  INV_X1 U442 ( .A(G953), .ZN(n400) );
  NAND2_X1 U443 ( .A1(n528), .A2(n540), .ZN(n387) );
  XNOR2_X1 U444 ( .A(G137), .B(G116), .ZN(n534) );
  NAND2_X1 U445 ( .A1(n382), .A2(KEYINPUT66), .ZN(n380) );
  NAND2_X1 U446 ( .A1(n397), .A2(n395), .ZN(n530) );
  NAND2_X1 U447 ( .A1(n398), .A2(KEYINPUT75), .ZN(n397) );
  NAND2_X1 U448 ( .A1(n771), .A2(n396), .ZN(n395) );
  NAND2_X1 U449 ( .A1(n400), .A2(n399), .ZN(n398) );
  XNOR2_X1 U450 ( .A(n518), .B(n517), .ZN(n421) );
  INV_X1 U451 ( .A(G134), .ZN(n517) );
  INV_X1 U452 ( .A(n656), .ZN(n438) );
  NAND2_X1 U453 ( .A1(n435), .A2(n434), .ZN(n433) );
  NAND2_X1 U454 ( .A1(G234), .A2(G237), .ZN(n467) );
  NOR2_X2 U455 ( .A1(n611), .A2(n612), .ZN(n643) );
  XNOR2_X1 U456 ( .A(G128), .B(KEYINPUT86), .ZN(n500) );
  INV_X1 U457 ( .A(KEYINPUT23), .ZN(n502) );
  XNOR2_X1 U458 ( .A(G119), .B(G110), .ZN(n503) );
  XNOR2_X1 U459 ( .A(G137), .B(G140), .ZN(n521) );
  XNOR2_X1 U460 ( .A(G110), .B(n373), .ZN(n523) );
  XNOR2_X1 U461 ( .A(n459), .B(KEYINPUT17), .ZN(n407) );
  XNOR2_X1 U462 ( .A(G146), .B(G125), .ZN(n459) );
  XNOR2_X1 U463 ( .A(KEYINPUT18), .B(KEYINPUT82), .ZN(n406) );
  NOR2_X1 U464 ( .A1(n706), .A2(n705), .ZN(n598) );
  INV_X1 U465 ( .A(KEYINPUT34), .ZN(n415) );
  INV_X1 U466 ( .A(KEYINPUT98), .ZN(n412) );
  INV_X1 U467 ( .A(KEYINPUT31), .ZN(n384) );
  BUF_X1 U468 ( .A(n584), .Z(n648) );
  INV_X1 U469 ( .A(KEYINPUT91), .ZN(n453) );
  XNOR2_X1 U470 ( .A(n401), .B(n478), .ZN(n404) );
  XNOR2_X1 U471 ( .A(n488), .B(n391), .ZN(n401) );
  XNOR2_X1 U472 ( .A(n392), .B(KEYINPUT16), .ZN(n391) );
  XNOR2_X1 U473 ( .A(n451), .B(n449), .ZN(n678) );
  XNOR2_X1 U474 ( .A(n490), .B(n450), .ZN(n449) );
  XNOR2_X1 U475 ( .A(n491), .B(n489), .ZN(n451) );
  XNOR2_X1 U476 ( .A(n477), .B(n411), .ZN(n485) );
  XNOR2_X1 U477 ( .A(n770), .B(n402), .ZN(n693) );
  XNOR2_X1 U478 ( .A(n461), .B(n371), .ZN(n402) );
  XNOR2_X1 U479 ( .A(n407), .B(n406), .ZN(n461) );
  XNOR2_X1 U480 ( .A(n519), .B(n460), .ZN(n371) );
  XNOR2_X1 U481 ( .A(n594), .B(KEYINPUT40), .ZN(n670) );
  NOR2_X1 U482 ( .A1(n620), .A2(n419), .ZN(n622) );
  NAND2_X1 U483 ( .A1(n452), .A2(n759), .ZN(n743) );
  NOR2_X2 U484 ( .A1(n567), .A2(n446), .ZN(n755) );
  INV_X1 U485 ( .A(n566), .ZN(n452) );
  XNOR2_X1 U486 ( .A(n577), .B(KEYINPUT97), .ZN(n789) );
  INV_X1 U487 ( .A(n439), .ZN(n699) );
  NOR2_X1 U488 ( .A1(n732), .A2(n419), .ZN(n365) );
  AND2_X1 U489 ( .A1(n409), .A2(n428), .ZN(n366) );
  XOR2_X1 U490 ( .A(n687), .B(n686), .Z(n367) );
  XOR2_X1 U491 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n368) );
  XOR2_X1 U492 ( .A(KEYINPUT70), .B(KEYINPUT48), .Z(n369) );
  XNOR2_X1 U493 ( .A(n404), .B(n537), .ZN(n770) );
  INV_X1 U494 ( .A(n529), .ZN(n370) );
  XNOR2_X2 U495 ( .A(n777), .B(G146), .ZN(n529) );
  OR2_X1 U496 ( .A1(n724), .A2(n372), .ZN(n385) );
  XNOR2_X1 U497 ( .A(n372), .B(KEYINPUT85), .ZN(n405) );
  XNOR2_X2 U498 ( .A(n476), .B(n475), .ZN(n372) );
  XNOR2_X1 U499 ( .A(n606), .B(n466), .ZN(n620) );
  NAND2_X1 U500 ( .A1(n374), .A2(n570), .ZN(n572) );
  NAND2_X1 U501 ( .A1(n566), .A2(n416), .ZN(n374) );
  AND2_X1 U502 ( .A1(n375), .A2(n789), .ZN(n376) );
  XNOR2_X1 U503 ( .A(n572), .B(n571), .ZN(n375) );
  NAND2_X1 U504 ( .A1(n378), .A2(n557), .ZN(n377) );
  NAND2_X1 U505 ( .A1(n556), .A2(n672), .ZN(n378) );
  NAND2_X1 U506 ( .A1(n381), .A2(n379), .ZN(n580) );
  NAND2_X1 U507 ( .A1(n366), .A2(n380), .ZN(n379) );
  NAND2_X1 U508 ( .A1(n672), .A2(n578), .ZN(n382) );
  NAND2_X1 U509 ( .A1(n383), .A2(KEYINPUT2), .ZN(n441) );
  OR2_X2 U510 ( .A1(n653), .A2(n654), .ZN(n383) );
  XNOR2_X2 U511 ( .A(n580), .B(n579), .ZN(n653) );
  INV_X1 U512 ( .A(n416), .ZN(n760) );
  XNOR2_X2 U513 ( .A(n558), .B(KEYINPUT1), .ZN(n717) );
  NOR2_X1 U514 ( .A1(n687), .A2(n387), .ZN(n386) );
  NAND2_X1 U515 ( .A1(n687), .A2(n420), .ZN(n390) );
  XNOR2_X2 U516 ( .A(n529), .B(n527), .ZN(n687) );
  XNOR2_X2 U517 ( .A(n393), .B(G116), .ZN(n488) );
  XNOR2_X1 U518 ( .A(n394), .B(KEYINPUT62), .ZN(n458) );
  XNOR2_X2 U519 ( .A(n408), .B(n422), .ZN(n519) );
  NAND2_X1 U520 ( .A1(n405), .A2(n561), .ZN(n562) );
  NAND2_X1 U521 ( .A1(n702), .A2(n405), .ZN(n551) );
  XNOR2_X1 U522 ( .A(n408), .B(G134), .ZN(n450) );
  XNOR2_X2 U523 ( .A(G143), .B(G128), .ZN(n408) );
  NAND2_X1 U524 ( .A1(n454), .A2(n409), .ZN(n455) );
  XNOR2_X1 U525 ( .A(n409), .B(G119), .ZN(G21) );
  NOR2_X1 U526 ( .A1(n425), .A2(n609), .ZN(n424) );
  XNOR2_X1 U527 ( .A(n616), .B(KEYINPUT36), .ZN(n617) );
  NOR2_X2 U528 ( .A1(n576), .A2(n546), .ZN(n666) );
  XNOR2_X1 U529 ( .A(n413), .B(n412), .ZN(n425) );
  NOR2_X1 U530 ( .A1(n573), .A2(n713), .ZN(n413) );
  NAND2_X1 U531 ( .A1(n717), .A2(n718), .ZN(n548) );
  NAND2_X2 U532 ( .A1(n414), .A2(n553), .ZN(n555) );
  XNOR2_X2 U533 ( .A(n551), .B(n415), .ZN(n414) );
  NAND2_X1 U534 ( .A1(n693), .A2(n656), .ZN(n427) );
  AND2_X2 U535 ( .A1(n441), .A2(n440), .ZN(n700) );
  NAND2_X1 U536 ( .A1(n655), .A2(n652), .ZN(n440) );
  NAND2_X1 U537 ( .A1(n670), .A2(n790), .ZN(n444) );
  XNOR2_X1 U538 ( .A(n444), .B(n368), .ZN(n443) );
  NOR2_X2 U539 ( .A1(n700), .A2(n432), .ZN(n659) );
  XNOR2_X1 U540 ( .A(n505), .B(n504), .ZN(n508) );
  INV_X1 U541 ( .A(n558), .ZN(n419) );
  INV_X1 U542 ( .A(n528), .ZN(n420) );
  XNOR2_X2 U543 ( .A(n519), .B(n421), .ZN(n777) );
  XNOR2_X2 U544 ( .A(KEYINPUT69), .B(G131), .ZN(n518) );
  XNOR2_X2 U545 ( .A(n427), .B(n464), .ZN(n584) );
  INV_X1 U546 ( .A(n666), .ZN(n428) );
  NAND2_X1 U547 ( .A1(n642), .A2(n755), .ZN(n594) );
  NOR2_X1 U548 ( .A1(n629), .A2(n591), .ZN(n430) );
  INV_X1 U549 ( .A(n630), .ZN(n431) );
  NAND2_X1 U550 ( .A1(n439), .A2(n438), .ZN(n437) );
  INV_X1 U551 ( .A(n653), .ZN(n765) );
  INV_X1 U552 ( .A(n657), .ZN(n434) );
  NOR2_X1 U553 ( .A1(n653), .A2(n656), .ZN(n435) );
  NAND2_X1 U554 ( .A1(n437), .A2(n657), .ZN(n436) );
  BUF_X2 U555 ( .A(n691), .Z(n673) );
  XNOR2_X1 U556 ( .A(n442), .B(n369), .ZN(n651) );
  NAND2_X1 U557 ( .A1(n445), .A2(n443), .ZN(n442) );
  NAND2_X1 U558 ( .A1(n567), .A2(n446), .ZN(n568) );
  INV_X1 U559 ( .A(n569), .ZN(n446) );
  NAND2_X1 U560 ( .A1(n452), .A2(n755), .ZN(n742) );
  XNOR2_X2 U561 ( .A(n562), .B(n453), .ZN(n566) );
  NOR2_X1 U562 ( .A1(n666), .A2(n578), .ZN(n454) );
  NAND2_X1 U563 ( .A1(n455), .A2(n456), .ZN(n556) );
  NOR2_X1 U564 ( .A1(n771), .A2(G952), .ZN(n696) );
  INV_X1 U565 ( .A(n582), .ZN(n563) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(n504) );
  INV_X1 U567 ( .A(KEYINPUT92), .ZN(n565) );
  XNOR2_X1 U568 ( .A(n514), .B(n513), .ZN(n515) );
  BUF_X1 U569 ( .A(n654), .Z(n779) );
  INV_X1 U570 ( .A(n696), .ZN(n661) );
  INV_X1 U571 ( .A(KEYINPUT63), .ZN(n663) );
  AND2_X1 U572 ( .A1(G224), .A2(n771), .ZN(n460) );
  INV_X1 U573 ( .A(G902), .ZN(n540) );
  NAND2_X1 U574 ( .A1(n540), .A2(n399), .ZN(n465) );
  AND2_X1 U575 ( .A1(n465), .A2(G210), .ZN(n464) );
  NAND2_X1 U576 ( .A1(n465), .A2(G214), .ZN(n703) );
  NAND2_X1 U577 ( .A1(n584), .A2(n703), .ZN(n606) );
  INV_X1 U578 ( .A(KEYINPUT19), .ZN(n466) );
  XNOR2_X1 U579 ( .A(n467), .B(KEYINPUT14), .ZN(n471) );
  AND2_X1 U580 ( .A1(n471), .A2(G952), .ZN(n730) );
  NAND2_X1 U581 ( .A1(n730), .A2(n771), .ZN(n469) );
  INV_X1 U582 ( .A(KEYINPUT83), .ZN(n468) );
  XNOR2_X1 U583 ( .A(n469), .B(n468), .ZN(n590) );
  AND2_X1 U584 ( .A1(G953), .A2(G902), .ZN(n470) );
  NAND2_X1 U585 ( .A1(n471), .A2(n470), .ZN(n586) );
  NOR2_X1 U586 ( .A1(G898), .A2(n586), .ZN(n472) );
  XOR2_X1 U587 ( .A(n472), .B(KEYINPUT84), .Z(n473) );
  AND2_X1 U588 ( .A1(n590), .A2(n473), .ZN(n474) );
  NOR2_X2 U589 ( .A1(n620), .A2(n474), .ZN(n476) );
  INV_X1 U590 ( .A(KEYINPUT0), .ZN(n475) );
  INV_X1 U591 ( .A(n499), .ZN(n477) );
  XOR2_X1 U592 ( .A(KEYINPUT93), .B(KEYINPUT12), .Z(n480) );
  XNOR2_X1 U593 ( .A(n480), .B(n479), .ZN(n483) );
  NAND2_X1 U594 ( .A1(n530), .A2(G214), .ZN(n481) );
  XNOR2_X1 U595 ( .A(n481), .B(n518), .ZN(n482) );
  XNOR2_X1 U596 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U597 ( .A(n485), .B(n484), .ZN(n680) );
  NAND2_X1 U598 ( .A1(n680), .A2(n540), .ZN(n487) );
  XOR2_X1 U599 ( .A(KEYINPUT13), .B(G475), .Z(n486) );
  XOR2_X1 U600 ( .A(KEYINPUT7), .B(n488), .Z(n491) );
  NAND2_X1 U601 ( .A1(G217), .A2(n506), .ZN(n489) );
  XOR2_X1 U602 ( .A(G122), .B(KEYINPUT9), .Z(n490) );
  NAND2_X1 U603 ( .A1(n678), .A2(n540), .ZN(n492) );
  NOR2_X1 U604 ( .A1(n569), .A2(n567), .ZN(n596) );
  NAND2_X1 U605 ( .A1(G234), .A2(n656), .ZN(n493) );
  XNOR2_X1 U606 ( .A(KEYINPUT20), .B(n493), .ZN(n510) );
  NAND2_X1 U607 ( .A1(n510), .A2(G221), .ZN(n495) );
  INV_X1 U608 ( .A(KEYINPUT21), .ZN(n494) );
  XNOR2_X1 U609 ( .A(n495), .B(n494), .ZN(n712) );
  NAND2_X1 U610 ( .A1(n596), .A2(n712), .ZN(n496) );
  XNOR2_X1 U611 ( .A(KEYINPUT67), .B(KEYINPUT22), .ZN(n497) );
  XNOR2_X1 U612 ( .A(n498), .B(n497), .ZN(n544) );
  INV_X1 U613 ( .A(n544), .ZN(n543) );
  XNOR2_X1 U614 ( .A(n499), .B(n521), .ZN(n775) );
  XOR2_X1 U615 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n501) );
  XNOR2_X1 U616 ( .A(n501), .B(n500), .ZN(n505) );
  AND2_X1 U617 ( .A1(n506), .A2(G221), .ZN(n507) );
  XNOR2_X1 U618 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U619 ( .A(n775), .B(n509), .ZN(n675) );
  NOR2_X1 U620 ( .A1(G902), .A2(n675), .ZN(n512) );
  NAND2_X1 U621 ( .A1(n510), .A2(G217), .ZN(n511) );
  XNOR2_X1 U622 ( .A(KEYINPUT76), .B(KEYINPUT88), .ZN(n514) );
  INV_X1 U623 ( .A(KEYINPUT25), .ZN(n513) );
  INV_X1 U624 ( .A(KEYINPUT96), .ZN(n516) );
  XNOR2_X1 U625 ( .A(n599), .B(n516), .ZN(n713) );
  NAND2_X1 U626 ( .A1(n771), .A2(G227), .ZN(n520) );
  XNOR2_X1 U627 ( .A(n520), .B(KEYINPUT77), .ZN(n522) );
  XNOR2_X1 U628 ( .A(n522), .B(n521), .ZN(n526) );
  XNOR2_X1 U629 ( .A(G104), .B(G101), .ZN(n524) );
  XNOR2_X1 U630 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U631 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U632 ( .A(KEYINPUT71), .B(G469), .ZN(n528) );
  NAND2_X1 U633 ( .A1(n530), .A2(G210), .ZN(n533) );
  XNOR2_X1 U634 ( .A(n531), .B(KEYINPUT74), .ZN(n532) );
  XNOR2_X1 U635 ( .A(n534), .B(KEYINPUT5), .ZN(n535) );
  XNOR2_X1 U636 ( .A(n538), .B(n537), .ZN(n539) );
  INV_X1 U637 ( .A(G472), .ZN(n541) );
  XNOR2_X2 U638 ( .A(n542), .B(n541), .ZN(n582) );
  BUF_X1 U639 ( .A(n544), .Z(n576) );
  AND2_X1 U640 ( .A1(n599), .A2(n582), .ZN(n545) );
  NAND2_X1 U641 ( .A1(n545), .A2(n573), .ZN(n546) );
  INV_X1 U642 ( .A(n712), .ZN(n547) );
  NOR2_X1 U643 ( .A1(n599), .A2(n547), .ZN(n718) );
  XNOR2_X1 U644 ( .A(n548), .B(KEYINPUT99), .ZN(n549) );
  NAND2_X1 U645 ( .A1(n549), .A2(n609), .ZN(n550) );
  NAND2_X1 U646 ( .A1(n569), .A2(n567), .ZN(n552) );
  XNOR2_X1 U647 ( .A(n552), .B(KEYINPUT100), .ZN(n633) );
  INV_X1 U648 ( .A(n633), .ZN(n553) );
  INV_X1 U649 ( .A(KEYINPUT35), .ZN(n554) );
  XNOR2_X2 U650 ( .A(n555), .B(n554), .ZN(n672) );
  INV_X1 U651 ( .A(KEYINPUT44), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n578), .A2(KEYINPUT66), .ZN(n557) );
  NAND2_X1 U653 ( .A1(n718), .A2(n558), .ZN(n560) );
  INV_X1 U654 ( .A(KEYINPUT89), .ZN(n559) );
  XNOR2_X1 U655 ( .A(n560), .B(n559), .ZN(n630) );
  NOR2_X1 U656 ( .A1(n630), .A2(n563), .ZN(n561) );
  NAND2_X1 U657 ( .A1(n718), .A2(n563), .ZN(n564) );
  XNOR2_X1 U658 ( .A(n568), .B(KEYINPUT94), .ZN(n747) );
  INV_X1 U659 ( .A(n755), .ZN(n612) );
  AND2_X1 U660 ( .A1(n747), .A2(n612), .ZN(n707) );
  INV_X1 U661 ( .A(KEYINPUT78), .ZN(n636) );
  XNOR2_X1 U662 ( .A(n707), .B(n636), .ZN(n570) );
  INV_X1 U663 ( .A(KEYINPUT95), .ZN(n571) );
  NAND2_X1 U664 ( .A1(n713), .A2(n573), .ZN(n574) );
  OR2_X1 U665 ( .A1(n574), .A2(n609), .ZN(n575) );
  NOR2_X1 U666 ( .A1(n576), .A2(n575), .ZN(n577) );
  INV_X1 U667 ( .A(KEYINPUT45), .ZN(n579) );
  INV_X1 U668 ( .A(n703), .ZN(n581) );
  OR2_X1 U669 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U670 ( .A(n583), .B(KEYINPUT30), .ZN(n629) );
  INV_X1 U671 ( .A(KEYINPUT38), .ZN(n585) );
  XNOR2_X1 U672 ( .A(n586), .B(KEYINPUT101), .ZN(n588) );
  INV_X1 U673 ( .A(G900), .ZN(n587) );
  NAND2_X1 U674 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U675 ( .A1(n590), .A2(n589), .ZN(n631) );
  NAND2_X1 U676 ( .A1(n595), .A2(n631), .ZN(n591) );
  INV_X1 U677 ( .A(KEYINPUT73), .ZN(n592) );
  XNOR2_X1 U678 ( .A(n592), .B(KEYINPUT39), .ZN(n593) );
  NAND2_X1 U679 ( .A1(n595), .A2(n703), .ZN(n706) );
  INV_X1 U680 ( .A(n596), .ZN(n705) );
  XNOR2_X1 U681 ( .A(KEYINPUT41), .B(KEYINPUT104), .ZN(n597) );
  XNOR2_X1 U682 ( .A(n598), .B(n597), .ZN(n732) );
  NAND2_X1 U683 ( .A1(n599), .A2(n712), .ZN(n607) );
  INV_X1 U684 ( .A(n631), .ZN(n608) );
  OR2_X1 U685 ( .A1(n608), .A2(n582), .ZN(n600) );
  OR2_X1 U686 ( .A1(n607), .A2(n600), .ZN(n602) );
  INV_X1 U687 ( .A(KEYINPUT28), .ZN(n601) );
  XNOR2_X1 U688 ( .A(n602), .B(n601), .ZN(n621) );
  NAND2_X1 U689 ( .A1(n365), .A2(n621), .ZN(n605) );
  INV_X1 U690 ( .A(KEYINPUT105), .ZN(n603) );
  XNOR2_X1 U691 ( .A(n603), .B(KEYINPUT42), .ZN(n604) );
  XNOR2_X1 U692 ( .A(n605), .B(n604), .ZN(n790) );
  BUF_X1 U693 ( .A(n606), .Z(n615) );
  INV_X1 U694 ( .A(KEYINPUT106), .ZN(n613) );
  NOR2_X1 U695 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U696 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U697 ( .A(n613), .B(n643), .ZN(n614) );
  NOR2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n616) );
  INV_X1 U699 ( .A(KEYINPUT107), .ZN(n618) );
  AND2_X1 U700 ( .A1(n622), .A2(n621), .ZN(n756) );
  INV_X1 U701 ( .A(n707), .ZN(n623) );
  AND2_X1 U702 ( .A1(n756), .A2(n623), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n624), .A2(KEYINPUT47), .ZN(n628) );
  INV_X1 U704 ( .A(KEYINPUT47), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n624), .A2(KEYINPUT78), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n640) );
  OR2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n648), .A2(n631), .ZN(n632) );
  OR2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n634) );
  OR2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n754) );
  AND2_X1 U712 ( .A1(n707), .A2(n636), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n756), .A2(n637), .ZN(n638) );
  AND2_X1 U714 ( .A1(n754), .A2(n638), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n641) );
  INV_X1 U716 ( .A(n747), .ZN(n759) );
  NAND2_X1 U717 ( .A1(n642), .A2(n759), .ZN(n665) );
  NAND2_X1 U718 ( .A1(n703), .A2(n643), .ZN(n644) );
  OR2_X1 U719 ( .A1(n717), .A2(n644), .ZN(n647) );
  XNOR2_X1 U720 ( .A(KEYINPUT43), .B(KEYINPUT102), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n645), .B(KEYINPUT103), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n647), .B(n646), .ZN(n649) );
  OR2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n764) );
  AND2_X1 U724 ( .A1(n665), .A2(n764), .ZN(n650) );
  NAND2_X1 U725 ( .A1(n651), .A2(n650), .ZN(n654) );
  INV_X1 U726 ( .A(KEYINPUT2), .ZN(n652) );
  INV_X1 U727 ( .A(n654), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n655), .A2(KEYINPUT79), .ZN(n657) );
  INV_X1 U729 ( .A(KEYINPUT65), .ZN(n658) );
  XNOR2_X2 U730 ( .A(n659), .B(n658), .ZN(n691) );
  NAND2_X1 U731 ( .A1(n691), .A2(G472), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n660), .B(n458), .ZN(n662) );
  XNOR2_X1 U733 ( .A(n664), .B(n663), .ZN(G57) );
  XNOR2_X1 U734 ( .A(n665), .B(G134), .ZN(G36) );
  XOR2_X1 U735 ( .A(n666), .B(G110), .Z(G12) );
  NAND2_X1 U736 ( .A1(n760), .A2(n755), .ZN(n668) );
  XOR2_X1 U737 ( .A(G113), .B(KEYINPUT113), .Z(n667) );
  XNOR2_X1 U738 ( .A(n668), .B(n667), .ZN(G15) );
  XOR2_X1 U739 ( .A(G131), .B(KEYINPUT127), .Z(n669) );
  XNOR2_X1 U740 ( .A(n670), .B(n669), .ZN(G33) );
  XNOR2_X1 U741 ( .A(G122), .B(KEYINPUT126), .ZN(n671) );
  XNOR2_X1 U742 ( .A(n672), .B(n671), .ZN(G24) );
  NAND2_X1 U743 ( .A1(n673), .A2(G217), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n676), .A2(n696), .ZN(G66) );
  NAND2_X1 U746 ( .A1(n673), .A2(G478), .ZN(n677) );
  XOR2_X1 U747 ( .A(n678), .B(n677), .Z(n679) );
  NOR2_X1 U748 ( .A1(n679), .A2(n696), .ZN(G63) );
  NAND2_X1 U749 ( .A1(n691), .A2(G475), .ZN(n682) );
  XNOR2_X1 U750 ( .A(n684), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U751 ( .A1(n691), .A2(G469), .ZN(n688) );
  XNOR2_X1 U752 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n685) );
  XNOR2_X1 U753 ( .A(n685), .B(KEYINPUT58), .ZN(n686) );
  XNOR2_X1 U754 ( .A(n688), .B(n367), .ZN(n689) );
  XNOR2_X1 U755 ( .A(n690), .B(KEYINPUT122), .ZN(G54) );
  NAND2_X1 U756 ( .A1(n691), .A2(G210), .ZN(n695) );
  XNOR2_X1 U757 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n692) );
  XNOR2_X1 U758 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U759 ( .A(n698), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X1 U760 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U761 ( .A(n701), .B(KEYINPUT80), .ZN(n738) );
  INV_X1 U762 ( .A(n702), .ZN(n733) );
  NOR2_X1 U763 ( .A1(n595), .A2(n703), .ZN(n704) );
  NOR2_X1 U764 ( .A1(n705), .A2(n704), .ZN(n710) );
  NOR2_X1 U765 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U766 ( .A(n708), .B(KEYINPUT118), .ZN(n709) );
  NOR2_X1 U767 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U768 ( .A1(n733), .A2(n711), .ZN(n728) );
  NOR2_X1 U769 ( .A1(n713), .A2(n712), .ZN(n715) );
  XNOR2_X1 U770 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n714) );
  XNOR2_X1 U771 ( .A(n715), .B(n714), .ZN(n716) );
  AND2_X1 U772 ( .A1(n716), .A2(n582), .ZN(n722) );
  NOR2_X1 U773 ( .A1(n718), .A2(n717), .ZN(n720) );
  XNOR2_X1 U774 ( .A(KEYINPUT117), .B(KEYINPUT50), .ZN(n719) );
  XNOR2_X1 U775 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U776 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U777 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U778 ( .A(n725), .B(KEYINPUT51), .ZN(n726) );
  NOR2_X1 U779 ( .A1(n726), .A2(n732), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U781 ( .A(KEYINPUT52), .B(n729), .Z(n731) );
  NAND2_X1 U782 ( .A1(n731), .A2(n730), .ZN(n736) );
  NOR2_X1 U783 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U784 ( .A1(n734), .A2(G953), .ZN(n735) );
  NAND2_X1 U785 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U786 ( .A1(n738), .A2(n737), .ZN(n741) );
  XNOR2_X1 U787 ( .A(KEYINPUT120), .B(KEYINPUT53), .ZN(n739) );
  XOR2_X1 U788 ( .A(n739), .B(KEYINPUT119), .Z(n740) );
  XNOR2_X1 U789 ( .A(n741), .B(n740), .ZN(G75) );
  XNOR2_X1 U790 ( .A(n742), .B(G104), .ZN(G6) );
  XNOR2_X1 U791 ( .A(n373), .B(KEYINPUT27), .ZN(n746) );
  XOR2_X1 U792 ( .A(KEYINPUT108), .B(KEYINPUT26), .Z(n744) );
  XNOR2_X1 U793 ( .A(n744), .B(n743), .ZN(n745) );
  XNOR2_X1 U794 ( .A(n746), .B(n745), .ZN(G9) );
  INV_X1 U795 ( .A(n756), .ZN(n748) );
  NOR2_X1 U796 ( .A1(n748), .A2(n747), .ZN(n752) );
  XOR2_X1 U797 ( .A(KEYINPUT109), .B(KEYINPUT29), .Z(n750) );
  XNOR2_X1 U798 ( .A(G128), .B(KEYINPUT110), .ZN(n749) );
  XNOR2_X1 U799 ( .A(n750), .B(n749), .ZN(n751) );
  XNOR2_X1 U800 ( .A(n752), .B(n751), .ZN(G30) );
  XOR2_X1 U801 ( .A(G143), .B(KEYINPUT111), .Z(n753) );
  XNOR2_X1 U802 ( .A(n754), .B(n753), .ZN(G45) );
  NAND2_X1 U803 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U804 ( .A(n757), .B(KEYINPUT112), .ZN(n758) );
  XNOR2_X1 U805 ( .A(G146), .B(n758), .ZN(G48) );
  NAND2_X1 U806 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U807 ( .A(n761), .B(KEYINPUT114), .ZN(n762) );
  XNOR2_X1 U808 ( .A(G116), .B(n762), .ZN(G18) );
  XOR2_X1 U809 ( .A(G140), .B(KEYINPUT115), .Z(n763) );
  XNOR2_X1 U810 ( .A(n764), .B(n763), .ZN(G42) );
  NAND2_X1 U811 ( .A1(n765), .A2(n771), .ZN(n769) );
  NAND2_X1 U812 ( .A1(G953), .A2(G224), .ZN(n766) );
  XNOR2_X1 U813 ( .A(KEYINPUT61), .B(n766), .ZN(n767) );
  NAND2_X1 U814 ( .A1(n767), .A2(G898), .ZN(n768) );
  NAND2_X1 U815 ( .A1(n769), .A2(n768), .ZN(n774) );
  NOR2_X1 U816 ( .A1(G898), .A2(n771), .ZN(n772) );
  NOR2_X1 U817 ( .A1(n770), .A2(n772), .ZN(n773) );
  XNOR2_X1 U818 ( .A(n774), .B(n773), .ZN(G69) );
  XNOR2_X1 U819 ( .A(n775), .B(KEYINPUT123), .ZN(n776) );
  XNOR2_X1 U820 ( .A(n777), .B(n776), .ZN(n782) );
  XOR2_X1 U821 ( .A(KEYINPUT124), .B(n782), .Z(n778) );
  XNOR2_X1 U822 ( .A(n779), .B(n778), .ZN(n780) );
  NOR2_X1 U823 ( .A1(n780), .A2(G953), .ZN(n781) );
  XNOR2_X1 U824 ( .A(n781), .B(KEYINPUT125), .ZN(n786) );
  XNOR2_X1 U825 ( .A(n782), .B(G227), .ZN(n783) );
  NAND2_X1 U826 ( .A1(n783), .A2(G900), .ZN(n784) );
  NAND2_X1 U827 ( .A1(G953), .A2(n784), .ZN(n785) );
  NAND2_X1 U828 ( .A1(n786), .A2(n785), .ZN(G72) );
  XNOR2_X1 U829 ( .A(n787), .B(G125), .ZN(n788) );
  XNOR2_X1 U830 ( .A(n788), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U831 ( .A(G101), .B(n789), .ZN(G3) );
  XNOR2_X1 U832 ( .A(G137), .B(n790), .ZN(G39) );
endmodule

