//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  XNOR2_X1  g000(.A(G110), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G107), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G104), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G101), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT74), .ZN(new_n193));
  AOI21_X1  g007(.A(KEYINPUT3), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n193), .A2(new_n188), .A3(KEYINPUT3), .A4(G104), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n190), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n193), .A2(new_n188), .A3(G104), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n189), .B1(new_n200), .B2(new_n195), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n197), .B(KEYINPUT4), .C1(new_n201), .C2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n195), .ZN(new_n204));
  INV_X1    g018(.A(new_n189), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n202), .A2(KEYINPUT4), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(G116), .B(G119), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT2), .B(G113), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n203), .A2(new_n208), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n209), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(new_n210), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT5), .ZN(new_n216));
  INV_X1    g030(.A(G119), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G116), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT80), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT80), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n220), .A2(new_n216), .A3(new_n217), .A4(G116), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(G113), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n209), .A2(KEYINPUT5), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n215), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G104), .B(G107), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT76), .B1(new_n226), .B2(new_n202), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT76), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n228), .B(G101), .C1(new_n189), .C2(new_n192), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n227), .A2(new_n229), .B1(new_n204), .B2(new_n190), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n187), .B1(new_n213), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT6), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT81), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n213), .A2(new_n231), .A3(new_n187), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT6), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n234), .B(new_n235), .C1(new_n237), .C2(new_n232), .ZN(new_n238));
  INV_X1    g052(.A(new_n232), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n239), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n236), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n242));
  XNOR2_X1  g056(.A(G143), .B(G146), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT0), .B(G128), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G143), .ZN(new_n247));
  INV_X1    g061(.A(G143), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G146), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  NOR2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n253), .A3(KEYINPUT64), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n247), .A2(new_n249), .A3(new_n251), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT65), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT65), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n247), .A2(new_n249), .A3(new_n251), .A4(new_n257), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n245), .A2(new_n254), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G125), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT1), .B1(new_n248), .B2(G146), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n250), .A2(G128), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G128), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n247), .B(new_n249), .C1(KEYINPUT1), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n261), .B1(new_n260), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G224), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(G953), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n267), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n241), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G210), .B1(G237), .B2(G902), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n273), .B(KEYINPUT84), .Z(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n269), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n276), .A2(KEYINPUT7), .ZN(new_n277));
  INV_X1    g091(.A(new_n261), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n278), .B2(KEYINPUT83), .ZN(new_n279));
  INV_X1    g093(.A(new_n266), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n278), .B1(G125), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OAI221_X1 g096(.A(new_n278), .B1(KEYINPUT83), .B2(new_n277), .C1(G125), .C2(new_n280), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n227), .A2(new_n229), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n197), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n225), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n187), .B(KEYINPUT8), .ZN(new_n287));
  OR2_X1    g101(.A1(new_n222), .A2(KEYINPUT82), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n222), .A2(KEYINPUT82), .B1(KEYINPUT5), .B2(new_n209), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n215), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n286), .B(new_n287), .C1(new_n290), .C2(new_n285), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n282), .A2(new_n283), .A3(new_n236), .A4(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n272), .A2(new_n275), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT85), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n270), .B1(new_n238), .B2(new_n240), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n293), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n274), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n295), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  OAI211_X1 g114(.A(KEYINPUT85), .B(new_n274), .C1(new_n297), .C2(new_n298), .ZN(new_n301));
  OAI21_X1  g115(.A(G214), .B1(G237), .B2(G902), .ZN(new_n302));
  INV_X1    g116(.A(G122), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT88), .B1(new_n303), .B2(G116), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT88), .ZN(new_n305));
  INV_X1    g119(.A(G116), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(G122), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT14), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n303), .A2(G116), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n308), .A2(KEYINPUT14), .ZN(new_n312));
  OAI21_X1  g126(.A(G107), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT89), .B1(new_n264), .B2(G143), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT89), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n248), .A3(G128), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n264), .A2(G143), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G134), .ZN(new_n320));
  INV_X1    g134(.A(G134), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n317), .A2(new_n321), .A3(new_n318), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n308), .A2(new_n188), .A3(new_n310), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n313), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT90), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT13), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n317), .B2(new_n327), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT90), .A4(KEYINPUT13), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n317), .A2(new_n327), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n328), .A2(new_n318), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n331), .A2(G134), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n308), .A2(new_n310), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G107), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n324), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n317), .A2(KEYINPUT91), .A3(new_n321), .A4(new_n318), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT91), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n322), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n325), .B1(new_n332), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT9), .B(G234), .ZN(new_n341));
  INV_X1    g155(.A(G217), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n341), .A2(new_n342), .A3(G953), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n331), .A2(G134), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n346), .A2(new_n336), .A3(new_n335), .A4(new_n338), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n325), .A3(new_n343), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n293), .ZN(new_n350));
  INV_X1    g164(.A(G478), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT92), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(KEYINPUT15), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(KEYINPUT15), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n356), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n349), .A2(new_n293), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(G125), .B(G140), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT16), .ZN(new_n362));
  OR3_X1    g176(.A1(new_n260), .A2(KEYINPUT16), .A3(G140), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n362), .A2(G146), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(G146), .B1(new_n362), .B2(new_n363), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G237), .ZN(new_n367));
  INV_X1    g181(.A(G953), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(G214), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT86), .A3(new_n248), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n248), .A2(KEYINPUT86), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n371), .A2(G214), .A3(new_n367), .A4(new_n368), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT66), .B(G131), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT17), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n370), .A2(new_n372), .A3(new_n374), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n373), .A2(KEYINPUT17), .A3(new_n375), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n366), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(KEYINPUT18), .A2(G131), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n370), .A2(new_n372), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n373), .A2(KEYINPUT18), .A3(G131), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n361), .A2(new_n246), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n361), .A2(new_n246), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT87), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n361), .A2(new_n246), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT87), .B1(new_n390), .B2(new_n385), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n383), .B(new_n384), .C1(new_n389), .C2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G113), .B(G122), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(new_n191), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n381), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n394), .B1(new_n381), .B2(new_n392), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n293), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G475), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n381), .A2(new_n392), .A3(new_n394), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n362), .A2(G146), .A3(new_n363), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT72), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n362), .A2(KEYINPUT72), .A3(G146), .A4(new_n363), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n361), .B(KEYINPUT19), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n376), .A2(new_n378), .B1(new_n405), .B2(new_n246), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n384), .A2(new_n383), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n388), .B1(new_n386), .B2(new_n387), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n390), .A2(new_n385), .A3(KEYINPUT87), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n404), .A2(new_n406), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n399), .B1(new_n411), .B2(new_n394), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n413));
  NOR2_X1   g227(.A1(G475), .A2(G902), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n413), .B1(new_n412), .B2(new_n414), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n398), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n368), .A2(G952), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n418), .B1(G234), .B2(G237), .ZN(new_n419));
  AOI211_X1 g233(.A(new_n293), .B(new_n368), .C1(G234), .C2(G237), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT21), .B(G898), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n360), .A2(new_n417), .A3(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n300), .A2(new_n301), .A3(new_n302), .A4(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G221), .B1(new_n341), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(G469), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT12), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n285), .A2(new_n266), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n230), .A2(new_n280), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT11), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n321), .B2(G137), .ZN(new_n432));
  INV_X1    g246(.A(G137), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(KEYINPUT11), .A3(G134), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n321), .A2(G137), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G131), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n374), .A2(new_n432), .A3(new_n434), .A4(new_n435), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n427), .B1(new_n430), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n440), .B1(new_n428), .B2(new_n429), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT12), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n197), .A2(KEYINPUT4), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n202), .B1(new_n204), .B2(new_n205), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n259), .B(new_n208), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT75), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT75), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n203), .A2(new_n449), .A3(new_n208), .A4(new_n259), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT67), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n262), .A2(G128), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(new_n243), .ZN(new_n454));
  INV_X1    g268(.A(new_n265), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n263), .A2(KEYINPUT67), .A3(new_n265), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n230), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT10), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT10), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n230), .A2(new_n460), .A3(new_n280), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n451), .A2(new_n440), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n444), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G110), .B(G140), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n368), .A2(G227), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n467), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n463), .A2(KEYINPUT77), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n451), .A2(new_n462), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n439), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT77), .B1(new_n463), .B2(new_n469), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n426), .B1(new_n475), .B2(new_n293), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT78), .B(G469), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n472), .A2(new_n463), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n467), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n448), .A2(new_n450), .B1(new_n459), .B2(new_n461), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n467), .B1(new_n481), .B2(new_n440), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n442), .A2(KEYINPUT12), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n427), .B(new_n440), .C1(new_n428), .C2(new_n429), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT79), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT79), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n441), .A2(new_n486), .A3(new_n443), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  AOI211_X1 g302(.A(G902), .B(new_n478), .C1(new_n480), .C2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n425), .B1(new_n476), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT93), .ZN(new_n491));
  OR3_X1    g305(.A1(new_n424), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n491), .B1(new_n424), .B2(new_n490), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n342), .B1(G234), .B2(new_n293), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT71), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT70), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n497), .B(KEYINPUT23), .C1(new_n264), .C2(G119), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n217), .A2(G128), .ZN(new_n499));
  OR2_X1    g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n498), .B(new_n499), .C1(new_n497), .C2(KEYINPUT23), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G110), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT24), .B(G110), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT69), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n264), .B2(G119), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n217), .A2(KEYINPUT69), .A3(G128), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n499), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n506), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n496), .B1(new_n504), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(G110), .B1(new_n500), .B2(new_n501), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n515), .A2(KEYINPUT71), .A3(new_n512), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n385), .B(new_n404), .C1(new_n514), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n510), .A2(new_n511), .ZN(new_n518));
  OAI22_X1  g332(.A1(new_n502), .A2(new_n503), .B1(new_n518), .B2(new_n505), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(new_n366), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n368), .A2(G221), .A3(G234), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT73), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT22), .B(G137), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n517), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n525), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n402), .A2(new_n385), .A3(new_n403), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n504), .A2(new_n496), .A3(new_n513), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT71), .B1(new_n515), .B2(new_n512), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n527), .B1(new_n531), .B2(new_n520), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n526), .A2(new_n293), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT25), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n526), .A2(new_n532), .A3(KEYINPUT25), .A4(new_n293), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n495), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n526), .A2(new_n532), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n494), .A2(G902), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n259), .A2(new_n439), .ZN(new_n543));
  INV_X1    g357(.A(new_n435), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n321), .A2(G137), .ZN(new_n545));
  OAI21_X1  g359(.A(G131), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n438), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n280), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n456), .A2(new_n547), .A3(new_n457), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n543), .A3(KEYINPUT30), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n212), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n543), .A3(new_n211), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n367), .A2(new_n368), .A3(G210), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT27), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT26), .B(G101), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n554), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT31), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT31), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n554), .A2(new_n562), .A3(new_n555), .A4(new_n559), .ZN(new_n563));
  INV_X1    g377(.A(new_n555), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(KEYINPUT28), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n439), .A2(new_n259), .B1(new_n280), .B2(new_n547), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT68), .B1(new_n566), .B2(new_n211), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT68), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n549), .A2(new_n568), .A3(new_n212), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n569), .A3(new_n555), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n565), .B1(new_n570), .B2(KEYINPUT28), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n561), .B(new_n563), .C1(new_n571), .C2(new_n559), .ZN(new_n572));
  NOR2_X1   g386(.A1(G472), .A2(G902), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT32), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT32), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n572), .A2(new_n576), .A3(new_n573), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G472), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n571), .A2(new_n559), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n554), .A2(new_n555), .ZN(new_n581));
  INV_X1    g395(.A(new_n559), .ZN(new_n582));
  AOI21_X1  g396(.A(KEYINPUT29), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n211), .B1(new_n552), .B2(new_n543), .ZN(new_n585));
  OR2_X1    g399(.A1(new_n564), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n565), .B1(new_n586), .B2(KEYINPUT28), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n559), .A2(KEYINPUT29), .ZN(new_n588));
  AOI21_X1  g402(.A(G902), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n579), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n542), .B1(new_n578), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n492), .A2(new_n493), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT94), .B(G101), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G3));
  NAND2_X1  g409(.A1(new_n561), .A2(new_n563), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n570), .A2(KEYINPUT28), .ZN(new_n597));
  INV_X1    g411(.A(new_n565), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n559), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n293), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G472), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n574), .A3(new_n541), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT95), .B1(new_n490), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n425), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n469), .B1(new_n444), .B2(new_n463), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n440), .B1(new_n451), .B2(new_n462), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n482), .B2(KEYINPUT77), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n463), .A2(new_n469), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT77), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n605), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(G469), .B1(new_n611), .B2(G902), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n469), .B1(new_n472), .B2(new_n463), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n293), .B(new_n477), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n604), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT95), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n579), .B1(new_n572), .B2(new_n293), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n572), .B2(new_n573), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n616), .A2(new_n617), .A3(new_n619), .A4(new_n541), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n603), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n275), .B1(new_n272), .B2(new_n294), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n297), .A2(new_n298), .A3(new_n274), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n302), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n293), .A2(G478), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT96), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n626), .A2(KEYINPUT96), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n349), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n345), .A2(new_n348), .A3(KEYINPUT96), .A4(new_n626), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(G478), .B1(new_n349), .B2(new_n293), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n417), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n624), .A2(new_n633), .A3(new_n422), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n621), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  INV_X1    g451(.A(new_n302), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n295), .B2(new_n299), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n412), .A2(new_n414), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT20), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n641), .A2(new_n642), .B1(G475), .B2(new_n397), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n360), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n422), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n621), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT97), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(new_n619), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n517), .A2(new_n521), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n527), .A2(KEYINPUT36), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n654), .A2(new_n539), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n537), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n492), .A2(new_n493), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT37), .B(G110), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  AOI21_X1  g476(.A(new_n656), .B1(new_n578), .B2(new_n591), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n358), .B1(new_n349), .B2(new_n293), .ZN(new_n664));
  AOI211_X1 g478(.A(G902), .B(new_n356), .C1(new_n345), .C2(new_n348), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n417), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n420), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n419), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(KEYINPUT100), .B1(new_n624), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n671), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n644), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n639), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n663), .A2(new_n673), .A3(new_n616), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  XOR2_X1   g493(.A(new_n671), .B(KEYINPUT39), .Z(new_n680));
  OAI21_X1  g494(.A(KEYINPUT40), .B1(new_n490), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n300), .A2(new_n301), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n682), .B(new_n684), .ZN(new_n685));
  OR3_X1    g499(.A1(new_n490), .A2(KEYINPUT40), .A3(new_n680), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n293), .B1(new_n586), .B2(new_n559), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n581), .A2(new_n559), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n579), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n575), .B2(new_n577), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n643), .A2(new_n666), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n302), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n655), .A2(new_n537), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT102), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT102), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n656), .A2(new_n692), .A3(new_n696), .A4(new_n302), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n691), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  AND4_X1   g512(.A1(new_n681), .A2(new_n685), .A3(new_n686), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n248), .ZN(G45));
  OAI211_X1 g514(.A(new_n417), .B(new_n671), .C1(new_n631), .C2(new_n632), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n624), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n663), .A2(new_n616), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  AOI21_X1  g518(.A(new_n590), .B1(new_n575), .B2(new_n577), .ZN(new_n705));
  AOI21_X1  g519(.A(G902), .B1(new_n480), .B2(new_n488), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n615), .B(new_n425), .C1(new_n706), .C2(new_n426), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n705), .A2(new_n542), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n634), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND2_X1  g525(.A1(new_n708), .A2(new_n646), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT103), .B(G116), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G18));
  INV_X1    g528(.A(new_n423), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n707), .A2(new_n624), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n663), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  OAI211_X1 g532(.A(new_n561), .B(new_n563), .C1(new_n587), .C2(new_n559), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n573), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n601), .A2(KEYINPUT104), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n618), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n541), .B(new_n720), .C1(new_n721), .C2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT105), .B1(new_n643), .B2(new_n666), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n360), .A2(new_n727), .A3(new_n417), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n707), .A2(new_n624), .A3(new_n729), .A4(new_n422), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT106), .B(G122), .Z(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G24));
  INV_X1    g547(.A(new_n720), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n601), .A2(KEYINPUT104), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n618), .A2(new_n722), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n707), .A2(new_n624), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n701), .B(KEYINPUT107), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n737), .A2(new_n738), .A3(new_n739), .A4(new_n694), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  AOI21_X1  g555(.A(new_n638), .B1(new_n300), .B2(new_n301), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n592), .A2(new_n616), .A3(new_n739), .A4(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n682), .A2(new_n302), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n490), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(KEYINPUT42), .A3(new_n592), .A4(new_n739), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT108), .B(G131), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G33));
  INV_X1    g565(.A(new_n592), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n752), .A2(new_n490), .A3(new_n746), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n675), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  NAND2_X1  g569(.A1(new_n611), .A2(KEYINPUT45), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n426), .B1(new_n475), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n761));
  AOI211_X1 g575(.A(KEYINPUT109), .B(new_n426), .C1(new_n475), .C2(new_n757), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n475), .A2(new_n757), .ZN(new_n764));
  OAI21_X1  g578(.A(G469), .B1(new_n611), .B2(KEYINPUT45), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n764), .B1(new_n765), .B2(KEYINPUT109), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n758), .A2(new_n759), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT110), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI22_X1  g582(.A1(new_n763), .A2(new_n768), .B1(new_n426), .B2(new_n293), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT46), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n426), .A2(new_n293), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n770), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(new_n763), .B2(new_n768), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n761), .B1(new_n760), .B2(new_n762), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n766), .A2(KEYINPUT110), .A3(new_n767), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(KEYINPUT111), .A3(new_n773), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n771), .A2(new_n776), .A3(new_n615), .A4(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n680), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n631), .A2(new_n632), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n417), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT43), .Z(new_n786));
  NAND2_X1  g600(.A1(new_n651), .A2(new_n694), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n742), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n786), .A2(new_n787), .A3(new_n783), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n781), .A2(new_n425), .A3(new_n782), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  AOI21_X1  g607(.A(new_n772), .B1(new_n777), .B2(new_n778), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n615), .B1(new_n794), .B2(KEYINPUT46), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT111), .B1(new_n779), .B2(new_n773), .ZN(new_n796));
  INV_X1    g610(.A(new_n773), .ZN(new_n797));
  AOI211_X1 g611(.A(new_n775), .B(new_n797), .C1(new_n777), .C2(new_n778), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n795), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT47), .B1(new_n799), .B2(new_n604), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n781), .A2(new_n801), .A3(new_n425), .ZN(new_n802));
  INV_X1    g616(.A(new_n705), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n746), .A2(new_n803), .A3(new_n541), .A4(new_n701), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n800), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  OR2_X1    g620(.A1(G952), .A2(G953), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n786), .A2(new_n670), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n746), .A2(new_n707), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n592), .A3(new_n809), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n810), .B(KEYINPUT48), .Z(new_n811));
  XOR2_X1   g625(.A(new_n418), .B(KEYINPUT118), .Z(new_n812));
  NAND4_X1  g626(.A1(new_n809), .A2(new_n419), .A3(new_n541), .A4(new_n691), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n808), .A2(new_n725), .ZN(new_n814));
  INV_X1    g628(.A(new_n738), .ZN(new_n815));
  OAI221_X1 g629(.A(new_n812), .B1(new_n813), .B2(new_n633), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n615), .B1(new_n706), .B2(new_n426), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(new_n425), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n796), .A2(new_n798), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n489), .B1(new_n769), .B2(new_n770), .ZN(new_n822));
  AOI211_X1 g636(.A(KEYINPUT47), .B(new_n604), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n801), .B1(new_n781), .B2(new_n425), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n814), .A2(new_n746), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n682), .B(new_n683), .ZN(new_n828));
  NOR2_X1   g642(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n707), .A2(new_n302), .A3(new_n829), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n828), .A2(new_n808), .A3(new_n725), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n784), .A2(new_n643), .ZN(new_n835));
  OR3_X1    g649(.A1(new_n813), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n834), .B1(new_n813), .B2(new_n835), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n808), .A2(new_n694), .A3(new_n737), .A4(new_n809), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n831), .A2(new_n832), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n833), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n818), .B1(new_n827), .B2(new_n842), .ZN(new_n843));
  AOI211_X1 g657(.A(KEYINPUT51), .B(new_n841), .C1(new_n825), .C2(new_n826), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n817), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n725), .A2(new_n730), .B1(new_n708), .B2(new_n646), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n708), .A2(new_n634), .B1(new_n716), .B2(new_n663), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n300), .A2(new_n301), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(KEYINPUT112), .A3(new_n302), .A4(new_n645), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n645), .A2(new_n300), .A3(new_n302), .A4(new_n301), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT112), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n850), .A2(new_n603), .A3(new_n620), .A4(new_n853), .ZN(new_n854));
  NOR4_X1   g668(.A1(new_n682), .A2(new_n638), .A3(new_n633), .A4(new_n422), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n603), .A3(new_n620), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n847), .A2(new_n848), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n492), .B(new_n493), .C1(new_n592), .C2(new_n657), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT113), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n360), .A2(new_n417), .A3(new_n674), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n682), .A2(new_n861), .A3(new_n302), .A4(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n863), .A2(new_n616), .A3(new_n663), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n742), .A2(new_n862), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT113), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n737), .A2(new_n694), .A3(new_n739), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n864), .A2(new_n866), .B1(new_n867), .B2(new_n747), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n868), .A2(new_n749), .A3(new_n754), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n678), .A2(new_n740), .A3(new_n703), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n624), .A2(new_n729), .A3(new_n694), .A4(new_n674), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  INV_X1    g686(.A(new_n690), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n578), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n871), .A2(new_n872), .A3(new_n616), .A4(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n624), .A2(new_n729), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n694), .A2(new_n674), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n874), .A2(new_n876), .A3(new_n616), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT114), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n870), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT52), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT52), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n870), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n860), .A2(new_n869), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n846), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n881), .B1(new_n678), .B2(new_n740), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n886), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n854), .A2(new_n856), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(new_n848), .A3(new_n847), .A4(new_n858), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n868), .A2(new_n749), .A3(new_n754), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n883), .B1(new_n870), .B2(new_n880), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n894), .A2(KEYINPUT115), .A3(KEYINPUT53), .A4(new_n884), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n887), .A2(new_n889), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT54), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT53), .B1(new_n885), .B2(new_n888), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n894), .A2(new_n886), .A3(new_n884), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT54), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n807), .B1(new_n845), .B2(new_n902), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n542), .A2(new_n604), .A3(new_n638), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n819), .A2(KEYINPUT49), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n905), .A3(new_n785), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n819), .A2(KEYINPUT49), .ZN(new_n907));
  OR4_X1    g721(.A1(new_n685), .A2(new_n906), .A3(new_n874), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n903), .A2(new_n908), .ZN(G75));
  NAND4_X1  g723(.A1(new_n898), .A2(G902), .A3(new_n899), .A4(new_n274), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT56), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n241), .A2(new_n271), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n297), .ZN(new_n913));
  XNOR2_X1  g727(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT120), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n913), .B(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n910), .A2(new_n911), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n916), .B1(new_n910), .B2(new_n911), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n368), .A2(G952), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(G51));
  XNOR2_X1  g734(.A(new_n772), .B(KEYINPUT57), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n898), .A2(KEYINPUT54), .A3(new_n899), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(new_n900), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(new_n614), .B2(new_n613), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n898), .A2(new_n899), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n925), .A2(G902), .A3(new_n777), .A4(new_n778), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n919), .B1(new_n924), .B2(new_n926), .ZN(G54));
  NAND2_X1  g741(.A1(KEYINPUT58), .A2(G475), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT121), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n925), .A2(G902), .A3(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n412), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n932), .A2(new_n933), .A3(new_n919), .ZN(G60));
  NAND2_X1  g748(.A1(new_n629), .A2(new_n630), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(G478), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT59), .Z(new_n938));
  NOR2_X1   g752(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n922), .B2(new_n900), .ZN(new_n940));
  INV_X1    g754(.A(new_n919), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n938), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n902), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n942), .B1(new_n936), .B2(new_n944), .ZN(G63));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT60), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n925), .A2(new_n654), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n898), .A2(new_n899), .A3(new_n948), .ZN(new_n950));
  INV_X1    g764(.A(new_n538), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n949), .A2(new_n941), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n949), .A2(KEYINPUT61), .A3(new_n941), .A4(new_n952), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(G66));
  OAI21_X1  g771(.A(G953), .B1(new_n421), .B2(new_n268), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n860), .B(KEYINPUT122), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n958), .B1(new_n960), .B2(G953), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n238), .B(new_n240), .C1(G898), .C2(new_n368), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  NAND2_X1  g777(.A1(new_n749), .A2(new_n754), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n678), .A2(new_n740), .A3(new_n703), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n678), .A2(new_n740), .A3(new_n703), .A4(KEYINPUT123), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n792), .A2(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n592), .A2(new_n876), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n781), .A2(new_n425), .A3(new_n782), .A4(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n970), .A2(new_n805), .A3(new_n368), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n551), .A2(new_n553), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(new_n405), .Z(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(G900), .B2(G953), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT125), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n368), .B1(G227), .B2(G900), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n699), .B1(new_n967), .B2(new_n968), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n680), .B1(new_n633), .B2(new_n644), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n753), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n792), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n967), .A2(new_n968), .ZN(new_n989));
  INV_X1    g803(.A(new_n699), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT124), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n983), .B2(new_n984), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n988), .A2(new_n805), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n975), .B1(new_n996), .B2(new_n368), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n973), .A2(new_n977), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n980), .B(new_n982), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n996), .A2(new_n368), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n976), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n1001), .B(new_n978), .C1(new_n979), .C2(new_n981), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n999), .A2(new_n1002), .ZN(G72));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  NAND3_X1  g819(.A1(new_n970), .A2(new_n805), .A3(new_n972), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1005), .B1(new_n1006), .B2(new_n959), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n581), .A2(new_n559), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n919), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1005), .B1(new_n996), .B2(new_n959), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1010), .A2(new_n559), .A3(new_n581), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT127), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1008), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1014), .A2(new_n689), .A3(new_n1005), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT126), .Z(new_n1016));
  AND3_X1   g830(.A1(new_n896), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1013), .B1(new_n896), .B2(new_n1016), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1012), .A2(new_n1019), .ZN(G57));
endmodule


