//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G104), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  AOI21_X1  g006(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(G107), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G101), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n197), .B(new_n191), .C1(new_n193), .C2(new_n194), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(KEYINPUT4), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n201), .A2(new_n203), .A3(G128), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT64), .B1(new_n202), .B2(G146), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n200), .A3(G143), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n207), .A3(new_n203), .ZN(new_n208));
  XOR2_X1   g022(.A(KEYINPUT0), .B(G128), .Z(new_n209));
  AOI22_X1  g023(.A1(KEYINPUT0), .A2(new_n204), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT4), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n195), .A2(new_n211), .A3(G101), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n199), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n214));
  OR2_X1    g028(.A1(KEYINPUT67), .A2(G128), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT67), .A2(G128), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n208), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n201), .A2(new_n203), .A3(new_n219), .A4(G128), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n190), .A2(G104), .ZN(new_n222));
  OAI21_X1  g036(.A(G101), .B1(new_n194), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n198), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n224), .A3(KEYINPUT10), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n213), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n214), .A2(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n201), .A2(new_n203), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n204), .A2(new_n219), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n198), .A2(new_n223), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT80), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G128), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n234));
  XNOR2_X1  g048(.A(G143), .B(G146), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n220), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT80), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n236), .A2(new_n237), .A3(new_n198), .A4(new_n223), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT10), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT11), .A2(G134), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(KEYINPUT65), .A2(G137), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT65), .A2(G137), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT66), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT65), .B(G137), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(new_n243), .ZN(new_n250));
  INV_X1    g064(.A(G137), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n251), .B1(KEYINPUT11), .B2(G134), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n242), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n247), .A2(new_n250), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G131), .ZN(new_n255));
  INV_X1    g069(.A(G131), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n247), .A2(new_n250), .A3(new_n256), .A4(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n227), .A2(new_n241), .A3(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G110), .B(G140), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n262), .A2(G227), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n261), .B(new_n263), .Z(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n218), .A2(new_n220), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n231), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n237), .B1(new_n224), .B2(new_n236), .ZN(new_n268));
  AND4_X1   g082(.A1(new_n237), .A2(new_n236), .A3(new_n198), .A4(new_n223), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT82), .ZN(new_n271));
  XOR2_X1   g085(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n270), .A2(new_n271), .A3(new_n258), .A4(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT12), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n232), .A2(new_n238), .B1(new_n266), .B2(new_n231), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(new_n259), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n239), .A2(new_n267), .B1(new_n255), .B2(new_n257), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n271), .B1(new_n279), .B2(new_n273), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n265), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT83), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n227), .A2(new_n241), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT10), .B1(new_n232), .B2(new_n238), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT83), .B1(new_n285), .B2(new_n226), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n258), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n264), .B1(new_n287), .B2(new_n260), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n187), .B(new_n188), .C1(new_n282), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n274), .A2(new_n277), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n260), .B1(new_n290), .B2(new_n280), .ZN(new_n291));
  INV_X1    g105(.A(new_n264), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n287), .A2(new_n264), .A3(new_n260), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(G469), .A3(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n187), .A2(new_n188), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n289), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G221), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT9), .B(G234), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n299), .B1(new_n301), .B2(new_n188), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT84), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT84), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n298), .A2(new_n306), .A3(new_n303), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(G237), .A2(G953), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G214), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(new_n202), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT18), .A3(G131), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n310), .A2(new_n202), .ZN(new_n313));
  AOI21_X1  g127(.A(G143), .B1(new_n309), .B2(G214), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(KEYINPUT18), .A2(G131), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G125), .ZN(new_n318));
  OAI21_X1  g132(.A(G140), .B1(new_n318), .B2(KEYINPUT75), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G146), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(G125), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n318), .A2(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n200), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n312), .A2(new_n317), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n311), .A2(G131), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n315), .A2(new_n256), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT17), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n321), .B1(new_n320), .B2(G125), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n318), .A2(KEYINPUT75), .A3(G140), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT16), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT16), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n325), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n200), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n337), .B1(new_n319), .B2(new_n322), .ZN(new_n340));
  INV_X1    g154(.A(new_n338), .ZN(new_n341));
  OAI21_X1  g155(.A(G146), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n339), .B(new_n342), .C1(new_n330), .C2(new_n332), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n329), .B1(new_n333), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G113), .B(G122), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(new_n192), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n317), .A2(new_n328), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(new_n312), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n323), .A2(KEYINPUT19), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT19), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n325), .A2(new_n326), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n200), .A3(new_n351), .ZN(new_n352));
  OR2_X1    g166(.A1(new_n352), .A2(KEYINPUT89), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n330), .A2(new_n331), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(KEYINPUT89), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n353), .A2(new_n354), .A3(new_n342), .A4(new_n355), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n344), .A2(new_n346), .B1(new_n348), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT20), .ZN(new_n358));
  NOR2_X1   g172(.A1(G475), .A2(G902), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT90), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n357), .A2(KEYINPUT90), .A3(new_n358), .A4(new_n359), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n357), .A2(new_n359), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT20), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  OR2_X1    g180(.A1(new_n346), .A2(KEYINPUT91), .ZN(new_n367));
  AOI21_X1  g181(.A(G902), .B1(new_n344), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(new_n367), .B2(new_n344), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G475), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT92), .ZN(new_n372));
  INV_X1    g186(.A(G122), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G116), .ZN(new_n374));
  INV_X1    g188(.A(G116), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G122), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n190), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n376), .A3(G107), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AND2_X1   g194(.A1(KEYINPUT67), .A2(G128), .ZN(new_n381));
  NOR2_X1   g195(.A1(KEYINPUT67), .A2(G128), .ZN(new_n382));
  OAI21_X1  g196(.A(G143), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G134), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n202), .A2(G128), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n383), .A2(KEYINPUT13), .A3(new_n385), .ZN(new_n387));
  OAI21_X1  g201(.A(G134), .B1(new_n385), .B2(KEYINPUT13), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n380), .B(new_n386), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n374), .A2(KEYINPUT14), .A3(G107), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n378), .A2(new_n379), .A3(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT14), .A4(G107), .ZN(new_n392));
  INV_X1    g206(.A(new_n386), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n384), .B1(new_n383), .B2(new_n385), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n391), .B(new_n392), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G217), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n300), .A2(new_n396), .A3(G953), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n389), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n397), .B1(new_n389), .B2(new_n395), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n372), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n399), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT92), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n188), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT15), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G478), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(KEYINPUT93), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(G902), .B1(new_n400), .B2(new_n402), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT93), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n405), .B(G478), .C1(new_n408), .C2(new_n409), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n407), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(G234), .A2(G237), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(G952), .A3(new_n262), .ZN(new_n415));
  XOR2_X1   g229(.A(KEYINPUT21), .B(G898), .Z(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(G902), .A3(G953), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT94), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n371), .A2(new_n413), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT86), .ZN(new_n421));
  AND2_X1   g235(.A1(KEYINPUT69), .A2(G119), .ZN(new_n422));
  NOR2_X1   g236(.A1(KEYINPUT69), .A2(G119), .ZN(new_n423));
  OAI21_X1  g237(.A(G116), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n375), .A2(G119), .ZN(new_n425));
  AND2_X1   g239(.A1(KEYINPUT85), .A2(KEYINPUT5), .ZN(new_n426));
  NOR2_X1   g240(.A1(KEYINPUT85), .A2(KEYINPUT5), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n424), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G113), .B1(new_n424), .B2(new_n428), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n421), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT2), .B(G113), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n424), .A3(new_n425), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n424), .A2(new_n425), .A3(new_n428), .ZN(new_n435));
  OR2_X1    g249(.A1(KEYINPUT69), .A2(G119), .ZN(new_n436));
  NAND2_X1  g250(.A1(KEYINPUT69), .A2(G119), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n375), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n435), .A2(new_n440), .A3(KEYINPUT86), .A4(G113), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n431), .A2(new_n434), .A3(new_n224), .A4(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n425), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n432), .B1(new_n438), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT70), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n434), .A3(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(KEYINPUT70), .B(new_n432), .C1(new_n438), .C2(new_n443), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n446), .A2(new_n199), .A3(new_n447), .A4(new_n212), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G110), .B(G122), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n442), .A2(new_n448), .A3(new_n450), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(KEYINPUT6), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n204), .A2(KEYINPUT0), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n208), .A2(new_n209), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G125), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n218), .A2(new_n318), .A3(new_n220), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G224), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(G953), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n460), .B(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT87), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n465));
  AND4_X1   g279(.A1(new_n464), .A2(new_n449), .A3(new_n465), .A4(new_n451), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n450), .B1(new_n442), .B2(new_n448), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n464), .B1(new_n467), .B2(new_n465), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n454), .B(new_n463), .C1(new_n466), .C2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(G210), .B1(G237), .B2(G902), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n450), .B(KEYINPUT8), .Z(new_n471));
  AND3_X1   g285(.A1(new_n424), .A2(KEYINPUT5), .A3(new_n425), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n434), .B1(new_n472), .B2(new_n430), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n471), .B1(new_n473), .B2(new_n224), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n431), .A2(new_n434), .A3(new_n441), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n474), .B1(new_n475), .B2(new_n224), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n477), .A2(KEYINPUT88), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n458), .A2(new_n459), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n477), .B2(new_n462), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n462), .A2(new_n477), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n458), .A2(new_n459), .A3(new_n478), .A4(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n476), .A2(new_n480), .A3(new_n453), .A4(new_n482), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n483), .A2(new_n188), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n469), .A2(new_n470), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n470), .B1(new_n469), .B2(new_n484), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(G214), .B1(G237), .B2(G902), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n420), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n446), .A2(new_n447), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n248), .A2(new_n384), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n493), .B(G131), .C1(new_n384), .C2(new_n251), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n257), .A2(new_n221), .A3(new_n494), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n258), .A2(new_n210), .B1(new_n495), .B2(KEYINPUT68), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT68), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n257), .A2(new_n221), .A3(new_n497), .A4(new_n494), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n492), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n257), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n246), .A2(KEYINPUT66), .B1(new_n242), .B2(new_n252), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n256), .B1(new_n501), .B2(new_n250), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n210), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n495), .A3(new_n492), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(KEYINPUT71), .B(KEYINPUT28), .C1(new_n499), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n309), .A2(G210), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(new_n197), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n508), .B(new_n509), .Z(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT28), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n495), .A2(KEYINPUT68), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n503), .A2(new_n513), .A3(new_n498), .ZN(new_n514));
  INV_X1    g328(.A(new_n492), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n512), .B1(new_n516), .B2(new_n504), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n504), .A2(new_n512), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT71), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n506), .B(new_n511), .C1(new_n517), .C2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n457), .B1(new_n255), .B2(new_n257), .ZN(new_n524));
  INV_X1    g338(.A(new_n495), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT30), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n515), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n510), .A3(new_n504), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT31), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT31), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n528), .A2(new_n531), .A3(new_n510), .A4(new_n504), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n521), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(G472), .A2(G902), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n533), .A2(KEYINPUT32), .A3(new_n534), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT74), .B1(new_n526), .B2(new_n492), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT74), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n541), .B(new_n515), .C1(new_n524), .C2(new_n525), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n504), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT28), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n544), .A2(KEYINPUT29), .A3(new_n510), .A4(new_n518), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n188), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT73), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n528), .A2(new_n504), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n547), .B1(new_n548), .B2(new_n511), .ZN(new_n549));
  AOI211_X1 g363(.A(KEYINPUT73), .B(new_n510), .C1(new_n528), .C2(new_n504), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n506), .B1(new_n517), .B2(new_n520), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT29), .B1(new_n552), .B2(new_n510), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n546), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G472), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n538), .B(new_n539), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT22), .B(G137), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n557), .B(new_n558), .Z(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n339), .A2(new_n342), .ZN(new_n561));
  OAI21_X1  g375(.A(G119), .B1(new_n381), .B2(new_n382), .ZN(new_n562));
  OAI21_X1  g376(.A(G128), .B1(new_n422), .B2(new_n423), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT23), .ZN(new_n564));
  NOR2_X1   g378(.A1(KEYINPUT23), .A2(G128), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n436), .A2(new_n437), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n566), .A3(G110), .ZN(new_n567));
  XOR2_X1   g381(.A(KEYINPUT24), .B(G110), .Z(new_n568));
  AND3_X1   g382(.A1(new_n568), .A2(new_n562), .A3(new_n563), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AND4_X1   g384(.A1(KEYINPUT76), .A2(new_n561), .A3(new_n567), .A4(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n569), .B1(new_n339), .B2(new_n342), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT76), .B1(new_n572), .B2(new_n567), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n342), .A2(new_n327), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n562), .A2(new_n563), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(new_n568), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n564), .A2(new_n566), .ZN(new_n578));
  INV_X1    g392(.A(G110), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT77), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(G110), .B1(new_n564), .B2(new_n566), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT77), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n575), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n560), .B1(new_n574), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n572), .A2(new_n567), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT76), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n572), .A2(KEYINPUT76), .A3(new_n567), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n584), .ZN(new_n592));
  OAI22_X1  g406(.A1(new_n583), .A2(KEYINPUT77), .B1(new_n576), .B2(new_n568), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n342), .B(new_n327), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n594), .A3(new_n559), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n586), .A2(new_n595), .A3(new_n188), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT25), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n586), .A2(new_n595), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n396), .B1(G234), .B2(new_n188), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT78), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n600), .A2(KEYINPUT78), .A3(new_n601), .ZN(new_n605));
  INV_X1    g419(.A(new_n601), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n188), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT79), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n586), .A2(new_n595), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n308), .A2(new_n491), .A3(new_n556), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  AND2_X1   g427(.A1(new_n533), .A2(new_n188), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n535), .B1(new_n614), .B2(new_n555), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n610), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n308), .ZN(new_n617));
  INV_X1    g431(.A(new_n419), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n469), .A2(new_n484), .ZN(new_n619));
  INV_X1    g433(.A(new_n470), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT95), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n485), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n469), .A2(KEYINPUT95), .A3(new_n470), .A4(new_n484), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n624), .A2(new_n489), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n617), .A2(new_n618), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT33), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n398), .A2(new_n399), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT96), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT96), .B1(new_n403), .B2(new_n628), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n631), .B1(new_n632), .B2(new_n629), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n188), .A2(G478), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT97), .B(G478), .Z(new_n635));
  OAI22_X1  g449(.A1(new_n633), .A2(new_n634), .B1(new_n408), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n366), .A2(new_n370), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n627), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT98), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT34), .B(G104), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  INV_X1    g457(.A(new_n413), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n365), .A2(new_n360), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n645), .A2(new_n370), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n627), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT35), .B(G107), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  AND2_X1   g465(.A1(new_n533), .A2(new_n534), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n555), .B1(new_n533), .B2(new_n188), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI22_X1  g468(.A1(new_n574), .A2(new_n585), .B1(KEYINPUT36), .B2(new_n560), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n560), .A2(KEYINPUT36), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n591), .A2(new_n594), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n655), .A2(new_n608), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT99), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n604), .A2(new_n605), .A3(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n308), .A2(new_n491), .A3(new_n654), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT37), .B(G110), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT100), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n661), .B(new_n663), .ZN(G12));
  XOR2_X1   g478(.A(new_n415), .B(KEYINPUT102), .Z(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT101), .B(G900), .Z(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(new_n417), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n647), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(KEYINPUT78), .B1(new_n600), .B2(new_n601), .ZN(new_n672));
  AOI211_X1 g486(.A(new_n603), .B(new_n606), .C1(new_n598), .C2(new_n599), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n626), .B1(new_n674), .B2(new_n659), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n308), .A2(new_n556), .A3(new_n671), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  XNOR2_X1  g491(.A(new_n669), .B(KEYINPUT39), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n308), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n681));
  INV_X1    g495(.A(new_n548), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n511), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n188), .B1(new_n543), .B2(new_n510), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n538), .A2(new_n539), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n488), .B(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n371), .A2(new_n413), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n489), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n687), .A2(new_n689), .A3(new_n691), .A4(new_n660), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n680), .A2(new_n681), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G143), .ZN(G45));
  NOR2_X1   g508(.A1(new_n638), .A2(new_n670), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n308), .A2(new_n556), .A3(new_n675), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  OAI21_X1  g511(.A(new_n188), .B1(new_n282), .B2(new_n288), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G469), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n303), .A3(new_n289), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n626), .A2(new_n700), .A3(new_n618), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n701), .A2(new_n556), .A3(new_n611), .A4(new_n639), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT41), .B(G113), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  NAND4_X1  g518(.A1(new_n701), .A2(new_n556), .A3(new_n611), .A4(new_n648), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  NOR2_X1   g520(.A1(new_n420), .A2(new_n700), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n556), .A2(new_n675), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  XNOR2_X1  g523(.A(new_n534), .B(KEYINPUT104), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n542), .A2(new_n504), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n512), .B1(new_n711), .B2(new_n540), .ZN(new_n712));
  INV_X1    g526(.A(new_n518), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT105), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n544), .A2(new_n715), .A3(new_n518), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n716), .A3(new_n511), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n530), .A2(new_n532), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n710), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n653), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n701), .A2(new_n611), .A3(new_n690), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NOR2_X1   g536(.A1(new_n626), .A2(new_n700), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n720), .A3(new_n695), .A4(new_n660), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  NAND2_X1  g539(.A1(new_n298), .A2(KEYINPUT106), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n486), .A2(new_n490), .A3(new_n487), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n289), .A2(new_n295), .A3(new_n728), .A4(new_n297), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n726), .A2(new_n303), .A3(new_n727), .A4(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n611), .A3(new_n556), .A4(new_n695), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n652), .A2(KEYINPUT32), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n735), .B(new_n539), .C1(new_n555), .C2(new_n554), .ZN(new_n736));
  INV_X1    g550(.A(new_n695), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n733), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n736), .A2(new_n738), .A3(new_n611), .A4(new_n731), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G131), .ZN(G33));
  NAND2_X1  g555(.A1(new_n556), .A2(new_n611), .ZN(new_n742));
  INV_X1    g556(.A(new_n671), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n742), .A2(new_n743), .A3(new_n730), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT107), .B(G134), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G36));
  AND2_X1   g560(.A1(new_n293), .A2(new_n294), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(KEYINPUT45), .ZN(new_n748));
  OAI21_X1  g562(.A(G469), .B1(new_n747), .B2(KEYINPUT45), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n296), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT46), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n289), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n751), .A2(KEYINPUT46), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n303), .B(new_n678), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n371), .A2(new_n636), .ZN(new_n757));
  XOR2_X1   g571(.A(new_n757), .B(KEYINPUT43), .Z(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n615), .A3(new_n660), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n727), .B(KEYINPUT108), .Z(new_n763));
  NAND4_X1  g577(.A1(new_n756), .A2(new_n761), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  OAI21_X1  g579(.A(new_n303), .B1(new_n753), .B2(new_n754), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(KEYINPUT47), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(KEYINPUT47), .ZN(new_n768));
  INV_X1    g582(.A(new_n727), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n737), .A2(new_n556), .A3(new_n611), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  NOR4_X1   g586(.A1(new_n610), .A2(new_n757), .A3(new_n302), .A4(new_n490), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n699), .A2(new_n289), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT49), .Z(new_n775));
  NAND4_X1  g589(.A1(new_n773), .A2(new_n775), .A3(new_n687), .A4(new_n689), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n645), .A2(new_n370), .A3(new_n669), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n413), .A2(KEYINPUT109), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n407), .B(new_n779), .C1(new_n412), .C2(new_n411), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n777), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(new_n660), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(new_n308), .A3(new_n556), .A4(new_n727), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n720), .A2(new_n660), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n695), .ZN(new_n785));
  OAI211_X1 g599(.A(KEYINPUT53), .B(new_n783), .C1(new_n785), .C2(new_n730), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n778), .A2(new_n371), .A3(new_n780), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n638), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n489), .B(new_n419), .C1(new_n486), .C2(new_n487), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n612), .B(new_n661), .C1(new_n617), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n786), .A2(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n721), .A2(new_n708), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n794), .A2(KEYINPUT113), .A3(new_n702), .A4(new_n705), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n744), .B1(new_n734), .B2(new_n739), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n702), .A2(new_n705), .A3(new_n721), .A4(new_n708), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n793), .A2(new_n795), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n676), .A2(new_n724), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n726), .A2(new_n303), .A3(new_n729), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n626), .A2(new_n371), .A3(new_n413), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n604), .A2(new_n605), .A3(new_n659), .A4(new_n669), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n686), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n801), .A2(new_n802), .A3(new_n696), .A4(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n676), .A2(new_n696), .A3(new_n806), .A4(new_n724), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT52), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n800), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n792), .A2(new_n797), .ZN(new_n812));
  INV_X1    g626(.A(new_n785), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n782), .A2(new_n556), .A3(new_n727), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n813), .A2(new_n731), .B1(new_n814), .B2(new_n308), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n812), .A2(new_n796), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n807), .A2(new_n817), .A3(new_n809), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n817), .B1(new_n807), .B2(new_n809), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  AOI211_X1 g635(.A(KEYINPUT54), .B(new_n811), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(KEYINPUT53), .B(new_n816), .C1(new_n818), .C2(new_n819), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n809), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n808), .A2(KEYINPUT52), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT111), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n807), .A2(new_n817), .A3(new_n809), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(KEYINPUT112), .A3(KEYINPUT53), .A4(new_n816), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT110), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n812), .A2(new_n796), .A3(new_n815), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n832), .B(new_n821), .C1(new_n833), .C2(new_n810), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n821), .B1(new_n833), .B2(new_n810), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT110), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n825), .A2(new_n831), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n822), .B1(new_n837), .B2(KEYINPUT54), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n758), .A2(new_n665), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n839), .A2(new_n611), .A3(new_n720), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n700), .A2(new_n489), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(new_n689), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT50), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n769), .A2(new_n700), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n839), .A2(new_n784), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n610), .A2(new_n415), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n687), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n847), .A2(new_n637), .A3(new_n636), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n843), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n840), .A2(new_n763), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n767), .A2(new_n768), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n699), .A2(new_n302), .A3(new_n289), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n842), .A2(KEYINPUT50), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n849), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n856), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n855), .B(new_n858), .Z(new_n859));
  NAND2_X1  g673(.A1(new_n262), .A2(G952), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n840), .B2(new_n723), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n861), .B1(new_n638), .B2(new_n847), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT115), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n736), .A2(new_n611), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n839), .A2(new_n844), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n864), .B(new_n865), .C1(new_n866), .C2(KEYINPUT48), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(KEYINPUT48), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n867), .B(new_n868), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n838), .A2(new_n859), .A3(new_n863), .A4(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(G952), .A2(G953), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n776), .B1(new_n870), .B2(new_n871), .ZN(G75));
  AOI21_X1  g686(.A(KEYINPUT53), .B1(new_n830), .B2(new_n816), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n811), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n188), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT56), .B1(new_n875), .B2(G210), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n454), .B1(new_n466), .B2(new_n468), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(new_n463), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT55), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n876), .A2(new_n879), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n262), .A2(G952), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(G51));
  XOR2_X1   g697(.A(new_n874), .B(KEYINPUT54), .Z(new_n884));
  XNOR2_X1  g698(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(new_n296), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n288), .B2(new_n282), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n875), .A2(new_n750), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n882), .B1(new_n888), .B2(new_n889), .ZN(G54));
  INV_X1    g704(.A(new_n882), .ZN(new_n891));
  NAND2_X1  g705(.A1(KEYINPUT58), .A2(G475), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT118), .Z(new_n893));
  AND2_X1   g707(.A1(new_n875), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n891), .B1(new_n894), .B2(new_n357), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n357), .B2(new_n894), .ZN(G60));
  XNOR2_X1  g710(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n897));
  NAND2_X1  g711(.A1(G478), .A2(G902), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n633), .B1(new_n838), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(KEYINPUT120), .B(new_n633), .C1(new_n838), .C2(new_n899), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n633), .A2(new_n899), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n882), .B1(new_n884), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n904), .A2(KEYINPUT121), .A3(new_n906), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(G63));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n912));
  NAND2_X1  g726(.A1(G217), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT60), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n912), .B1(new_n874), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n586), .A2(new_n595), .ZN(new_n916));
  INV_X1    g730(.A(new_n914), .ZN(new_n917));
  OAI211_X1 g731(.A(KEYINPUT122), .B(new_n917), .C1(new_n873), .C2(new_n811), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n919), .A2(new_n891), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n655), .A2(new_n657), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n915), .B2(new_n918), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n922), .A2(KEYINPUT123), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(KEYINPUT123), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g741(.A(KEYINPUT61), .B(new_n920), .C1(new_n923), .C2(new_n924), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(G66));
  INV_X1    g743(.A(new_n416), .ZN(new_n930));
  OAI21_X1  g744(.A(G953), .B1(new_n930), .B2(new_n461), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n812), .B2(G953), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT124), .Z(new_n933));
  OAI21_X1  g747(.A(new_n877), .B1(G898), .B2(new_n262), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G69));
  AOI21_X1  g749(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n771), .A2(new_n764), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n788), .A2(new_n727), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n679), .A2(new_n742), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n801), .A2(new_n696), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n693), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT62), .Z(new_n944));
  NAND2_X1  g758(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n941), .A2(new_n944), .A3(KEYINPUT125), .ZN(new_n948));
  AOI21_X1  g762(.A(G953), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n523), .A2(new_n527), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n349), .A2(new_n351), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n950), .B(new_n951), .Z(new_n952));
  OR2_X1    g766(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n954));
  NAND2_X1  g768(.A1(G900), .A2(G953), .ZN(new_n955));
  INV_X1    g769(.A(new_n942), .ZN(new_n956));
  INV_X1    g770(.A(new_n804), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n755), .A2(new_n864), .A3(new_n957), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n938), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n796), .A2(KEYINPUT126), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n796), .A2(KEYINPUT126), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n952), .B(new_n955), .C1(new_n962), .C2(G953), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n953), .A2(new_n954), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n954), .B1(new_n953), .B2(new_n963), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n937), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n953), .A2(new_n963), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n953), .A2(new_n954), .A3(new_n963), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n936), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n966), .A2(new_n970), .ZN(G72));
  NAND3_X1  g785(.A1(new_n947), .A2(new_n812), .A3(new_n948), .ZN(new_n972));
  NAND2_X1  g786(.A1(G472), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT63), .Z(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n683), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n551), .A2(new_n529), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n837), .A2(new_n974), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n812), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n974), .B1(new_n962), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n980), .A2(new_n511), .A3(new_n682), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n891), .A2(new_n976), .A3(new_n978), .A4(new_n981), .ZN(G57));
endmodule


