

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U551 ( .A1(n686), .A2(n799), .ZN(n735) );
  NOR2_X1 U552 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  AND2_X1 U553 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U554 ( .A1(G651), .A2(n629), .ZN(n640) );
  AND2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n887) );
  NAND2_X1 U556 ( .A1(G113), .A2(n887), .ZN(n518) );
  INV_X1 U557 ( .A(G2105), .ZN(n521) );
  NOR2_X1 U558 ( .A1(G2104), .A2(n521), .ZN(n888) );
  NAND2_X1 U559 ( .A1(G125), .A2(n888), .ZN(n517) );
  AND2_X1 U560 ( .A1(n518), .A2(n517), .ZN(n682) );
  XOR2_X2 U561 ( .A(KEYINPUT17), .B(n519), .Z(n884) );
  NAND2_X1 U562 ( .A1(G137), .A2(n884), .ZN(n520) );
  XNOR2_X1 U563 ( .A(n520), .B(KEYINPUT64), .ZN(n524) );
  AND2_X1 U564 ( .A1(n521), .A2(G2104), .ZN(n883) );
  NAND2_X1 U565 ( .A1(G101), .A2(n883), .ZN(n522) );
  XOR2_X1 U566 ( .A(KEYINPUT23), .B(n522), .Z(n523) );
  AND2_X1 U567 ( .A1(n524), .A2(n523), .ZN(n684) );
  AND2_X1 U568 ( .A1(n682), .A2(n684), .ZN(G160) );
  NOR2_X1 U569 ( .A1(G651), .A2(G543), .ZN(n636) );
  NAND2_X1 U570 ( .A1(G85), .A2(n636), .ZN(n526) );
  XOR2_X1 U571 ( .A(KEYINPUT0), .B(G543), .Z(n629) );
  INV_X1 U572 ( .A(G651), .ZN(n527) );
  NOR2_X1 U573 ( .A1(n629), .A2(n527), .ZN(n637) );
  NAND2_X1 U574 ( .A1(G72), .A2(n637), .ZN(n525) );
  NAND2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n532) );
  NOR2_X1 U576 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n528), .Z(n642) );
  NAND2_X1 U578 ( .A1(G60), .A2(n642), .ZN(n530) );
  NAND2_X1 U579 ( .A1(G47), .A2(n640), .ZN(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n531) );
  OR2_X1 U581 ( .A1(n532), .A2(n531), .ZN(G290) );
  XOR2_X1 U582 ( .A(G2446), .B(G2430), .Z(n534) );
  XNOR2_X1 U583 ( .A(G2451), .B(G2454), .ZN(n533) );
  XNOR2_X1 U584 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U585 ( .A(n535), .B(G2427), .Z(n537) );
  XNOR2_X1 U586 ( .A(G1341), .B(G1348), .ZN(n536) );
  XNOR2_X1 U587 ( .A(n537), .B(n536), .ZN(n541) );
  XOR2_X1 U588 ( .A(G2443), .B(KEYINPUT104), .Z(n539) );
  XNOR2_X1 U589 ( .A(G2438), .B(G2435), .ZN(n538) );
  XNOR2_X1 U590 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U591 ( .A(n541), .B(n540), .Z(n542) );
  AND2_X1 U592 ( .A1(G14), .A2(n542), .ZN(G401) );
  AND2_X1 U593 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U594 ( .A(G132), .ZN(G219) );
  INV_X1 U595 ( .A(G82), .ZN(G220) );
  NAND2_X1 U596 ( .A1(G90), .A2(n636), .ZN(n544) );
  NAND2_X1 U597 ( .A1(G77), .A2(n637), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U599 ( .A(KEYINPUT9), .B(n545), .ZN(n549) );
  NAND2_X1 U600 ( .A1(G64), .A2(n642), .ZN(n547) );
  NAND2_X1 U601 ( .A1(G52), .A2(n640), .ZN(n546) );
  AND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U603 ( .A1(n549), .A2(n548), .ZN(G301) );
  INV_X1 U604 ( .A(G301), .ZN(G171) );
  NAND2_X1 U605 ( .A1(n636), .A2(G89), .ZN(n550) );
  XOR2_X1 U606 ( .A(KEYINPUT4), .B(n550), .Z(n553) );
  NAND2_X1 U607 ( .A1(n637), .A2(G76), .ZN(n551) );
  XOR2_X1 U608 ( .A(KEYINPUT70), .B(n551), .Z(n552) );
  NOR2_X1 U609 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U610 ( .A(KEYINPUT5), .B(n554), .ZN(n555) );
  XNOR2_X1 U611 ( .A(n555), .B(KEYINPUT71), .ZN(n560) );
  NAND2_X1 U612 ( .A1(G63), .A2(n642), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G51), .A2(n640), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U615 ( .A(KEYINPUT6), .B(n558), .Z(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U617 ( .A(KEYINPUT7), .B(n561), .ZN(G168) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U620 ( .A(n562), .B(KEYINPUT66), .ZN(n563) );
  XNOR2_X1 U621 ( .A(KEYINPUT10), .B(n563), .ZN(G223) );
  INV_X1 U622 ( .A(G223), .ZN(n831) );
  NAND2_X1 U623 ( .A1(n831), .A2(G567), .ZN(n564) );
  XOR2_X1 U624 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  NAND2_X1 U625 ( .A1(n636), .A2(G81), .ZN(n565) );
  XNOR2_X1 U626 ( .A(n565), .B(KEYINPUT12), .ZN(n567) );
  NAND2_X1 U627 ( .A1(G68), .A2(n637), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT13), .B(n568), .Z(n572) );
  NAND2_X1 U630 ( .A1(G56), .A2(n642), .ZN(n569) );
  XNOR2_X1 U631 ( .A(n569), .B(KEYINPUT67), .ZN(n570) );
  XNOR2_X1 U632 ( .A(n570), .B(KEYINPUT14), .ZN(n571) );
  NOR2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U634 ( .A(n573), .B(KEYINPUT68), .ZN(n575) );
  NAND2_X1 U635 ( .A1(G43), .A2(n640), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n575), .A2(n574), .ZN(n976) );
  INV_X1 U637 ( .A(G860), .ZN(n840) );
  OR2_X1 U638 ( .A1(n976), .A2(n840), .ZN(G153) );
  NAND2_X1 U639 ( .A1(G92), .A2(n636), .ZN(n577) );
  NAND2_X1 U640 ( .A1(G79), .A2(n637), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G66), .A2(n642), .ZN(n579) );
  NAND2_X1 U643 ( .A1(G54), .A2(n640), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT15), .B(n582), .Z(n977) );
  NOR2_X1 U647 ( .A1(n977), .A2(G868), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(KEYINPUT69), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G868), .A2(G301), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U651 ( .A1(G65), .A2(n642), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G53), .A2(n640), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U654 ( .A1(G91), .A2(n636), .ZN(n589) );
  NAND2_X1 U655 ( .A1(G78), .A2(n637), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n713) );
  INV_X1 U658 ( .A(n713), .ZN(G299) );
  NOR2_X1 U659 ( .A1(G868), .A2(G299), .ZN(n592) );
  XOR2_X1 U660 ( .A(KEYINPUT73), .B(n592), .Z(n595) );
  INV_X1 U661 ( .A(G868), .ZN(n658) );
  NOR2_X1 U662 ( .A1(G286), .A2(n658), .ZN(n593) );
  XNOR2_X1 U663 ( .A(KEYINPUT72), .B(n593), .ZN(n594) );
  NOR2_X1 U664 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U665 ( .A1(n840), .A2(G559), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n596), .A2(n977), .ZN(n597) );
  XNOR2_X1 U667 ( .A(n597), .B(KEYINPUT74), .ZN(n598) );
  XNOR2_X1 U668 ( .A(KEYINPUT16), .B(n598), .ZN(G148) );
  NOR2_X1 U669 ( .A1(G868), .A2(n976), .ZN(n601) );
  NAND2_X1 U670 ( .A1(G868), .A2(n977), .ZN(n599) );
  NOR2_X1 U671 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U672 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U673 ( .A1(G99), .A2(n883), .ZN(n603) );
  NAND2_X1 U674 ( .A1(G111), .A2(n887), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n609) );
  NAND2_X1 U676 ( .A1(n888), .A2(G123), .ZN(n604) );
  XNOR2_X1 U677 ( .A(n604), .B(KEYINPUT18), .ZN(n606) );
  NAND2_X1 U678 ( .A1(G135), .A2(n884), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U680 ( .A(KEYINPUT75), .B(n607), .Z(n608) );
  NOR2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n934) );
  XNOR2_X1 U682 ( .A(n934), .B(G2096), .ZN(n611) );
  INV_X1 U683 ( .A(G2100), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n611), .A2(n610), .ZN(G156) );
  NAND2_X1 U685 ( .A1(G62), .A2(n642), .ZN(n613) );
  NAND2_X1 U686 ( .A1(G50), .A2(n640), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U688 ( .A(KEYINPUT81), .B(n614), .ZN(n620) );
  NAND2_X1 U689 ( .A1(G88), .A2(n636), .ZN(n615) );
  XOR2_X1 U690 ( .A(KEYINPUT82), .B(n615), .Z(n618) );
  NAND2_X1 U691 ( .A1(G75), .A2(n637), .ZN(n616) );
  XNOR2_X1 U692 ( .A(KEYINPUT83), .B(n616), .ZN(n617) );
  NOR2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n620), .A2(n619), .ZN(G303) );
  INV_X1 U695 ( .A(G303), .ZN(G166) );
  NAND2_X1 U696 ( .A1(G48), .A2(n640), .ZN(n627) );
  NAND2_X1 U697 ( .A1(G86), .A2(n636), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G61), .A2(n642), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n637), .A2(G73), .ZN(n623) );
  XOR2_X1 U701 ( .A(KEYINPUT2), .B(n623), .Z(n624) );
  NOR2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n628), .B(KEYINPUT80), .ZN(G305) );
  NAND2_X1 U705 ( .A1(G49), .A2(n640), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G87), .A2(n629), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U708 ( .A1(n642), .A2(n632), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G651), .A2(G74), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G559), .A2(n977), .ZN(n635) );
  XOR2_X1 U712 ( .A(n976), .B(n635), .Z(n839) );
  XNOR2_X1 U713 ( .A(G166), .B(G305), .ZN(n656) );
  NAND2_X1 U714 ( .A1(G93), .A2(n636), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G80), .A2(n637), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n640), .A2(G55), .ZN(n641) );
  XNOR2_X1 U718 ( .A(KEYINPUT77), .B(n641), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n642), .A2(G67), .ZN(n643) );
  XOR2_X1 U720 ( .A(KEYINPUT76), .B(n643), .Z(n644) );
  NOR2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U722 ( .A(KEYINPUT78), .B(n646), .Z(n647) );
  NOR2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U724 ( .A(KEYINPUT79), .B(n649), .ZN(n841) );
  XNOR2_X1 U725 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n651) );
  XNOR2_X1 U726 ( .A(G288), .B(KEYINPUT85), .ZN(n650) );
  XNOR2_X1 U727 ( .A(n651), .B(n650), .ZN(n652) );
  XOR2_X1 U728 ( .A(n841), .B(n652), .Z(n654) );
  XNOR2_X1 U729 ( .A(G290), .B(n713), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U731 ( .A(n656), .B(n655), .ZN(n908) );
  XNOR2_X1 U732 ( .A(n839), .B(n908), .ZN(n657) );
  NAND2_X1 U733 ( .A1(n657), .A2(G868), .ZN(n660) );
  NAND2_X1 U734 ( .A1(n658), .A2(n841), .ZN(n659) );
  NAND2_X1 U735 ( .A1(n660), .A2(n659), .ZN(G295) );
  NAND2_X1 U736 ( .A1(G2084), .A2(G2078), .ZN(n661) );
  XOR2_X1 U737 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XNOR2_X1 U739 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U740 ( .A1(n664), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U741 ( .A(KEYINPUT65), .B(G57), .ZN(G237) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U743 ( .A1(G108), .A2(G120), .ZN(n665) );
  NOR2_X1 U744 ( .A1(G237), .A2(n665), .ZN(n666) );
  NAND2_X1 U745 ( .A1(G69), .A2(n666), .ZN(n838) );
  NAND2_X1 U746 ( .A1(n838), .A2(G567), .ZN(n672) );
  NOR2_X1 U747 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U749 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U750 ( .A1(G96), .A2(n669), .ZN(n837) );
  NAND2_X1 U751 ( .A1(G2106), .A2(n837), .ZN(n670) );
  XNOR2_X1 U752 ( .A(KEYINPUT86), .B(n670), .ZN(n671) );
  NAND2_X1 U753 ( .A1(n672), .A2(n671), .ZN(n843) );
  NAND2_X1 U754 ( .A1(G483), .A2(G661), .ZN(n673) );
  NOR2_X1 U755 ( .A1(n843), .A2(n673), .ZN(n836) );
  NAND2_X1 U756 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U757 ( .A1(G102), .A2(n883), .ZN(n675) );
  NAND2_X1 U758 ( .A1(G138), .A2(n884), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n675), .A2(n674), .ZN(n679) );
  NAND2_X1 U760 ( .A1(G114), .A2(n887), .ZN(n677) );
  NAND2_X1 U761 ( .A1(G126), .A2(n888), .ZN(n676) );
  NAND2_X1 U762 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U763 ( .A1(n679), .A2(n678), .ZN(G164) );
  NOR2_X1 U764 ( .A1(G2090), .A2(G303), .ZN(n680) );
  XOR2_X1 U765 ( .A(KEYINPUT101), .B(n680), .Z(n681) );
  NAND2_X1 U766 ( .A1(G8), .A2(n681), .ZN(n751) );
  AND2_X1 U767 ( .A1(n682), .A2(G40), .ZN(n683) );
  NAND2_X1 U768 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U769 ( .A(KEYINPUT87), .B(n685), .Z(n798) );
  XNOR2_X1 U770 ( .A(KEYINPUT95), .B(n798), .ZN(n686) );
  NOR2_X1 U771 ( .A1(G164), .A2(G1384), .ZN(n799) );
  NOR2_X1 U772 ( .A1(G2084), .A2(n735), .ZN(n721) );
  NAND2_X1 U773 ( .A1(G8), .A2(n721), .ZN(n734) );
  NAND2_X1 U774 ( .A1(G8), .A2(n735), .ZN(n771) );
  NOR2_X1 U775 ( .A1(G1966), .A2(n771), .ZN(n732) );
  AND2_X1 U776 ( .A1(n735), .A2(G1961), .ZN(n688) );
  XNOR2_X1 U777 ( .A(G2078), .B(KEYINPUT25), .ZN(n951) );
  NOR2_X1 U778 ( .A1(n735), .A2(n951), .ZN(n687) );
  NOR2_X1 U779 ( .A1(n688), .A2(n687), .ZN(n725) );
  NAND2_X1 U780 ( .A1(n725), .A2(G171), .ZN(n720) );
  INV_X1 U781 ( .A(n735), .ZN(n694) );
  NAND2_X1 U782 ( .A1(n694), .A2(G2072), .ZN(n689) );
  XNOR2_X1 U783 ( .A(KEYINPUT27), .B(n689), .ZN(n692) );
  NAND2_X1 U784 ( .A1(G1956), .A2(n735), .ZN(n690) );
  XOR2_X1 U785 ( .A(KEYINPUT96), .B(n690), .Z(n691) );
  NOR2_X1 U786 ( .A1(n692), .A2(n691), .ZN(n712) );
  NOR2_X1 U787 ( .A1(n713), .A2(n712), .ZN(n693) );
  XOR2_X1 U788 ( .A(n693), .B(KEYINPUT28), .Z(n717) );
  NOR2_X1 U789 ( .A1(n694), .A2(G1348), .ZN(n696) );
  NOR2_X1 U790 ( .A1(G2067), .A2(n735), .ZN(n695) );
  NOR2_X1 U791 ( .A1(n696), .A2(n695), .ZN(n706) );
  INV_X1 U792 ( .A(G1996), .ZN(n949) );
  NOR2_X1 U793 ( .A1(n735), .A2(n949), .ZN(n698) );
  INV_X1 U794 ( .A(KEYINPUT26), .ZN(n697) );
  NAND2_X1 U795 ( .A1(n698), .A2(n697), .ZN(n701) );
  INV_X1 U796 ( .A(n698), .ZN(n699) );
  NAND2_X1 U797 ( .A1(n699), .A2(KEYINPUT26), .ZN(n700) );
  NAND2_X1 U798 ( .A1(n701), .A2(n700), .ZN(n704) );
  AND2_X1 U799 ( .A1(n735), .A2(G1341), .ZN(n702) );
  NOR2_X1 U800 ( .A1(n702), .A2(n976), .ZN(n703) );
  AND2_X1 U801 ( .A1(n704), .A2(n703), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n977), .A2(n709), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n706), .A2(n705), .ZN(n708) );
  INV_X1 U804 ( .A(KEYINPUT97), .ZN(n707) );
  XNOR2_X1 U805 ( .A(n708), .B(n707), .ZN(n711) );
  OR2_X1 U806 ( .A1(n977), .A2(n709), .ZN(n710) );
  NAND2_X1 U807 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U809 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U811 ( .A(n718), .B(KEYINPUT29), .Z(n719) );
  NAND2_X1 U812 ( .A1(n720), .A2(n719), .ZN(n743) );
  INV_X1 U813 ( .A(KEYINPUT98), .ZN(n729) );
  NOR2_X1 U814 ( .A1(n732), .A2(n721), .ZN(n722) );
  NAND2_X1 U815 ( .A1(G8), .A2(n722), .ZN(n723) );
  XNOR2_X1 U816 ( .A(n723), .B(KEYINPUT30), .ZN(n724) );
  NOR2_X1 U817 ( .A1(G168), .A2(n724), .ZN(n727) );
  NOR2_X1 U818 ( .A1(G171), .A2(n725), .ZN(n726) );
  NOR2_X1 U819 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U820 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U821 ( .A(n730), .B(KEYINPUT31), .ZN(n742) );
  AND2_X1 U822 ( .A1(n743), .A2(n742), .ZN(n731) );
  NOR2_X1 U823 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n753) );
  INV_X1 U825 ( .A(G8), .ZN(n741) );
  NOR2_X1 U826 ( .A1(G1971), .A2(n771), .ZN(n737) );
  NOR2_X1 U827 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U828 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U829 ( .A1(n738), .A2(G303), .ZN(n739) );
  XOR2_X1 U830 ( .A(KEYINPUT99), .B(n739), .Z(n740) );
  OR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n745) );
  AND2_X1 U832 ( .A1(n742), .A2(n745), .ZN(n744) );
  NAND2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n748) );
  INV_X1 U834 ( .A(n745), .ZN(n746) );
  OR2_X1 U835 ( .A1(n746), .A2(G286), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U837 ( .A(n749), .B(KEYINPUT32), .ZN(n760) );
  NAND2_X1 U838 ( .A1(n753), .A2(n760), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n752), .A2(n771), .ZN(n777) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n981) );
  AND2_X1 U842 ( .A1(n753), .A2(n981), .ZN(n758) );
  XOR2_X1 U843 ( .A(G1981), .B(G305), .Z(n973) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n754) );
  XOR2_X1 U845 ( .A(KEYINPUT100), .B(n754), .Z(n761) );
  NOR2_X1 U846 ( .A1(n771), .A2(n761), .ZN(n755) );
  NAND2_X1 U847 ( .A1(KEYINPUT33), .A2(n755), .ZN(n756) );
  NAND2_X1 U848 ( .A1(n973), .A2(n756), .ZN(n768) );
  INV_X1 U849 ( .A(n768), .ZN(n757) );
  AND2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n775) );
  INV_X1 U852 ( .A(KEYINPUT33), .ZN(n766) );
  INV_X1 U853 ( .A(n981), .ZN(n763) );
  NOR2_X1 U854 ( .A1(G1971), .A2(G303), .ZN(n979) );
  INV_X1 U855 ( .A(n761), .ZN(n987) );
  NOR2_X1 U856 ( .A1(n979), .A2(n987), .ZN(n762) );
  OR2_X1 U857 ( .A1(n763), .A2(n762), .ZN(n764) );
  OR2_X1 U858 ( .A1(n771), .A2(n764), .ZN(n765) );
  AND2_X1 U859 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n773) );
  NOR2_X1 U861 ( .A1(G1981), .A2(G305), .ZN(n769) );
  XOR2_X1 U862 ( .A(n769), .B(KEYINPUT24), .Z(n770) );
  NOR2_X1 U863 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n774) );
  AND2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U867 ( .A(n778), .B(KEYINPUT102), .ZN(n815) );
  NAND2_X1 U868 ( .A1(n883), .A2(G105), .ZN(n780) );
  XNOR2_X1 U869 ( .A(KEYINPUT38), .B(KEYINPUT92), .ZN(n779) );
  XNOR2_X1 U870 ( .A(n780), .B(n779), .ZN(n787) );
  NAND2_X1 U871 ( .A1(G141), .A2(n884), .ZN(n782) );
  NAND2_X1 U872 ( .A1(G129), .A2(n888), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G117), .A2(n887), .ZN(n783) );
  XNOR2_X1 U875 ( .A(KEYINPUT91), .B(n783), .ZN(n784) );
  NOR2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n896) );
  NAND2_X1 U878 ( .A1(G1996), .A2(n896), .ZN(n788) );
  XNOR2_X1 U879 ( .A(n788), .B(KEYINPUT93), .ZN(n797) );
  XOR2_X1 U880 ( .A(KEYINPUT90), .B(G1991), .Z(n957) );
  NAND2_X1 U881 ( .A1(n883), .A2(G95), .ZN(n791) );
  NAND2_X1 U882 ( .A1(G107), .A2(n887), .ZN(n789) );
  XOR2_X1 U883 ( .A(KEYINPUT89), .B(n789), .Z(n790) );
  NAND2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n795) );
  NAND2_X1 U885 ( .A1(G131), .A2(n884), .ZN(n793) );
  NAND2_X1 U886 ( .A1(G119), .A2(n888), .ZN(n792) );
  NAND2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n897) );
  NOR2_X1 U889 ( .A1(n957), .A2(n897), .ZN(n796) );
  NOR2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n928) );
  NOR2_X1 U891 ( .A1(n799), .A2(n798), .ZN(n826) );
  XOR2_X1 U892 ( .A(n826), .B(KEYINPUT94), .Z(n800) );
  NOR2_X1 U893 ( .A1(n928), .A2(n800), .ZN(n819) );
  NAND2_X1 U894 ( .A1(n884), .A2(G140), .ZN(n801) );
  XNOR2_X1 U895 ( .A(n801), .B(KEYINPUT88), .ZN(n803) );
  NAND2_X1 U896 ( .A1(G104), .A2(n883), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U898 ( .A(KEYINPUT34), .B(n804), .ZN(n809) );
  NAND2_X1 U899 ( .A1(G116), .A2(n887), .ZN(n806) );
  NAND2_X1 U900 ( .A1(G128), .A2(n888), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U902 ( .A(KEYINPUT35), .B(n807), .Z(n808) );
  NOR2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U904 ( .A(KEYINPUT36), .B(n810), .ZN(n904) );
  XNOR2_X1 U905 ( .A(G2067), .B(KEYINPUT37), .ZN(n824) );
  NOR2_X1 U906 ( .A1(n904), .A2(n824), .ZN(n930) );
  NAND2_X1 U907 ( .A1(n826), .A2(n930), .ZN(n822) );
  INV_X1 U908 ( .A(n822), .ZN(n811) );
  NOR2_X1 U909 ( .A1(n819), .A2(n811), .ZN(n813) );
  XNOR2_X1 U910 ( .A(G1986), .B(G290), .ZN(n986) );
  NAND2_X1 U911 ( .A1(n986), .A2(n826), .ZN(n812) );
  NAND2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n829) );
  NOR2_X1 U913 ( .A1(G1996), .A2(n896), .ZN(n925) );
  AND2_X1 U914 ( .A1(n957), .A2(n897), .ZN(n816) );
  XOR2_X1 U915 ( .A(KEYINPUT103), .B(n816), .Z(n929) );
  NOR2_X1 U916 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U917 ( .A1(n929), .A2(n817), .ZN(n818) );
  NOR2_X1 U918 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U919 ( .A1(n925), .A2(n820), .ZN(n821) );
  XNOR2_X1 U920 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U921 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n904), .A2(n824), .ZN(n937) );
  NAND2_X1 U923 ( .A1(n825), .A2(n937), .ZN(n827) );
  NAND2_X1 U924 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U926 ( .A(KEYINPUT40), .B(n830), .ZN(G329) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n831), .ZN(G217) );
  NAND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n833) );
  INV_X1 U929 ( .A(G661), .ZN(n832) );
  NOR2_X1 U930 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n834), .B(KEYINPUT105), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U933 ( .A1(n836), .A2(n835), .ZN(G188) );
  XOR2_X1 U934 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G108), .ZN(G238) );
  INV_X1 U938 ( .A(G69), .ZN(G235) );
  NOR2_X1 U939 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  NAND2_X1 U941 ( .A1(n840), .A2(n839), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(G145) );
  INV_X1 U943 ( .A(n843), .ZN(G319) );
  XOR2_X1 U944 ( .A(KEYINPUT110), .B(G2474), .Z(n845) );
  XNOR2_X1 U945 ( .A(KEYINPUT108), .B(KEYINPUT107), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U947 ( .A(n846), .B(KEYINPUT41), .Z(n848) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n856) );
  XOR2_X1 U950 ( .A(G1976), .B(G1971), .Z(n850) );
  XNOR2_X1 U951 ( .A(G1986), .B(G1956), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U953 ( .A(KEYINPUT109), .B(G1981), .Z(n852) );
  XNOR2_X1 U954 ( .A(G1966), .B(G1961), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U956 ( .A(n854), .B(n853), .Z(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(G229) );
  XOR2_X1 U958 ( .A(G2100), .B(G2096), .Z(n858) );
  XNOR2_X1 U959 ( .A(KEYINPUT42), .B(G2678), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U961 ( .A(KEYINPUT43), .B(G2090), .Z(n860) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2072), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U964 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U965 ( .A(G2084), .B(G2078), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n864), .B(n863), .ZN(G227) );
  NAND2_X1 U967 ( .A1(G124), .A2(n888), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n887), .A2(G112), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G100), .A2(n883), .ZN(n869) );
  NAND2_X1 U972 ( .A1(G136), .A2(n884), .ZN(n868) );
  NAND2_X1 U973 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U974 ( .A1(n871), .A2(n870), .ZN(G162) );
  XOR2_X1 U975 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n882) );
  NAND2_X1 U976 ( .A1(G118), .A2(n887), .ZN(n873) );
  NAND2_X1 U977 ( .A1(G130), .A2(n888), .ZN(n872) );
  NAND2_X1 U978 ( .A1(n873), .A2(n872), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G106), .A2(n883), .ZN(n875) );
  NAND2_X1 U980 ( .A1(G142), .A2(n884), .ZN(n874) );
  NAND2_X1 U981 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U982 ( .A(KEYINPUT111), .B(n876), .ZN(n877) );
  XNOR2_X1 U983 ( .A(KEYINPUT45), .B(n877), .ZN(n878) );
  NOR2_X1 U984 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U985 ( .A(G164), .B(n880), .ZN(n881) );
  XNOR2_X1 U986 ( .A(n882), .B(n881), .ZN(n903) );
  NAND2_X1 U987 ( .A1(G103), .A2(n883), .ZN(n886) );
  NAND2_X1 U988 ( .A1(G139), .A2(n884), .ZN(n885) );
  NAND2_X1 U989 ( .A1(n886), .A2(n885), .ZN(n895) );
  XNOR2_X1 U990 ( .A(KEYINPUT114), .B(KEYINPUT47), .ZN(n893) );
  NAND2_X1 U991 ( .A1(n887), .A2(G115), .ZN(n891) );
  NAND2_X1 U992 ( .A1(n888), .A2(G127), .ZN(n889) );
  XOR2_X1 U993 ( .A(KEYINPUT113), .B(n889), .Z(n890) );
  NAND2_X1 U994 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U995 ( .A(n893), .B(n892), .Z(n894) );
  NOR2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n919) );
  XNOR2_X1 U997 ( .A(n919), .B(n896), .ZN(n898) );
  XOR2_X1 U998 ( .A(n898), .B(n897), .Z(n899) );
  XOR2_X1 U999 ( .A(n899), .B(G162), .Z(n901) );
  XNOR2_X1 U1000 ( .A(G160), .B(n934), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n904), .B(KEYINPUT48), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n907), .ZN(G395) );
  XOR2_X1 U1006 ( .A(n908), .B(G286), .Z(n910) );
  XNOR2_X1 U1007 ( .A(G171), .B(n977), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1009 ( .A(n911), .B(n976), .Z(n912) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n912), .ZN(G397) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n913) );
  XOR2_X1 U1012 ( .A(KEYINPUT49), .B(n913), .Z(n914) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n914), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n915), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n916) );
  XOR2_X1 U1016 ( .A(KEYINPUT115), .B(n916), .Z(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(KEYINPUT55), .ZN(n968) );
  XNOR2_X1 U1020 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n944) );
  XOR2_X1 U1021 ( .A(G2072), .B(n919), .Z(n921) );
  XOR2_X1 U1022 ( .A(G164), .B(G2078), .Z(n920) );
  NOR2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1024 ( .A(KEYINPUT50), .B(n922), .ZN(n941) );
  XNOR2_X1 U1025 ( .A(G2090), .B(G162), .ZN(n923) );
  XNOR2_X1 U1026 ( .A(n923), .B(KEYINPUT117), .ZN(n924) );
  NOR2_X1 U1027 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1028 ( .A(KEYINPUT51), .B(n926), .Z(n927) );
  NAND2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n939) );
  XNOR2_X1 U1030 ( .A(G160), .B(G2084), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(n935), .B(KEYINPUT116), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(n942), .B(KEYINPUT52), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(n944), .B(n943), .ZN(n945) );
  NAND2_X1 U1040 ( .A1(n968), .A2(n945), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n946), .A2(G29), .ZN(n1029) );
  XNOR2_X1 U1042 ( .A(G2090), .B(G35), .ZN(n963) );
  XNOR2_X1 U1043 ( .A(G2067), .B(G26), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(G33), .B(G2072), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n956) );
  XNOR2_X1 U1046 ( .A(G32), .B(n949), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n950), .A2(G28), .ZN(n954) );
  XOR2_X1 U1048 ( .A(G27), .B(n951), .Z(n952) );
  XNOR2_X1 U1049 ( .A(KEYINPUT120), .B(n952), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1052 ( .A(G25), .B(n957), .Z(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1054 ( .A(KEYINPUT53), .B(n960), .Z(n961) );
  XNOR2_X1 U1055 ( .A(n961), .B(KEYINPUT121), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1057 ( .A(G2084), .B(G34), .Z(n964) );
  XNOR2_X1 U1058 ( .A(KEYINPUT54), .B(n964), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(n968), .B(n967), .ZN(n970) );
  INV_X1 U1061 ( .A(G29), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n971), .ZN(n1027) );
  INV_X1 U1064 ( .A(G16), .ZN(n1023) );
  XOR2_X1 U1065 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n972) );
  XNOR2_X1 U1066 ( .A(n1023), .B(n972), .ZN(n998) );
  XNOR2_X1 U1067 ( .A(G1966), .B(G168), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(n975), .B(KEYINPUT57), .ZN(n996) );
  XNOR2_X1 U1070 ( .A(n976), .B(G1341), .ZN(n994) );
  XOR2_X1 U1071 ( .A(G1348), .B(n977), .Z(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n985) );
  NAND2_X1 U1073 ( .A1(G1971), .A2(G303), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(G1956), .B(G299), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n991) );
  XNOR2_X1 U1078 ( .A(G171), .B(G1961), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(KEYINPUT123), .B(n992), .ZN(n993) );
  NOR2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n1025) );
  XOR2_X1 U1086 ( .A(G4), .B(KEYINPUT126), .Z(n1000) );
  XNOR2_X1 U1087 ( .A(G1348), .B(KEYINPUT59), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(n1000), .B(n999), .ZN(n1008) );
  XNOR2_X1 U1089 ( .A(G1341), .B(G19), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(G1981), .B(G6), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(KEYINPUT124), .B(n1003), .Z(n1005) );
  XNOR2_X1 U1093 ( .A(G1956), .B(G20), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(n1006), .B(KEYINPUT125), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1009), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(G1966), .B(G21), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(G5), .B(G1961), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1020) );
  XNOR2_X1 U1102 ( .A(G1971), .B(G22), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(G23), .B(G1976), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XOR2_X1 U1105 ( .A(G1986), .B(G24), .Z(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(KEYINPUT58), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1109 ( .A(KEYINPUT61), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

