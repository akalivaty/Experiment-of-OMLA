//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G226), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  OAI22_X1  g0008(.A1(new_n202), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n209), .B(new_n215), .C1(G116), .C2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G1), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT64), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n223), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n230), .A2(new_n221), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(new_n224), .B2(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n226), .A2(new_n229), .A3(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G264), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G226), .B(G232), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n238), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G107), .ZN(new_n247));
  INV_X1    g0047(.A(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n207), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G200), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G77), .ZN(new_n258));
  OAI211_X1 g0058(.A(G223), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  OAI211_X1 g0060(.A(G222), .B(new_n260), .C1(new_n255), .C2(new_n256), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT69), .ZN(new_n263));
  AND2_X1   g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n231), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT69), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n258), .A2(new_n266), .A3(new_n259), .A4(new_n261), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n263), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  AOI21_X1  g0070(.A(G1), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT68), .B1(new_n264), .B2(new_n231), .ZN(new_n272));
  AND2_X1   g0072(.A1(G1), .A2(G13), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT68), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n271), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n278), .B1(new_n272), .B2(new_n276), .ZN(new_n279));
  AOI22_X1  g0079(.A1(G226), .A2(new_n277), .B1(new_n279), .B2(new_n271), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n254), .B1(new_n268), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT76), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n281), .B(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(KEYINPUT10), .B1(new_n283), .B2(KEYINPUT77), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G150), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT70), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n287), .B1(new_n288), .B2(G20), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n221), .A2(KEYINPUT70), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT8), .B(G58), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n286), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT71), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n203), .A2(G20), .ZN(new_n296));
  OAI211_X1 g0096(.A(KEYINPUT71), .B(new_n286), .C1(new_n291), .C2(new_n292), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n273), .B1(new_n222), .B2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n220), .A2(G13), .A3(G20), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n202), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n299), .B1(G1), .B2(new_n221), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G50), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n301), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n268), .A2(G190), .A3(new_n280), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n301), .A2(KEYINPUT9), .A3(new_n304), .A4(new_n307), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n284), .B(new_n314), .C1(KEYINPUT77), .C2(new_n283), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT78), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n316), .B(KEYINPUT10), .C1(new_n313), .C2(new_n283), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n268), .A2(new_n280), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n282), .B1(new_n319), .B2(G200), .ZN(new_n320));
  AOI211_X1 g0120(.A(KEYINPUT76), .B(new_n254), .C1(new_n268), .C2(new_n280), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n322), .A2(new_n311), .A3(new_n310), .A4(new_n312), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n316), .B1(new_n323), .B2(KEYINPUT10), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n315), .B1(new_n318), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n279), .A2(new_n271), .ZN(new_n326));
  INV_X1    g0126(.A(new_n277), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(new_n208), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT72), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT73), .B(G107), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n257), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT3), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n288), .ZN(new_n333));
  NAND2_X1  g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n260), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(G1698), .ZN(new_n337));
  OAI221_X1 g0137(.A(new_n331), .B1(new_n336), .B2(new_n218), .C1(new_n212), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n265), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n328), .A2(KEYINPUT72), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n329), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n341), .A2(G179), .ZN(new_n342));
  INV_X1    g0142(.A(G169), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G20), .A2(G77), .ZN(new_n345));
  INV_X1    g0145(.A(new_n285), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT15), .B(G87), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n345), .B1(new_n292), .B2(new_n346), .C1(new_n291), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n300), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT74), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n303), .A2(new_n207), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n306), .A2(G77), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n342), .A2(new_n344), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n308), .B1(G179), .B2(new_n319), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n355), .B1(new_n343), .B2(new_n319), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G190), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n341), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT75), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n353), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n350), .A2(KEYINPUT75), .A3(new_n351), .A4(new_n352), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n341), .A2(G200), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n359), .A2(new_n361), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n325), .A2(new_n354), .A3(new_n357), .A4(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT79), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT10), .B1(new_n313), .B2(new_n283), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT78), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n317), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n356), .B1(new_n370), .B2(new_n315), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n371), .A2(KEYINPUT79), .A3(new_n354), .A4(new_n364), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT13), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G97), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n374), .B1(new_n336), .B2(new_n206), .C1(new_n218), .C2(new_n337), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(new_n265), .B1(new_n271), .B2(new_n279), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n277), .A2(G238), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n373), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(new_n373), .A3(new_n377), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(G190), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n375), .A2(new_n265), .ZN(new_n382));
  AND4_X1   g0182(.A1(new_n373), .A2(new_n382), .A3(new_n326), .A4(new_n377), .ZN(new_n383));
  OAI21_X1  g0183(.A(G200), .B1(new_n383), .B2(new_n378), .ZN(new_n384));
  OAI22_X1  g0184(.A1(new_n291), .A2(new_n207), .B1(new_n221), .B2(G68), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n346), .A2(new_n202), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n300), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT11), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n387), .A2(new_n388), .B1(new_n305), .B2(new_n211), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n387), .A2(new_n388), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n302), .A2(G68), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n391), .B(KEYINPUT12), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n381), .A2(new_n384), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(G169), .B1(new_n383), .B2(new_n378), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT80), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(KEYINPUT14), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(KEYINPUT14), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n379), .A2(G179), .A3(new_n380), .ZN(new_n402));
  OAI211_X1 g0202(.A(G169), .B(new_n398), .C1(new_n383), .C2(new_n378), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n400), .A2(new_n401), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n393), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n395), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT7), .B1(new_n257), .B2(new_n221), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n333), .A2(KEYINPUT7), .A3(new_n221), .A4(new_n334), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(G68), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT81), .B1(G58), .B2(G68), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(KEYINPUT81), .A2(G58), .A3(G68), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(new_n413), .C1(G58), .C2(G68), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(G20), .B1(G159), .B2(new_n285), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT82), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n410), .B(new_n415), .C1(new_n416), .C2(KEYINPUT16), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT16), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n285), .A2(G159), .ZN(new_n419));
  AND3_X1   g0219(.A1(KEYINPUT81), .A2(G58), .A3(G68), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n420), .A2(new_n411), .A3(new_n201), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n416), .B(new_n419), .C1(new_n421), .C2(new_n221), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n333), .A2(new_n221), .A3(new_n334), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT7), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n211), .B1(new_n425), .B2(new_n408), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n419), .B1(new_n421), .B2(new_n221), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n418), .B(new_n422), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n417), .A2(new_n428), .A3(new_n300), .ZN(new_n429));
  INV_X1    g0229(.A(new_n292), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(new_n302), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n306), .B2(new_n430), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(G226), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n434));
  OAI211_X1 g0234(.A(G223), .B(new_n260), .C1(new_n255), .C2(new_n256), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G87), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n265), .A2(new_n437), .B1(new_n279), .B2(new_n271), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n277), .A2(G232), .ZN(new_n439));
  AOI21_X1  g0239(.A(G200), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n265), .ZN(new_n441));
  AND4_X1   g0241(.A1(new_n358), .A2(new_n441), .A3(new_n326), .A4(new_n439), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT17), .B1(new_n433), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n326), .A3(new_n439), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n254), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n438), .A2(new_n358), .A3(new_n439), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT17), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(new_n429), .A4(new_n432), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT84), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n445), .A2(G169), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n438), .A2(G179), .A3(new_n439), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n429), .A2(KEYINPUT83), .A3(new_n432), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT83), .B1(new_n429), .B2(new_n432), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT18), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n444), .A2(KEYINPUT84), .A3(new_n450), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT18), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(new_n456), .C1(new_n457), .C2(new_n458), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n453), .A2(new_n460), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n367), .A2(new_n372), .A3(new_n406), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT24), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n221), .A2(G33), .A3(G116), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT23), .ZN(new_n469));
  INV_X1    g0269(.A(G107), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(G20), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(KEYINPUT73), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT73), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G107), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n221), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n468), .B(new_n471), .C1(new_n475), .C2(new_n469), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT89), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT23), .B1(new_n330), .B2(new_n221), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n479), .A2(KEYINPUT89), .A3(new_n468), .A4(new_n471), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n221), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n335), .A2(KEYINPUT22), .A3(new_n221), .A4(G87), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT88), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT88), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n481), .A2(new_n490), .A3(new_n487), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n467), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n490), .B1(new_n481), .B2(new_n487), .ZN(new_n493));
  AOI211_X1 g0293(.A(KEYINPUT88), .B(new_n486), .C1(new_n478), .C2(new_n480), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT24), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n300), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n302), .A2(G107), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT25), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n299), .B(new_n302), .C1(G1), .C2(new_n288), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(G107), .B1(new_n498), .B2(new_n497), .ZN(new_n503));
  OAI21_X1  g0303(.A(KEYINPUT90), .B1(new_n337), .B2(new_n214), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n335), .A2(G250), .A3(new_n260), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G294), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n260), .B1(new_n333), .B2(new_n334), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT90), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n508), .A3(G257), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n504), .A2(new_n505), .A3(new_n506), .A4(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n220), .B(G45), .C1(new_n269), .C2(KEYINPUT5), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(KEYINPUT5), .B2(new_n269), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n272), .B2(new_n276), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n510), .A2(new_n265), .B1(G264), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT87), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n269), .A2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g0316(.A(new_n276), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n274), .B1(new_n273), .B2(new_n275), .ZN(new_n518));
  OAI211_X1 g0318(.A(G274), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT86), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n511), .B(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n515), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n511), .B(KEYINPUT86), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n523), .A2(KEYINPUT87), .A3(new_n279), .A4(new_n516), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n514), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n254), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(G190), .B2(new_n526), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n496), .A2(new_n500), .A3(new_n503), .A4(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n302), .A2(G97), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n470), .A2(KEYINPUT6), .A3(G97), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n213), .A2(new_n470), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n531), .B1(new_n534), .B2(KEYINPUT6), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G20), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n330), .B1(new_n407), .B2(new_n409), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n285), .A2(G77), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n530), .B1(new_n539), .B2(new_n300), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n502), .A2(G97), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(G244), .B(new_n260), .C1(new_n255), .C2(new_n256), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT85), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT4), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n507), .A2(G250), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT4), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(KEYINPUT85), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G283), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n545), .A2(new_n546), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n265), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n513), .A2(G257), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n525), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G200), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n551), .A2(new_n525), .A3(G190), .A4(new_n552), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n542), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n507), .A2(G244), .B1(G33), .B2(G116), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n335), .A2(G238), .A3(new_n260), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n265), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n220), .A2(KEYINPUT68), .A3(G45), .A4(G274), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n220), .A2(G45), .ZN(new_n562));
  OAI211_X1 g0362(.A(G250), .B(new_n562), .C1(new_n517), .C2(new_n518), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n560), .A2(G190), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n291), .B2(new_n213), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n335), .A2(new_n221), .A3(G68), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n330), .A2(G87), .A3(G97), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n374), .A2(new_n565), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n569), .A2(G20), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(new_n300), .B1(new_n347), .B2(new_n303), .ZN(new_n572));
  INV_X1    g0372(.A(new_n265), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n557), .B2(new_n558), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n563), .A2(new_n561), .ZN(new_n575));
  OAI21_X1  g0375(.A(G200), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n502), .A2(G87), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n564), .A2(new_n572), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n571), .A2(new_n300), .ZN(new_n579));
  OR2_X1    g0379(.A1(new_n501), .A2(new_n347), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n347), .A2(new_n303), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G179), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n560), .A2(new_n583), .A3(new_n561), .A4(new_n563), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n343), .B1(new_n574), .B2(new_n575), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n578), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n553), .A2(new_n343), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n551), .A2(new_n525), .A3(new_n583), .A4(new_n552), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n540), .A2(new_n541), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n556), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n529), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n513), .A2(G270), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n507), .A2(G264), .B1(new_n257), .B2(G303), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n214), .B2(new_n336), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n265), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n525), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n303), .A2(new_n248), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n502), .A2(G116), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n299), .B1(G20), .B2(new_n248), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n549), .B(new_n221), .C1(G33), .C2(new_n213), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n601), .A2(KEYINPUT20), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT20), .B1(new_n601), .B2(new_n602), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n599), .B(new_n600), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n598), .A2(new_n605), .A3(G169), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n605), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n525), .A2(new_n597), .A3(G190), .A4(new_n594), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n525), .A2(new_n594), .A3(new_n597), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n254), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(G179), .A3(new_n605), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n598), .A2(new_n605), .A3(KEYINPUT21), .A4(G169), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n608), .A2(new_n612), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n489), .A2(new_n467), .A3(new_n491), .ZN(new_n616));
  OAI21_X1  g0416(.A(KEYINPUT24), .B1(new_n493), .B2(new_n494), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n299), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n503), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n618), .A2(new_n499), .A3(new_n619), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n526), .A2(KEYINPUT91), .A3(new_n583), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT91), .B1(new_n526), .B2(G169), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n526), .A2(new_n583), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n621), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n615), .B1(new_n620), .B2(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n466), .A2(new_n593), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g0428(.A(new_n628), .B(KEYINPUT92), .Z(G372));
  AOI221_X4 g0429(.A(new_n462), .B1(new_n454), .B2(new_n455), .C1(new_n429), .C2(new_n432), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT18), .B1(new_n433), .B2(new_n456), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n354), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n404), .A2(new_n405), .B1(new_n633), .B2(new_n394), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n453), .A2(new_n461), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n356), .B1(new_n636), .B2(new_n325), .ZN(new_n637));
  XOR2_X1   g0437(.A(new_n637), .B(KEYINPUT94), .Z(new_n638));
  NAND3_X1  g0438(.A1(new_n608), .A2(new_n613), .A3(new_n614), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n496), .A2(new_n500), .A3(new_n503), .ZN(new_n640));
  INV_X1    g0440(.A(new_n621), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n624), .B2(new_n622), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n639), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n586), .B1(new_n643), .B2(new_n593), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT93), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n590), .A2(new_n589), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n587), .A2(new_n646), .A3(new_n588), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n578), .A2(new_n586), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n591), .B2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n587), .A2(new_n646), .A3(KEYINPUT26), .A4(new_n588), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n649), .B1(new_n645), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n644), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n638), .B1(new_n466), .B2(new_n655), .ZN(G369));
  NOR2_X1   g0456(.A1(new_n620), .A2(new_n626), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G13), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G20), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n220), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n639), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n658), .A2(new_n529), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n658), .A2(new_n529), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n620), .A2(new_n667), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n670), .A2(new_n671), .B1(new_n658), .B2(new_n667), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n669), .B1(new_n672), .B2(new_n668), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n609), .A2(new_n667), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n639), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n612), .A2(new_n608), .A3(new_n613), .A4(new_n614), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n674), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n657), .A2(new_n667), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n669), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n227), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G1), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n568), .A2(new_n248), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n687), .A2(new_n688), .B1(new_n230), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n667), .B1(new_n644), .B2(new_n654), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(KEYINPUT96), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT29), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT96), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n694), .B(new_n667), .C1(new_n644), .C2(new_n654), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n653), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n667), .B1(new_n644), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT29), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G330), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n574), .A2(new_n575), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n611), .A2(G179), .A3(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n514), .A2(new_n552), .A3(new_n525), .A4(new_n551), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n706), .B1(new_n703), .B2(new_n704), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n611), .A2(G179), .ZN(new_n709));
  INV_X1    g0509(.A(new_n702), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(new_n710), .A3(new_n553), .A4(new_n526), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n666), .B1(new_n707), .B2(new_n712), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n627), .A2(new_n593), .A3(new_n666), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n712), .A2(KEYINPUT95), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n705), .A2(new_n706), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT95), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n708), .A2(new_n711), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n666), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n701), .B1(new_n716), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n700), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n690), .B1(new_n726), .B2(G1), .ZN(G364));
  AOI21_X1  g0527(.A(new_n220), .B1(new_n660), .B2(G45), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n685), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n677), .B2(G330), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G330), .B2(new_n677), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n231), .B1(G20), .B2(new_n343), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n733), .B(KEYINPUT98), .Z(new_n734));
  NOR2_X1   g0534(.A1(new_n221), .A2(new_n583), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n736), .A2(new_n358), .A3(G200), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G322), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n736), .A2(G190), .A3(G200), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G311), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n738), .A2(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n735), .A2(new_n358), .A3(G200), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT99), .Z(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(KEYINPUT33), .B(G317), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(G20), .A2(G190), .A3(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n583), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G326), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n749), .A2(G179), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G303), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n221), .A2(G190), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(new_n583), .A3(new_n254), .ZN(new_n755));
  INV_X1    g0555(.A(G329), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n754), .A2(new_n583), .A3(G200), .ZN(new_n757));
  INV_X1    g0557(.A(G283), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n755), .A2(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n358), .A2(G179), .A3(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n221), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n335), .B(new_n759), .C1(G294), .C2(new_n762), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n748), .A2(new_n751), .A3(new_n753), .A4(new_n763), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n738), .A2(new_n217), .B1(new_n741), .B2(new_n207), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n746), .B2(G68), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n750), .A2(G50), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n761), .A2(new_n213), .ZN(new_n768));
  INV_X1    g0568(.A(new_n752), .ZN(new_n769));
  INV_X1    g0569(.A(G87), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n757), .A2(new_n470), .ZN(new_n772));
  NOR4_X1   g0572(.A1(new_n768), .A2(new_n771), .A3(new_n772), .A4(new_n257), .ZN(new_n773));
  INV_X1    g0573(.A(G159), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n755), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT32), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n766), .A2(new_n767), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n734), .B1(new_n764), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n230), .A2(G45), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n252), .A2(new_n270), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT97), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n684), .A2(new_n335), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n782), .B(new_n783), .C1(new_n781), .C2(new_n780), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n684), .A2(new_n257), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G355), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n784), .B(new_n786), .C1(G116), .C2(new_n227), .ZN(new_n787));
  INV_X1    g0587(.A(new_n734), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G13), .A2(G33), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n778), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n791), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n793), .B(new_n730), .C1(new_n677), .C2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n732), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  NOR2_X1   g0597(.A1(new_n354), .A2(new_n666), .ZN(new_n798));
  INV_X1    g0598(.A(new_n353), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n364), .B1(new_n799), .B2(new_n667), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n798), .B1(new_n800), .B2(new_n354), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n667), .B(new_n801), .C1(new_n644), .C2(new_n654), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n692), .A2(new_n695), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n803), .B2(new_n801), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n804), .A2(new_n724), .ZN(new_n805));
  INV_X1    g0605(.A(new_n730), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n724), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G143), .A2(new_n737), .B1(new_n740), .B2(G159), .ZN(new_n809));
  INV_X1    g0609(.A(G137), .ZN(new_n810));
  INV_X1    g0610(.A(new_n750), .ZN(new_n811));
  INV_X1    g0611(.A(G150), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n809), .B1(new_n810), .B2(new_n811), .C1(new_n745), .C2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT34), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n761), .A2(new_n217), .B1(new_n757), .B2(new_n211), .ZN(new_n815));
  INV_X1    g0615(.A(new_n755), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n257), .B(new_n815), .C1(G132), .C2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n814), .B(new_n817), .C1(new_n202), .C2(new_n769), .ZN(new_n818));
  INV_X1    g0618(.A(G303), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n741), .A2(new_n248), .B1(new_n811), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n746), .B2(G283), .ZN(new_n821));
  INV_X1    g0621(.A(G294), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n257), .B1(new_n738), .B2(new_n822), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n755), .A2(new_n742), .B1(new_n757), .B2(new_n770), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n823), .A2(new_n768), .A3(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n821), .B(new_n825), .C1(new_n470), .C2(new_n769), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n734), .B1(new_n818), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n788), .A2(new_n789), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n827), .B1(new_n207), .B2(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n829), .B(new_n730), .C1(new_n790), .C2(new_n801), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n808), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G384));
  NOR2_X1   g0632(.A1(new_n393), .A2(new_n667), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n406), .B(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n712), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n667), .B1(new_n718), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n556), .A2(new_n587), .A3(new_n591), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n620), .B2(new_n528), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n676), .B1(new_n640), .B2(new_n642), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n839), .A2(new_n840), .A3(new_n667), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n837), .B1(new_n841), .B2(KEYINPUT31), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n713), .A2(new_n715), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n835), .B(new_n801), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n664), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n457), .A2(new_n458), .B1(new_n456), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n429), .A2(new_n432), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT37), .B1(new_n848), .B2(new_n448), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n410), .A2(new_n415), .A3(KEYINPUT16), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n418), .B1(new_n426), .B2(new_n427), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n850), .A2(new_n851), .A3(new_n300), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n432), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n456), .B2(new_n846), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n448), .A2(new_n432), .A3(new_n429), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n847), .A2(new_n849), .B1(new_n856), .B2(KEYINPUT37), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n664), .B1(new_n852), .B2(new_n432), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(new_n464), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n859), .A2(KEYINPUT38), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n861), .B(new_n857), .C1(new_n464), .C2(new_n858), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT102), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n859), .A2(KEYINPUT102), .A3(KEYINPUT38), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT40), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n845), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n464), .A2(new_n858), .ZN(new_n869));
  INV_X1    g0669(.A(new_n857), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT105), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n859), .A2(KEYINPUT105), .A3(KEYINPUT38), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT104), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n846), .B1(new_n457), .B2(new_n458), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n433), .A2(new_n456), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT103), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n448), .A2(new_n878), .A3(new_n429), .A4(new_n432), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT103), .B1(new_n433), .B2(new_n443), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n876), .A2(new_n877), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .B1(new_n849), .B2(new_n847), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n876), .B1(new_n632), .B2(new_n451), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n875), .B(new_n861), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n880), .A2(new_n877), .A3(new_n879), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT83), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n433), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n429), .A2(KEYINPUT83), .A3(new_n432), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n664), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT37), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n847), .A2(new_n849), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n449), .B1(new_n848), .B2(new_n448), .ZN(new_n892));
  INV_X1    g0692(.A(new_n450), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n892), .A2(new_n893), .B1(new_n630), .B2(new_n631), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n890), .A2(new_n891), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT104), .B1(new_n895), .B2(KEYINPUT38), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n873), .A2(new_n874), .B1(new_n884), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT40), .B1(new_n844), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n868), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(G330), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n372), .A2(new_n406), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n464), .B1(new_n365), .B2(new_n366), .ZN(new_n902));
  INV_X1    g0702(.A(new_n843), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n716), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n901), .A2(G330), .A3(new_n902), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT106), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n842), .A2(new_n843), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n466), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n907), .B1(new_n909), .B2(new_n899), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT39), .B1(new_n864), .B2(new_n865), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n896), .A2(new_n884), .ZN(new_n912));
  AND4_X1   g0712(.A1(KEYINPUT105), .A2(new_n869), .A3(KEYINPUT38), .A4(new_n870), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT105), .B1(new_n859), .B2(KEYINPUT38), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n404), .A2(new_n405), .A3(new_n667), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n911), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n406), .B(new_n833), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n798), .B(KEYINPUT101), .Z(new_n922));
  AOI21_X1  g0722(.A(new_n921), .B1(new_n802), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n866), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n632), .A2(new_n846), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n920), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n466), .B1(new_n696), .B2(new_n699), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n637), .B(KEYINPUT94), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n927), .B(new_n930), .Z(new_n931));
  XNOR2_X1  g0731(.A(new_n910), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n220), .B2(new_n660), .ZN(new_n933));
  OAI211_X1 g0733(.A(G20), .B(new_n273), .C1(new_n535), .C2(KEYINPUT35), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n248), .B(new_n934), .C1(KEYINPUT35), .C2(new_n535), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT36), .Z(new_n936));
  NOR4_X1   g0736(.A1(new_n411), .A2(new_n420), .A3(new_n230), .A4(new_n207), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n211), .A2(G50), .ZN(new_n938));
  OAI211_X1 g0738(.A(G1), .B(new_n659), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT100), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n933), .A2(new_n936), .A3(new_n940), .ZN(G367));
  OAI211_X1 g0741(.A(new_n556), .B(new_n591), .C1(new_n542), .C2(new_n667), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n646), .A2(new_n588), .A3(new_n666), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n669), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT42), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n591), .B1(new_n658), .B2(new_n942), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n667), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n572), .A2(new_n577), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n666), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n587), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n586), .B2(new_n950), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n946), .A2(new_n948), .B1(KEYINPUT43), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n944), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n679), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n953), .B(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n956), .B(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n673), .B(new_n678), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n682), .A2(new_n954), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT44), .Z(new_n962));
  NAND2_X1  g0762(.A1(new_n682), .A2(new_n954), .ZN(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n726), .B(new_n960), .C1(new_n962), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n726), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n685), .B(KEYINPUT41), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n958), .B1(new_n969), .B2(new_n729), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n738), .A2(new_n812), .B1(new_n769), .B2(new_n217), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n746), .B2(G159), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n750), .A2(G143), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n740), .A2(G50), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n757), .A2(new_n207), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n335), .B1(new_n755), .B2(new_n810), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n975), .B(new_n976), .C1(G68), .C2(new_n762), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n972), .A2(new_n973), .A3(new_n974), .A4(new_n977), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n257), .B1(new_n742), .B2(new_n811), .C1(new_n741), .C2(new_n758), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G294), .B2(new_n746), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n752), .A2(G116), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT46), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT108), .Z(new_n984));
  INV_X1    g0784(.A(new_n757), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(G97), .ZN(new_n986));
  INV_X1    g0786(.A(G317), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n986), .B1(new_n987), .B2(new_n755), .C1(new_n981), .C2(new_n982), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n330), .B2(new_n762), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n980), .A2(new_n984), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n738), .A2(new_n819), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n978), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT109), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT47), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n806), .B1(new_n994), .B2(new_n788), .ZN(new_n995));
  INV_X1    g0795(.A(new_n783), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n792), .B1(new_n227), .B2(new_n347), .C1(new_n238), .C2(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n995), .B(new_n997), .C1(new_n794), .C2(new_n952), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n970), .A2(new_n998), .ZN(G387));
  NAND2_X1  g0799(.A1(new_n726), .A2(new_n960), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n725), .A2(new_n959), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(new_n685), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n257), .B1(new_n757), .B2(new_n248), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n737), .A2(G317), .B1(new_n750), .B2(G322), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n819), .B2(new_n741), .C1(new_n745), .C2(new_n742), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT48), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n758), .B2(new_n761), .C1(new_n822), .C2(new_n769), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT49), .Z(new_n1008));
  AOI211_X1 g0808(.A(new_n1003), .B(new_n1008), .C1(G326), .C2(new_n816), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n740), .A2(G68), .B1(new_n750), .B2(G159), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n745), .B2(new_n292), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n761), .A2(new_n347), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(KEYINPUT111), .B(G150), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1012), .B1(new_n816), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n737), .A2(G50), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1014), .A2(new_n335), .A3(new_n986), .A4(new_n1015), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1011), .B(new_n1016), .C1(G77), .C2(new_n752), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n788), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n996), .B1(new_n243), .B2(G45), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n688), .B2(new_n785), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n292), .A2(G50), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n211), .B2(new_n207), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1023), .A2(G45), .A3(new_n688), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n1020), .A2(new_n1024), .B1(G107), .B2(new_n227), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n806), .B1(new_n1025), .B2(new_n792), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT110), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1018), .B(new_n1027), .C1(new_n672), .C2(new_n794), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1002), .B(new_n1028), .C1(new_n728), .C2(new_n959), .ZN(G393));
  NOR2_X1   g0829(.A1(new_n962), .A2(new_n965), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(KEYINPUT112), .B2(new_n680), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n680), .A2(KEYINPUT112), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n728), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n792), .B1(new_n213), .B2(new_n227), .C1(new_n249), .C2(new_n996), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n954), .A2(new_n794), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n257), .B1(new_n822), .B2(new_n741), .C1(new_n745), .C2(new_n819), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n737), .A2(G311), .B1(new_n750), .B2(G317), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT52), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n772), .B1(G116), .B2(new_n762), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n739), .B2(new_n755), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1039), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n758), .B2(new_n769), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n737), .A2(G159), .B1(new_n750), .B2(G150), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT51), .Z(new_n1047));
  NOR2_X1   g0847(.A1(new_n761), .A2(new_n207), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n257), .B(new_n1048), .C1(new_n430), .C2(new_n740), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n746), .A2(G50), .B1(G87), .B2(new_n985), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n816), .A2(G143), .B1(G68), .B2(new_n752), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT113), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1045), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT114), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n806), .B(new_n1038), .C1(new_n788), .C2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1036), .B1(new_n1037), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1034), .A2(new_n1000), .A3(new_n1035), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1058), .A2(new_n685), .A3(new_n966), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(G390));
  NAND2_X1  g0860(.A1(new_n716), .A2(new_n722), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1061), .A2(G330), .A3(new_n801), .A4(new_n835), .ZN(new_n1062));
  OAI211_X1 g0862(.A(G330), .B(new_n801), .C1(new_n842), .C2(new_n843), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n921), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n667), .B(new_n801), .C1(new_n644), .C2(new_n697), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1065), .A2(new_n922), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1062), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n904), .A2(G330), .A3(new_n801), .A4(new_n835), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n666), .ZN(new_n1069));
  OAI211_X1 g0869(.A(G330), .B(new_n801), .C1(new_n842), .C2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n921), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n802), .A2(new_n922), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1067), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n466), .A2(new_n701), .A3(new_n908), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n928), .A2(new_n1076), .A3(new_n929), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1068), .A2(KEYINPUT115), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1073), .A2(new_n835), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n911), .A2(new_n917), .B1(new_n1080), .B2(new_n918), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n921), .B1(new_n1065), .B2(new_n922), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n1082), .A2(new_n897), .A3(new_n919), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1079), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1070), .A2(new_n921), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT115), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1085), .B1(new_n1068), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n873), .A2(new_n874), .ZN(new_n1088));
  AOI21_X1  g0888(.A(KEYINPUT39), .B1(new_n1088), .B2(new_n912), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n869), .A2(new_n870), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n861), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n863), .B1(new_n859), .B2(KEYINPUT38), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n865), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n916), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1089), .A2(new_n1095), .B1(new_n923), .B2(new_n919), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n918), .B(new_n915), .C1(new_n1066), .C2(new_n921), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1087), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1084), .A2(new_n1098), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1078), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1078), .A2(new_n1099), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(new_n685), .A3(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1099), .A2(new_n728), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n789), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n738), .A2(new_n248), .B1(new_n811), .B2(new_n758), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n746), .B2(new_n330), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n740), .A2(G97), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n335), .B1(new_n985), .B2(G68), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n771), .B(new_n1048), .C1(G294), .C2(new_n816), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  XOR2_X1   g0910(.A(KEYINPUT54), .B(G143), .Z(new_n1111));
  AOI21_X1  g0911(.A(new_n257), .B1(new_n740), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(G132), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1112), .B1(new_n1113), .B2(new_n738), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1013), .A2(new_n752), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT53), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1114), .B(new_n1116), .C1(G137), .C2(new_n746), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n762), .A2(G159), .B1(new_n816), .B2(G125), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(new_n202), .C2(new_n757), .ZN(new_n1119));
  INV_X1    g0919(.A(G128), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n811), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1110), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1122), .A2(new_n788), .B1(new_n292), .B2(new_n828), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1104), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1103), .B1(new_n730), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1102), .A2(new_n1125), .ZN(G378));
  INV_X1    g0926(.A(KEYINPUT56), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n371), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n308), .A2(new_n846), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT55), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1131), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1127), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1135), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(KEYINPUT56), .A3(new_n1133), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n701), .B1(new_n868), .B2(new_n898), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1140), .A2(new_n927), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n927), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1139), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n927), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n900), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1139), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1140), .A2(new_n927), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1143), .A2(new_n1148), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1062), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1074), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1077), .B1(new_n1099), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT118), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(KEYINPUT118), .B(new_n1077), .C1(new_n1099), .C2(new_n1152), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1149), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT57), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1149), .A2(new_n1155), .A3(KEYINPUT57), .A4(new_n1156), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n685), .A3(new_n1160), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n788), .A2(G50), .A3(new_n789), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n745), .A2(new_n213), .B1(new_n347), .B2(new_n741), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT116), .Z(new_n1164));
  AOI22_X1  g0964(.A1(new_n737), .A2(G107), .B1(new_n750), .B2(G116), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n207), .B2(new_n769), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n757), .A2(new_n217), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n1166), .A2(G41), .A3(new_n335), .A4(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n762), .A2(G68), .B1(new_n816), .B2(G283), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1164), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT58), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n202), .B1(new_n255), .B2(G41), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n741), .A2(new_n810), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1111), .A2(new_n752), .B1(G125), .B2(new_n750), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1174), .B1(new_n812), .B2(new_n761), .C1(new_n738), .C2(new_n1120), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(G132), .C2(new_n746), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT59), .ZN(new_n1177));
  AOI21_X1  g0977(.A(G41), .B1(new_n816), .B2(G124), .ZN(new_n1178));
  AOI21_X1  g0978(.A(G33), .B1(new_n985), .B2(G159), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1171), .A2(new_n1172), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n788), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n730), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1162), .B(new_n1183), .C1(new_n1146), .C2(new_n789), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1184), .A2(KEYINPUT117), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(KEYINPUT117), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1185), .A2(new_n1186), .B1(new_n729), .B2(new_n1149), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1161), .A2(new_n1187), .ZN(G375));
  OAI211_X1 g0988(.A(new_n638), .B(new_n905), .C1(new_n700), .C2(new_n466), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1152), .A2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n968), .B(KEYINPUT119), .Z(new_n1191));
  NAND3_X1  g0991(.A1(new_n1078), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n738), .A2(new_n758), .B1(new_n769), .B2(new_n213), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n746), .B2(G116), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n740), .A2(new_n330), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n335), .B1(new_n750), .B2(G294), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n975), .B(new_n1012), .C1(G303), .C2(new_n816), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n738), .A2(new_n810), .B1(new_n811), .B2(new_n1113), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n746), .B2(new_n1111), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1167), .A2(new_n257), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n761), .A2(new_n202), .B1(new_n755), .B2(new_n1120), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G150), .B2(new_n740), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n769), .A2(new_n774), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1198), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1206), .A2(new_n788), .B1(new_n211), .B2(new_n828), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n730), .B(new_n1207), .C1(new_n835), .C2(new_n790), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n1152), .B2(new_n728), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1192), .A2(new_n1210), .ZN(G381));
  INV_X1    g1011(.A(KEYINPUT121), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(G375), .A2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(G393), .A2(G396), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT120), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(G378), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1102), .A2(new_n1125), .A3(KEYINPUT120), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1161), .A2(KEYINPUT121), .A3(new_n1187), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1213), .A2(new_n1214), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(G390), .A2(G387), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1221), .A2(new_n831), .A3(new_n1210), .A4(new_n1192), .ZN(new_n1222));
  OR3_X1    g1022(.A1(new_n1220), .A2(new_n1222), .A3(KEYINPUT122), .ZN(new_n1223));
  OAI21_X1  g1023(.A(KEYINPUT122), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(G407));
  NAND4_X1  g1025(.A1(new_n1213), .A2(new_n665), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(G407), .A2(G213), .A3(new_n1226), .ZN(G409));
  OR2_X1    g1027(.A1(G390), .A2(G387), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(G390), .A2(G387), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(G393), .B(new_n796), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(KEYINPUT126), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1230), .A2(KEYINPUT126), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1228), .B(new_n1229), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1229), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1231), .B1(new_n1235), .B2(new_n1221), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1152), .A2(KEYINPUT60), .A3(new_n1189), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n685), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT60), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT123), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT60), .B1(new_n1152), .B2(new_n1189), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT123), .B1(new_n1246), .B2(new_n1190), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1240), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT124), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1244), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1246), .A2(KEYINPUT123), .A3(new_n1190), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(new_n1253), .A3(new_n1240), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1249), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G384), .B1(new_n1255), .B2(new_n1210), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1253), .B1(new_n1252), .B2(new_n1240), .ZN(new_n1257));
  AOI211_X1 g1057(.A(KEYINPUT124), .B(new_n1239), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G384), .B(new_n1210), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1161), .A2(G378), .A3(new_n1187), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1184), .B1(new_n1149), .B2(new_n729), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1191), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1157), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1218), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n665), .A2(G213), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1261), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1262), .A2(new_n1266), .B1(G213), .B2(new_n665), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT62), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1273), .A3(new_n1261), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1210), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n831), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1259), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n665), .A2(G213), .A3(G2897), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1278), .A2(new_n1259), .A3(new_n1280), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1276), .B1(new_n1284), .B2(new_n1272), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1237), .B1(new_n1275), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT125), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1269), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT63), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1278), .A2(new_n1259), .A3(new_n1280), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1280), .B1(new_n1278), .B2(new_n1259), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1272), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT61), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1269), .A2(new_n1287), .A3(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1289), .A2(new_n1294), .A3(new_n1295), .A4(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1286), .A2(new_n1298), .ZN(G405));
  NAND2_X1  g1099(.A1(G375), .A2(new_n1218), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1262), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(new_n1261), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(new_n1237), .ZN(G402));
endmodule


