

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  INV_X1 U322 ( .A(KEYINPUT91), .ZN(n396) );
  XOR2_X1 U323 ( .A(n377), .B(n402), .Z(n449) );
  XNOR2_X1 U324 ( .A(n373), .B(n372), .ZN(n377) );
  XNOR2_X1 U325 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U326 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U327 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n444) );
  XNOR2_X1 U328 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U329 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U330 ( .A(n441), .B(n393), .Z(n290) );
  XNOR2_X1 U331 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n386) );
  INV_X1 U332 ( .A(KEYINPUT22), .ZN(n428) );
  XNOR2_X1 U333 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U334 ( .A(n390), .B(KEYINPUT48), .ZN(n523) );
  XNOR2_X1 U335 ( .A(n431), .B(n430), .ZN(n433) );
  INV_X1 U336 ( .A(KEYINPUT37), .ZN(n467) );
  XNOR2_X1 U337 ( .A(n437), .B(n436), .ZN(n438) );
  NOR2_X1 U338 ( .A1(n426), .A2(n511), .ZN(n427) );
  INV_X1 U339 ( .A(n523), .ZN(n525) );
  XNOR2_X1 U340 ( .A(n439), .B(n438), .ZN(n443) );
  XNOR2_X1 U341 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U342 ( .A(n403), .B(n402), .ZN(n513) );
  XNOR2_X1 U343 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n447) );
  XNOR2_X1 U344 ( .A(n474), .B(G43GAT), .ZN(n475) );
  XNOR2_X1 U345 ( .A(n448), .B(n447), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n476), .B(n475), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n292) );
  XNOR2_X1 U348 ( .A(KEYINPUT11), .B(KEYINPUT76), .ZN(n291) );
  XNOR2_X1 U349 ( .A(n292), .B(n291), .ZN(n302) );
  XOR2_X1 U350 ( .A(G99GAT), .B(G85GAT), .Z(n367) );
  XOR2_X1 U351 ( .A(KEYINPUT10), .B(n367), .Z(n294) );
  XOR2_X1 U352 ( .A(G50GAT), .B(G162GAT), .Z(n432) );
  XNOR2_X1 U353 ( .A(G218GAT), .B(n432), .ZN(n293) );
  XNOR2_X1 U354 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U355 ( .A(G92GAT), .B(G106GAT), .Z(n296) );
  NAND2_X1 U356 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U357 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U358 ( .A(n298), .B(n297), .Z(n300) );
  XOR2_X1 U359 ( .A(G36GAT), .B(G190GAT), .Z(n393) );
  XNOR2_X1 U360 ( .A(G134GAT), .B(n393), .ZN(n299) );
  XNOR2_X1 U361 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U362 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U363 ( .A(KEYINPUT7), .B(KEYINPUT67), .Z(n304) );
  XNOR2_X1 U364 ( .A(G43GAT), .B(G29GAT), .ZN(n303) );
  XNOR2_X1 U365 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U366 ( .A(KEYINPUT8), .B(n305), .ZN(n336) );
  XNOR2_X1 U367 ( .A(n306), .B(n336), .ZN(n552) );
  XOR2_X1 U368 ( .A(G190GAT), .B(G43GAT), .Z(n308) );
  NAND2_X1 U369 ( .A1(G227GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U370 ( .A(n308), .B(n307), .ZN(n311) );
  XOR2_X1 U371 ( .A(G127GAT), .B(KEYINPUT0), .Z(n310) );
  XNOR2_X1 U372 ( .A(G113GAT), .B(G134GAT), .ZN(n309) );
  XNOR2_X1 U373 ( .A(n310), .B(n309), .ZN(n405) );
  XOR2_X1 U374 ( .A(n311), .B(n405), .Z(n319) );
  XOR2_X1 U375 ( .A(G176GAT), .B(G120GAT), .Z(n313) );
  XNOR2_X1 U376 ( .A(G169GAT), .B(G99GAT), .ZN(n312) );
  XNOR2_X1 U377 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U378 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n315) );
  XNOR2_X1 U379 ( .A(G15GAT), .B(G71GAT), .ZN(n314) );
  XNOR2_X1 U380 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U381 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U382 ( .A(n319), .B(n318), .ZN(n324) );
  XOR2_X1 U383 ( .A(G183GAT), .B(KEYINPUT80), .Z(n321) );
  XNOR2_X1 U384 ( .A(KEYINPUT19), .B(KEYINPUT81), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n321), .B(n320), .ZN(n323) );
  XOR2_X1 U386 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n322) );
  XOR2_X1 U387 ( .A(n323), .B(n322), .Z(n401) );
  XOR2_X1 U388 ( .A(n324), .B(n401), .Z(n528) );
  XOR2_X1 U389 ( .A(G169GAT), .B(G8GAT), .Z(n395) );
  XOR2_X1 U390 ( .A(G15GAT), .B(G22GAT), .Z(n326) );
  XNOR2_X1 U391 ( .A(G1GAT), .B(KEYINPUT68), .ZN(n325) );
  XNOR2_X1 U392 ( .A(n326), .B(n325), .ZN(n352) );
  XOR2_X1 U393 ( .A(n395), .B(n352), .Z(n328) );
  NAND2_X1 U394 ( .A1(G229GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U395 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U396 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n330) );
  XNOR2_X1 U397 ( .A(G197GAT), .B(KEYINPUT30), .ZN(n329) );
  XNOR2_X1 U398 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U399 ( .A(n332), .B(n331), .Z(n338) );
  XOR2_X1 U400 ( .A(G113GAT), .B(G141GAT), .Z(n334) );
  XNOR2_X1 U401 ( .A(G50GAT), .B(G36GAT), .ZN(n333) );
  XNOR2_X1 U402 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U403 ( .A(n336), .B(n335), .Z(n337) );
  XOR2_X1 U404 ( .A(n338), .B(n337), .Z(n541) );
  INV_X1 U405 ( .A(n541), .ZN(n567) );
  XNOR2_X1 U406 ( .A(KEYINPUT36), .B(KEYINPUT100), .ZN(n339) );
  XNOR2_X1 U407 ( .A(n339), .B(n552), .ZN(n576) );
  XOR2_X1 U408 ( .A(KEYINPUT78), .B(G211GAT), .Z(n341) );
  XNOR2_X1 U409 ( .A(G8GAT), .B(G183GAT), .ZN(n340) );
  XNOR2_X1 U410 ( .A(n341), .B(n340), .ZN(n356) );
  XOR2_X1 U411 ( .A(G64GAT), .B(G57GAT), .Z(n343) );
  XNOR2_X1 U412 ( .A(G127GAT), .B(G155GAT), .ZN(n342) );
  XNOR2_X1 U413 ( .A(n343), .B(n342), .ZN(n348) );
  XNOR2_X1 U414 ( .A(G71GAT), .B(KEYINPUT69), .ZN(n344) );
  XNOR2_X1 U415 ( .A(n344), .B(KEYINPUT13), .ZN(n364) );
  XOR2_X1 U416 ( .A(n364), .B(KEYINPUT12), .Z(n346) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U418 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U419 ( .A(n348), .B(n347), .Z(n354) );
  XOR2_X1 U420 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n350) );
  XNOR2_X1 U421 ( .A(G78GAT), .B(KEYINPUT14), .ZN(n349) );
  XNOR2_X1 U422 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U423 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U424 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U425 ( .A(n356), .B(n355), .ZN(n477) );
  INV_X1 U426 ( .A(n477), .ZN(n574) );
  NAND2_X1 U427 ( .A1(n576), .A2(n574), .ZN(n358) );
  XNOR2_X1 U428 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n357) );
  XNOR2_X1 U429 ( .A(n358), .B(n357), .ZN(n378) );
  XOR2_X1 U430 ( .A(KEYINPUT70), .B(KEYINPUT31), .Z(n360) );
  NAND2_X1 U431 ( .A1(G230GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U432 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U433 ( .A(n361), .B(KEYINPUT75), .Z(n366) );
  XOR2_X1 U434 ( .A(KEYINPUT72), .B(G78GAT), .Z(n363) );
  XNOR2_X1 U435 ( .A(G148GAT), .B(G106GAT), .ZN(n362) );
  XNOR2_X1 U436 ( .A(n363), .B(n362), .ZN(n440) );
  XNOR2_X1 U437 ( .A(n440), .B(n364), .ZN(n365) );
  XNOR2_X1 U438 ( .A(n366), .B(n365), .ZN(n373) );
  XOR2_X1 U439 ( .A(G120GAT), .B(G57GAT), .Z(n406) );
  XOR2_X1 U440 ( .A(n406), .B(n367), .Z(n371) );
  XOR2_X1 U441 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n369) );
  XNOR2_X1 U442 ( .A(KEYINPUT32), .B(KEYINPUT74), .ZN(n368) );
  XNOR2_X1 U443 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U444 ( .A(G92GAT), .B(G64GAT), .Z(n375) );
  XNOR2_X1 U445 ( .A(G176GAT), .B(G204GAT), .ZN(n374) );
  XNOR2_X1 U446 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U447 ( .A(KEYINPUT73), .B(n376), .ZN(n402) );
  NAND2_X1 U448 ( .A1(n378), .A2(n449), .ZN(n379) );
  NOR2_X1 U449 ( .A1(n567), .A2(n379), .ZN(n380) );
  XNOR2_X1 U450 ( .A(KEYINPUT115), .B(n380), .ZN(n389) );
  INV_X1 U451 ( .A(n449), .ZN(n570) );
  XOR2_X1 U452 ( .A(KEYINPUT41), .B(n570), .Z(n544) );
  NAND2_X1 U453 ( .A1(n544), .A2(n567), .ZN(n382) );
  INV_X1 U454 ( .A(KEYINPUT46), .ZN(n381) );
  XNOR2_X1 U455 ( .A(n382), .B(n381), .ZN(n383) );
  NOR2_X1 U456 ( .A1(n383), .A2(n574), .ZN(n384) );
  XNOR2_X1 U457 ( .A(n384), .B(KEYINPUT113), .ZN(n385) );
  NOR2_X1 U458 ( .A1(n552), .A2(n385), .ZN(n387) );
  XNOR2_X1 U459 ( .A(n387), .B(n386), .ZN(n388) );
  NAND2_X1 U460 ( .A1(n389), .A2(n388), .ZN(n390) );
  XOR2_X1 U461 ( .A(G211GAT), .B(KEYINPUT21), .Z(n392) );
  XNOR2_X1 U462 ( .A(G197GAT), .B(G218GAT), .ZN(n391) );
  XNOR2_X1 U463 ( .A(n392), .B(n391), .ZN(n441) );
  NAND2_X1 U464 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U465 ( .A(n290), .B(n394), .ZN(n399) );
  XNOR2_X1 U466 ( .A(n395), .B(KEYINPUT90), .ZN(n397) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n403) );
  NAND2_X1 U468 ( .A1(n523), .A2(n513), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n404), .B(KEYINPUT54), .ZN(n426) );
  XOR2_X1 U470 ( .A(n406), .B(n405), .Z(n408) );
  NAND2_X1 U471 ( .A1(G225GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U472 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U473 ( .A(n409), .B(G148GAT), .Z(n413) );
  XOR2_X1 U474 ( .A(G155GAT), .B(KEYINPUT2), .Z(n411) );
  XNOR2_X1 U475 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n411), .B(n410), .ZN(n431) );
  XNOR2_X1 U477 ( .A(n431), .B(KEYINPUT5), .ZN(n412) );
  XNOR2_X1 U478 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U479 ( .A(KEYINPUT86), .B(G85GAT), .Z(n415) );
  XNOR2_X1 U480 ( .A(G29GAT), .B(G162GAT), .ZN(n414) );
  XNOR2_X1 U481 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U482 ( .A(n417), .B(n416), .Z(n425) );
  XOR2_X1 U483 ( .A(KEYINPUT89), .B(KEYINPUT4), .Z(n419) );
  XNOR2_X1 U484 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n418) );
  XNOR2_X1 U485 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U486 ( .A(KEYINPUT85), .B(KEYINPUT6), .Z(n421) );
  XNOR2_X1 U487 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n420) );
  XNOR2_X1 U488 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U489 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n511) );
  XNOR2_X1 U491 ( .A(n427), .B(KEYINPUT64), .ZN(n565) );
  NAND2_X1 U492 ( .A1(G228GAT), .A2(G233GAT), .ZN(n429) );
  XOR2_X1 U493 ( .A(n433), .B(n432), .Z(n439) );
  XOR2_X1 U494 ( .A(KEYINPUT84), .B(KEYINPUT24), .Z(n435) );
  XNOR2_X1 U495 ( .A(KEYINPUT83), .B(KEYINPUT23), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U497 ( .A(G22GAT), .B(G204GAT), .ZN(n436) );
  XOR2_X1 U498 ( .A(n441), .B(n440), .Z(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n460) );
  NAND2_X1 U500 ( .A1(n565), .A2(n460), .ZN(n445) );
  NOR2_X1 U501 ( .A1(n528), .A2(n446), .ZN(n561) );
  NAND2_X1 U502 ( .A1(n552), .A2(n561), .ZN(n448) );
  NAND2_X1 U503 ( .A1(n567), .A2(n449), .ZN(n481) );
  INV_X1 U504 ( .A(n528), .ZN(n516) );
  NAND2_X1 U505 ( .A1(n516), .A2(n513), .ZN(n450) );
  XNOR2_X1 U506 ( .A(KEYINPUT94), .B(n450), .ZN(n451) );
  NAND2_X1 U507 ( .A1(n451), .A2(n460), .ZN(n452) );
  XNOR2_X1 U508 ( .A(KEYINPUT25), .B(n452), .ZN(n457) );
  NOR2_X1 U509 ( .A1(n460), .A2(n516), .ZN(n454) );
  XNOR2_X1 U510 ( .A(KEYINPUT26), .B(KEYINPUT92), .ZN(n453) );
  XNOR2_X1 U511 ( .A(n454), .B(n453), .ZN(n566) );
  XNOR2_X1 U512 ( .A(KEYINPUT27), .B(n513), .ZN(n461) );
  NAND2_X1 U513 ( .A1(n566), .A2(n461), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n455), .B(KEYINPUT93), .ZN(n456) );
  NOR2_X1 U515 ( .A1(n457), .A2(n456), .ZN(n458) );
  XOR2_X1 U516 ( .A(KEYINPUT95), .B(n458), .Z(n459) );
  NOR2_X1 U517 ( .A1(n511), .A2(n459), .ZN(n464) );
  XOR2_X1 U518 ( .A(n460), .B(KEYINPUT28), .Z(n519) );
  INV_X1 U519 ( .A(n519), .ZN(n526) );
  NAND2_X1 U520 ( .A1(n528), .A2(n526), .ZN(n462) );
  NAND2_X1 U521 ( .A1(n511), .A2(n461), .ZN(n524) );
  NOR2_X1 U522 ( .A1(n462), .A2(n524), .ZN(n463) );
  NOR2_X1 U523 ( .A1(n464), .A2(n463), .ZN(n465) );
  XOR2_X1 U524 ( .A(KEYINPUT96), .B(n465), .Z(n479) );
  NAND2_X1 U525 ( .A1(n479), .A2(n576), .ZN(n466) );
  NOR2_X1 U526 ( .A1(n574), .A2(n466), .ZN(n470) );
  XNOR2_X1 U527 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n470), .B(n469), .ZN(n510) );
  NOR2_X1 U529 ( .A1(n481), .A2(n510), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT38), .ZN(n495) );
  NAND2_X1 U531 ( .A1(n495), .A2(n513), .ZN(n473) );
  XNOR2_X1 U532 ( .A(G36GAT), .B(KEYINPUT104), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n473), .B(n472), .ZN(G1329GAT) );
  NAND2_X1 U534 ( .A1(n495), .A2(n516), .ZN(n476) );
  XOR2_X1 U535 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n474) );
  NOR2_X1 U536 ( .A1(n552), .A2(n477), .ZN(n478) );
  XNOR2_X1 U537 ( .A(KEYINPUT16), .B(n478), .ZN(n480) );
  NAND2_X1 U538 ( .A1(n480), .A2(n479), .ZN(n497) );
  NOR2_X1 U539 ( .A1(n481), .A2(n497), .ZN(n489) );
  NAND2_X1 U540 ( .A1(n489), .A2(n511), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT34), .ZN(n483) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U543 ( .A1(n513), .A2(n489), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT35), .B(KEYINPUT98), .Z(n486) );
  NAND2_X1 U546 ( .A1(n489), .A2(n516), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(n488) );
  XOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT97), .Z(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  NAND2_X1 U550 ( .A1(n489), .A2(n519), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U552 ( .A1(n495), .A2(n511), .ZN(n494) );
  XOR2_X1 U553 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n492) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT99), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n519), .A2(n495), .ZN(n496) );
  XNOR2_X1 U558 ( .A(G50GAT), .B(n496), .ZN(G1331GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n499) );
  XOR2_X1 U560 ( .A(n544), .B(KEYINPUT107), .Z(n558) );
  NAND2_X1 U561 ( .A1(n558), .A2(n541), .ZN(n509) );
  NOR2_X1 U562 ( .A1(n509), .A2(n497), .ZN(n504) );
  NAND2_X1 U563 ( .A1(n504), .A2(n511), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U565 ( .A(G57GAT), .B(n500), .Z(G1332GAT) );
  NAND2_X1 U566 ( .A1(n513), .A2(n504), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n501), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U568 ( .A1(n516), .A2(n504), .ZN(n502) );
  XNOR2_X1 U569 ( .A(n502), .B(KEYINPUT108), .ZN(n503) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(n503), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n506) );
  NAND2_X1 U572 ( .A1(n504), .A2(n519), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(n508) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT110), .Z(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  NOR2_X1 U576 ( .A1(n510), .A2(n509), .ZN(n520) );
  NAND2_X1 U577 ( .A1(n511), .A2(n520), .ZN(n512) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n512), .ZN(G1336GAT) );
  XOR2_X1 U579 ( .A(G92GAT), .B(KEYINPUT111), .Z(n515) );
  NAND2_X1 U580 ( .A1(n520), .A2(n513), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(G1337GAT) );
  NAND2_X1 U582 ( .A1(n516), .A2(n520), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(KEYINPUT112), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G99GAT), .B(n518), .ZN(G1338GAT) );
  NAND2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(KEYINPUT44), .ZN(n522) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  XNOR2_X1 U588 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n530) );
  NOR2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n540) );
  NAND2_X1 U590 ( .A1(n540), .A2(n526), .ZN(n527) );
  NOR2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n567), .A2(n537), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n530), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n532) );
  NAND2_X1 U595 ( .A1(n537), .A2(n558), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n534) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT117), .Z(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n537), .A2(n574), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n535), .B(KEYINPUT50), .ZN(n536) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U603 ( .A1(n537), .A2(n552), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U605 ( .A1(n566), .A2(n540), .ZN(n543) );
  NOR2_X1 U606 ( .A1(n541), .A2(n543), .ZN(n542) );
  XOR2_X1 U607 ( .A(G141GAT), .B(n542), .Z(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n546) );
  INV_X1 U609 ( .A(n543), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n551), .A2(n544), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U612 ( .A(n547), .B(KEYINPUT119), .Z(n549) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n551), .A2(n574), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U619 ( .A1(n561), .A2(n567), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n556) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(n557), .Z(n560) );
  NAND2_X1 U625 ( .A1(n558), .A2(n561), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n574), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(KEYINPUT60), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT59), .B(n564), .Z(n569) );
  AND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n577) );
  NAND2_X1 U633 ( .A1(n577), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U636 ( .A1(n577), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(G204GAT), .B(n573), .Z(G1353GAT) );
  NAND2_X1 U639 ( .A1(n577), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1355GAT) );
endmodule

