

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U546 ( .A1(n522), .A2(G2105), .ZN(n861) );
  INV_X2 U547 ( .A(G2104), .ZN(n522) );
  OR2_X1 U548 ( .A1(n693), .A2(n692), .ZN(n694) );
  OR2_X1 U549 ( .A1(n524), .A2(n510), .ZN(n525) );
  AND2_X1 U550 ( .A1(n862), .A2(G113), .ZN(n510) );
  XOR2_X1 U551 ( .A(KEYINPUT14), .B(n594), .Z(n511) );
  NOR2_X1 U552 ( .A1(n620), .A2(n619), .ZN(n632) );
  INV_X1 U553 ( .A(KEYINPUT96), .ZN(n646) );
  INV_X1 U554 ( .A(KEYINPUT97), .ZN(n649) );
  NOR2_X1 U555 ( .A1(G651), .A2(n568), .ZN(n776) );
  XOR2_X1 U556 ( .A(KEYINPUT68), .B(n596), .Z(n992) );
  NOR2_X1 U557 ( .A1(n526), .A2(n525), .ZN(n531) );
  XOR2_X1 U558 ( .A(G543), .B(KEYINPUT0), .Z(n568) );
  NAND2_X1 U559 ( .A1(G52), .A2(n776), .ZN(n514) );
  INV_X1 U560 ( .A(G651), .ZN(n515) );
  NOR2_X1 U561 ( .A1(G543), .A2(n515), .ZN(n512) );
  XOR2_X2 U562 ( .A(KEYINPUT1), .B(n512), .Z(n779) );
  NAND2_X1 U563 ( .A1(G64), .A2(n779), .ZN(n513) );
  NAND2_X1 U564 ( .A1(n514), .A2(n513), .ZN(n520) );
  NOR2_X1 U565 ( .A1(G651), .A2(G543), .ZN(n770) );
  NAND2_X1 U566 ( .A1(G90), .A2(n770), .ZN(n517) );
  NOR2_X1 U567 ( .A1(n568), .A2(n515), .ZN(n772) );
  NAND2_X1 U568 ( .A1(G77), .A2(n772), .ZN(n516) );
  NAND2_X1 U569 ( .A1(n517), .A2(n516), .ZN(n518) );
  XOR2_X1 U570 ( .A(KEYINPUT9), .B(n518), .Z(n519) );
  NOR2_X1 U571 ( .A1(n520), .A2(n519), .ZN(G171) );
  INV_X1 U572 ( .A(G171), .ZN(G301) );
  NOR2_X2 U573 ( .A1(G2105), .A2(n522), .ZN(n866) );
  NAND2_X1 U574 ( .A1(G101), .A2(n866), .ZN(n521) );
  XNOR2_X1 U575 ( .A(n521), .B(KEYINPUT23), .ZN(n526) );
  AND2_X1 U576 ( .A1(G125), .A2(n861), .ZN(n523) );
  XNOR2_X1 U577 ( .A(KEYINPUT64), .B(n523), .ZN(n524) );
  AND2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n862) );
  INV_X1 U579 ( .A(KEYINPUT65), .ZN(n529) );
  NOR2_X1 U580 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XOR2_X2 U581 ( .A(KEYINPUT17), .B(n527), .Z(n865) );
  NAND2_X1 U582 ( .A1(G137), .A2(n865), .ZN(n528) );
  XNOR2_X1 U583 ( .A(n529), .B(n528), .ZN(n530) );
  AND2_X2 U584 ( .A1(n531), .A2(n530), .ZN(G160) );
  NAND2_X1 U585 ( .A1(G138), .A2(n865), .ZN(n533) );
  NAND2_X1 U586 ( .A1(G102), .A2(n866), .ZN(n532) );
  NAND2_X1 U587 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U588 ( .A(KEYINPUT82), .B(n534), .ZN(n538) );
  NAND2_X1 U589 ( .A1(G126), .A2(n861), .ZN(n536) );
  NAND2_X1 U590 ( .A1(G114), .A2(n862), .ZN(n535) );
  NAND2_X1 U591 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U592 ( .A1(n538), .A2(n537), .ZN(G164) );
  NAND2_X1 U593 ( .A1(n770), .A2(G89), .ZN(n539) );
  XNOR2_X1 U594 ( .A(n539), .B(KEYINPUT4), .ZN(n541) );
  NAND2_X1 U595 ( .A1(G76), .A2(n772), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U597 ( .A(n542), .B(KEYINPUT5), .ZN(n547) );
  NAND2_X1 U598 ( .A1(G51), .A2(n776), .ZN(n544) );
  NAND2_X1 U599 ( .A1(G63), .A2(n779), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U601 ( .A(KEYINPUT6), .B(n545), .Z(n546) );
  NAND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U603 ( .A(n548), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U604 ( .A1(G88), .A2(n770), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G75), .A2(n772), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U607 ( .A1(G50), .A2(n776), .ZN(n552) );
  NAND2_X1 U608 ( .A1(G62), .A2(n779), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U610 ( .A1(n554), .A2(n553), .ZN(G166) );
  INV_X1 U611 ( .A(G166), .ZN(G303) );
  XOR2_X1 U612 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U613 ( .A1(G48), .A2(n776), .ZN(n555) );
  XNOR2_X1 U614 ( .A(n555), .B(KEYINPUT78), .ZN(n562) );
  NAND2_X1 U615 ( .A1(G86), .A2(n770), .ZN(n557) );
  NAND2_X1 U616 ( .A1(G61), .A2(n779), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n772), .A2(G73), .ZN(n558) );
  XOR2_X1 U619 ( .A(KEYINPUT2), .B(n558), .Z(n559) );
  NOR2_X1 U620 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n562), .A2(n561), .ZN(G305) );
  NAND2_X1 U622 ( .A1(G651), .A2(G74), .ZN(n563) );
  XOR2_X1 U623 ( .A(KEYINPUT76), .B(n563), .Z(n564) );
  NOR2_X1 U624 ( .A1(n779), .A2(n564), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n776), .A2(G49), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U627 ( .A(n567), .B(KEYINPUT77), .ZN(n570) );
  NAND2_X1 U628 ( .A1(G87), .A2(n568), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n570), .A2(n569), .ZN(G288) );
  NAND2_X1 U630 ( .A1(G85), .A2(n770), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G72), .A2(n772), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U633 ( .A1(G47), .A2(n776), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G60), .A2(n779), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n575) );
  OR2_X1 U636 ( .A1(n576), .A2(n575), .ZN(G290) );
  NAND2_X1 U637 ( .A1(G160), .A2(G40), .ZN(n696) );
  XNOR2_X1 U638 ( .A(KEYINPUT87), .B(n696), .ZN(n577) );
  NOR2_X1 U639 ( .A1(G164), .A2(G1384), .ZN(n697) );
  AND2_X2 U640 ( .A1(n577), .A2(n697), .ZN(n628) );
  XOR2_X1 U641 ( .A(KEYINPUT25), .B(G2078), .Z(n910) );
  NAND2_X1 U642 ( .A1(n628), .A2(n910), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n697), .ZN(n598) );
  INV_X1 U644 ( .A(n628), .ZN(n655) );
  NAND2_X1 U645 ( .A1(G1961), .A2(n655), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n580), .B(KEYINPUT88), .ZN(n640) );
  AND2_X1 U648 ( .A1(G301), .A2(n640), .ZN(n581) );
  XNOR2_X1 U649 ( .A(n581), .B(KEYINPUT94), .ZN(n586) );
  NOR2_X1 U650 ( .A1(G2084), .A2(n655), .ZN(n651) );
  NAND2_X1 U651 ( .A1(G8), .A2(n598), .ZN(n669) );
  NOR2_X1 U652 ( .A1(G1966), .A2(n669), .ZN(n647) );
  NOR2_X1 U653 ( .A1(n651), .A2(n647), .ZN(n582) );
  NAND2_X1 U654 ( .A1(G8), .A2(n582), .ZN(n583) );
  XNOR2_X1 U655 ( .A(KEYINPUT30), .B(n583), .ZN(n584) );
  NOR2_X1 U656 ( .A1(n584), .A2(G168), .ZN(n585) );
  NOR2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U658 ( .A(n587), .B(KEYINPUT31), .ZN(n644) );
  NAND2_X1 U659 ( .A1(n770), .A2(G81), .ZN(n588) );
  XNOR2_X1 U660 ( .A(n588), .B(KEYINPUT12), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G68), .A2(n772), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U663 ( .A(n591), .B(KEYINPUT13), .ZN(n593) );
  NAND2_X1 U664 ( .A1(G43), .A2(n776), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n779), .A2(G56), .ZN(n594) );
  NOR2_X1 U667 ( .A1(n595), .A2(n511), .ZN(n596) );
  XOR2_X1 U668 ( .A(G1996), .B(KEYINPUT91), .Z(n909) );
  XNOR2_X1 U669 ( .A(KEYINPUT26), .B(KEYINPUT92), .ZN(n612) );
  NOR2_X1 U670 ( .A1(n909), .A2(n612), .ZN(n597) );
  NOR2_X1 U671 ( .A1(n992), .A2(n597), .ZN(n609) );
  NAND2_X1 U672 ( .A1(G1348), .A2(n598), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G2067), .A2(n628), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n618) );
  NAND2_X1 U675 ( .A1(G54), .A2(n776), .ZN(n602) );
  NAND2_X1 U676 ( .A1(G66), .A2(n779), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U678 ( .A1(G92), .A2(n770), .ZN(n604) );
  NAND2_X1 U679 ( .A1(G79), .A2(n772), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U682 ( .A(n607), .B(KEYINPUT15), .ZN(n987) );
  NAND2_X1 U683 ( .A1(n618), .A2(n987), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n617) );
  INV_X1 U685 ( .A(G1341), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n610), .A2(n612), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n611), .A2(n655), .ZN(n615) );
  AND2_X1 U688 ( .A1(n628), .A2(n909), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n620) );
  NOR2_X1 U692 ( .A1(n987), .A2(n618), .ZN(n619) );
  NAND2_X1 U693 ( .A1(G53), .A2(n776), .ZN(n622) );
  NAND2_X1 U694 ( .A1(G65), .A2(n779), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U696 ( .A1(G91), .A2(n770), .ZN(n624) );
  NAND2_X1 U697 ( .A1(G78), .A2(n772), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U699 ( .A1(n626), .A2(n625), .ZN(n787) );
  NAND2_X1 U700 ( .A1(n628), .A2(G2072), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(KEYINPUT27), .ZN(n630) );
  XNOR2_X1 U702 ( .A(G1956), .B(KEYINPUT89), .ZN(n936) );
  NOR2_X1 U703 ( .A1(n936), .A2(n628), .ZN(n629) );
  NOR2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n787), .A2(n633), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n637) );
  NOR2_X1 U707 ( .A1(n787), .A2(n633), .ZN(n635) );
  XOR2_X1 U708 ( .A(KEYINPUT28), .B(KEYINPUT90), .Z(n634) );
  XNOR2_X1 U709 ( .A(n635), .B(n634), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n637), .A2(n636), .ZN(n639) );
  XOR2_X1 U711 ( .A(KEYINPUT93), .B(KEYINPUT29), .Z(n638) );
  XNOR2_X1 U712 ( .A(n639), .B(n638), .ZN(n642) );
  NOR2_X1 U713 ( .A1(n640), .A2(G301), .ZN(n641) );
  NOR2_X1 U714 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U715 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n645), .B(KEYINPUT95), .ZN(n659) );
  XNOR2_X1 U717 ( .A(n659), .B(n646), .ZN(n648) );
  NOR2_X1 U718 ( .A1(n648), .A2(n647), .ZN(n650) );
  XNOR2_X1 U719 ( .A(n650), .B(n649), .ZN(n653) );
  NAND2_X1 U720 ( .A1(G8), .A2(n651), .ZN(n652) );
  NAND2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U722 ( .A(KEYINPUT98), .B(n654), .Z(n687) );
  NOR2_X1 U723 ( .A1(G1971), .A2(n669), .ZN(n657) );
  NOR2_X1 U724 ( .A1(G2090), .A2(n655), .ZN(n656) );
  NOR2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U726 ( .A1(n658), .A2(G303), .ZN(n661) );
  NAND2_X1 U727 ( .A1(G286), .A2(n659), .ZN(n660) );
  NAND2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U729 ( .A1(G8), .A2(n662), .ZN(n663) );
  XOR2_X1 U730 ( .A(KEYINPUT32), .B(n663), .Z(n685) );
  INV_X1 U731 ( .A(n669), .ZN(n668) );
  OR2_X1 U732 ( .A1(n685), .A2(n668), .ZN(n664) );
  OR2_X2 U733 ( .A1(n687), .A2(n664), .ZN(n681) );
  NOR2_X1 U734 ( .A1(G2090), .A2(G303), .ZN(n665) );
  XNOR2_X1 U735 ( .A(n665), .B(KEYINPUT100), .ZN(n666) );
  NAND2_X1 U736 ( .A1(n666), .A2(G8), .ZN(n667) );
  NOR2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n675) );
  XOR2_X1 U738 ( .A(G1981), .B(G305), .Z(n983) );
  INV_X1 U739 ( .A(n983), .ZN(n672) );
  NOR2_X1 U740 ( .A1(G1976), .A2(G288), .ZN(n1003) );
  NAND2_X1 U741 ( .A1(n1003), .A2(KEYINPUT33), .ZN(n670) );
  NOR2_X1 U742 ( .A1(n670), .A2(n669), .ZN(n671) );
  OR2_X1 U743 ( .A1(n672), .A2(n671), .ZN(n682) );
  INV_X1 U744 ( .A(n682), .ZN(n673) );
  AND2_X1 U745 ( .A1(n673), .A2(KEYINPUT33), .ZN(n674) );
  OR2_X1 U746 ( .A1(n675), .A2(n674), .ZN(n679) );
  NOR2_X1 U747 ( .A1(G1981), .A2(G305), .ZN(n676) );
  XOR2_X1 U748 ( .A(n676), .B(KEYINPUT24), .Z(n677) );
  NOR2_X1 U749 ( .A1(n669), .A2(n677), .ZN(n678) );
  NOR2_X1 U750 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U751 ( .A1(n681), .A2(n680), .ZN(n695) );
  NOR2_X1 U752 ( .A1(n669), .A2(n682), .ZN(n683) );
  NAND2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n1001) );
  AND2_X1 U754 ( .A1(n683), .A2(n1001), .ZN(n691) );
  INV_X1 U755 ( .A(n691), .ZN(n684) );
  OR2_X1 U756 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n693) );
  NOR2_X1 U758 ( .A1(G1971), .A2(G303), .ZN(n688) );
  XOR2_X1 U759 ( .A(KEYINPUT99), .B(n688), .Z(n689) );
  OR2_X1 U760 ( .A1(n689), .A2(n1003), .ZN(n690) );
  AND2_X1 U761 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n729) );
  XNOR2_X1 U763 ( .A(G1986), .B(G290), .ZN(n1000) );
  NOR2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n740) );
  AND2_X1 U765 ( .A1(n1000), .A2(n740), .ZN(n727) );
  XNOR2_X1 U766 ( .A(G2067), .B(KEYINPUT37), .ZN(n738) );
  NAND2_X1 U767 ( .A1(n865), .A2(G140), .ZN(n698) );
  XOR2_X1 U768 ( .A(KEYINPUT83), .B(n698), .Z(n700) );
  NAND2_X1 U769 ( .A1(n866), .A2(G104), .ZN(n699) );
  NAND2_X1 U770 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U771 ( .A(KEYINPUT34), .B(n701), .ZN(n706) );
  NAND2_X1 U772 ( .A1(G128), .A2(n861), .ZN(n703) );
  NAND2_X1 U773 ( .A1(G116), .A2(n862), .ZN(n702) );
  NAND2_X1 U774 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U775 ( .A(KEYINPUT35), .B(n704), .Z(n705) );
  NOR2_X1 U776 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U777 ( .A(KEYINPUT36), .B(n707), .ZN(n884) );
  NOR2_X1 U778 ( .A1(n738), .A2(n884), .ZN(n961) );
  NAND2_X1 U779 ( .A1(n740), .A2(n961), .ZN(n736) );
  XOR2_X1 U780 ( .A(KEYINPUT84), .B(G1991), .Z(n916) );
  NAND2_X1 U781 ( .A1(G131), .A2(n865), .ZN(n709) );
  NAND2_X1 U782 ( .A1(G119), .A2(n861), .ZN(n708) );
  NAND2_X1 U783 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U784 ( .A1(G95), .A2(n866), .ZN(n711) );
  NAND2_X1 U785 ( .A1(G107), .A2(n862), .ZN(n710) );
  NAND2_X1 U786 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U787 ( .A1(n713), .A2(n712), .ZN(n873) );
  NOR2_X1 U788 ( .A1(n916), .A2(n873), .ZN(n714) );
  XOR2_X1 U789 ( .A(KEYINPUT85), .B(n714), .Z(n723) );
  NAND2_X1 U790 ( .A1(G141), .A2(n865), .ZN(n716) );
  NAND2_X1 U791 ( .A1(G129), .A2(n861), .ZN(n715) );
  NAND2_X1 U792 ( .A1(n716), .A2(n715), .ZN(n719) );
  NAND2_X1 U793 ( .A1(n866), .A2(G105), .ZN(n717) );
  XOR2_X1 U794 ( .A(KEYINPUT38), .B(n717), .Z(n718) );
  NOR2_X1 U795 ( .A1(n719), .A2(n718), .ZN(n721) );
  NAND2_X1 U796 ( .A1(n862), .A2(G117), .ZN(n720) );
  NAND2_X1 U797 ( .A1(n721), .A2(n720), .ZN(n877) );
  AND2_X1 U798 ( .A1(G1996), .A2(n877), .ZN(n722) );
  NOR2_X1 U799 ( .A1(n723), .A2(n722), .ZN(n965) );
  XOR2_X1 U800 ( .A(n740), .B(KEYINPUT86), .Z(n724) );
  NOR2_X1 U801 ( .A1(n965), .A2(n724), .ZN(n732) );
  INV_X1 U802 ( .A(n732), .ZN(n725) );
  NAND2_X1 U803 ( .A1(n736), .A2(n725), .ZN(n726) );
  OR2_X1 U804 ( .A1(n727), .A2(n726), .ZN(n728) );
  OR2_X2 U805 ( .A1(n729), .A2(n728), .ZN(n743) );
  NOR2_X1 U806 ( .A1(G1996), .A2(n877), .ZN(n968) );
  NOR2_X1 U807 ( .A1(G1986), .A2(G290), .ZN(n730) );
  AND2_X1 U808 ( .A1(n916), .A2(n873), .ZN(n960) );
  NOR2_X1 U809 ( .A1(n730), .A2(n960), .ZN(n731) );
  NOR2_X1 U810 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U811 ( .A(KEYINPUT101), .B(n733), .Z(n734) );
  NOR2_X1 U812 ( .A1(n968), .A2(n734), .ZN(n735) );
  XNOR2_X1 U813 ( .A(KEYINPUT39), .B(n735), .ZN(n737) );
  NAND2_X1 U814 ( .A1(n737), .A2(n736), .ZN(n739) );
  NAND2_X1 U815 ( .A1(n738), .A2(n884), .ZN(n979) );
  NAND2_X1 U816 ( .A1(n739), .A2(n979), .ZN(n741) );
  NAND2_X1 U817 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U818 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U819 ( .A(n744), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U820 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U821 ( .A(G860), .ZN(n753) );
  OR2_X1 U822 ( .A1(n753), .A2(n992), .ZN(G153) );
  INV_X1 U823 ( .A(G132), .ZN(G219) );
  INV_X1 U824 ( .A(n787), .ZN(G299) );
  NAND2_X1 U825 ( .A1(G7), .A2(G661), .ZN(n745) );
  XNOR2_X1 U826 ( .A(n745), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U827 ( .A(G223), .ZN(n814) );
  NAND2_X1 U828 ( .A1(n814), .A2(G567), .ZN(n746) );
  XOR2_X1 U829 ( .A(KEYINPUT11), .B(n746), .Z(G234) );
  INV_X1 U830 ( .A(G868), .ZN(n750) );
  INV_X1 U831 ( .A(n987), .ZN(n888) );
  NAND2_X1 U832 ( .A1(n750), .A2(n888), .ZN(n748) );
  NAND2_X1 U833 ( .A1(G171), .A2(G868), .ZN(n747) );
  NAND2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U835 ( .A(n749), .B(KEYINPUT69), .ZN(G284) );
  NOR2_X1 U836 ( .A1(G286), .A2(n750), .ZN(n752) );
  NOR2_X1 U837 ( .A1(G868), .A2(G299), .ZN(n751) );
  NOR2_X1 U838 ( .A1(n752), .A2(n751), .ZN(G297) );
  NAND2_X1 U839 ( .A1(n753), .A2(G559), .ZN(n754) );
  NAND2_X1 U840 ( .A1(n754), .A2(n888), .ZN(n755) );
  XNOR2_X1 U841 ( .A(n755), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U842 ( .A1(n888), .A2(G868), .ZN(n756) );
  NOR2_X1 U843 ( .A1(G559), .A2(n756), .ZN(n757) );
  XNOR2_X1 U844 ( .A(n757), .B(KEYINPUT70), .ZN(n759) );
  NOR2_X1 U845 ( .A1(n992), .A2(G868), .ZN(n758) );
  NOR2_X1 U846 ( .A1(n759), .A2(n758), .ZN(G282) );
  NAND2_X1 U847 ( .A1(G123), .A2(n861), .ZN(n760) );
  XOR2_X1 U848 ( .A(KEYINPUT71), .B(n760), .Z(n761) );
  XNOR2_X1 U849 ( .A(n761), .B(KEYINPUT18), .ZN(n763) );
  NAND2_X1 U850 ( .A1(G99), .A2(n866), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n767) );
  NAND2_X1 U852 ( .A1(G135), .A2(n865), .ZN(n765) );
  NAND2_X1 U853 ( .A1(G111), .A2(n862), .ZN(n764) );
  NAND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U855 ( .A1(n767), .A2(n766), .ZN(n959) );
  XNOR2_X1 U856 ( .A(G2096), .B(n959), .ZN(n769) );
  INV_X1 U857 ( .A(G2100), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(G156) );
  NAND2_X1 U859 ( .A1(G93), .A2(n770), .ZN(n771) );
  XNOR2_X1 U860 ( .A(n771), .B(KEYINPUT73), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G80), .A2(n772), .ZN(n773) );
  XOR2_X1 U862 ( .A(KEYINPUT74), .B(n773), .Z(n774) );
  NOR2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n776), .A2(G55), .ZN(n777) );
  NAND2_X1 U865 ( .A1(n778), .A2(n777), .ZN(n782) );
  NAND2_X1 U866 ( .A1(G67), .A2(n779), .ZN(n780) );
  XNOR2_X1 U867 ( .A(KEYINPUT75), .B(n780), .ZN(n781) );
  NOR2_X1 U868 ( .A1(n782), .A2(n781), .ZN(n791) );
  NAND2_X1 U869 ( .A1(G559), .A2(n888), .ZN(n783) );
  XNOR2_X1 U870 ( .A(n783), .B(KEYINPUT72), .ZN(n795) );
  XNOR2_X1 U871 ( .A(n992), .B(n795), .ZN(n784) );
  NOR2_X1 U872 ( .A1(G860), .A2(n784), .ZN(n785) );
  XNOR2_X1 U873 ( .A(n791), .B(n785), .ZN(G145) );
  NOR2_X1 U874 ( .A1(G868), .A2(n791), .ZN(n786) );
  XNOR2_X1 U875 ( .A(n786), .B(KEYINPUT79), .ZN(n798) );
  XNOR2_X1 U876 ( .A(n992), .B(G288), .ZN(n794) );
  XNOR2_X1 U877 ( .A(G166), .B(KEYINPUT19), .ZN(n789) );
  XNOR2_X1 U878 ( .A(G290), .B(n787), .ZN(n788) );
  XNOR2_X1 U879 ( .A(n789), .B(n788), .ZN(n790) );
  XNOR2_X1 U880 ( .A(n791), .B(n790), .ZN(n792) );
  XNOR2_X1 U881 ( .A(n792), .B(G305), .ZN(n793) );
  XNOR2_X1 U882 ( .A(n794), .B(n793), .ZN(n887) );
  XNOR2_X1 U883 ( .A(n887), .B(n795), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G868), .A2(n796), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n798), .A2(n797), .ZN(G295) );
  NAND2_X1 U886 ( .A1(G2084), .A2(G2078), .ZN(n799) );
  XOR2_X1 U887 ( .A(KEYINPUT20), .B(n799), .Z(n800) );
  NAND2_X1 U888 ( .A1(n800), .A2(G2090), .ZN(n801) );
  XNOR2_X1 U889 ( .A(n801), .B(KEYINPUT21), .ZN(n802) );
  XNOR2_X1 U890 ( .A(KEYINPUT80), .B(n802), .ZN(n803) );
  NAND2_X1 U891 ( .A1(G2072), .A2(n803), .ZN(G158) );
  XOR2_X1 U892 ( .A(KEYINPUT66), .B(G57), .Z(G237) );
  XNOR2_X1 U893 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U894 ( .A(KEYINPUT67), .B(G82), .ZN(G220) );
  NAND2_X1 U895 ( .A1(G120), .A2(G108), .ZN(n804) );
  NOR2_X1 U896 ( .A1(G237), .A2(n804), .ZN(n805) );
  NAND2_X1 U897 ( .A1(G69), .A2(n805), .ZN(n819) );
  NAND2_X1 U898 ( .A1(G567), .A2(n819), .ZN(n810) );
  NOR2_X1 U899 ( .A1(G219), .A2(G220), .ZN(n806) );
  XOR2_X1 U900 ( .A(KEYINPUT22), .B(n806), .Z(n807) );
  NOR2_X1 U901 ( .A1(G218), .A2(n807), .ZN(n808) );
  NAND2_X1 U902 ( .A1(G96), .A2(n808), .ZN(n820) );
  NAND2_X1 U903 ( .A1(G2106), .A2(n820), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U905 ( .A(KEYINPUT81), .B(n811), .ZN(G319) );
  INV_X1 U906 ( .A(G319), .ZN(n813) );
  NAND2_X1 U907 ( .A1(G661), .A2(G483), .ZN(n812) );
  NOR2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n818), .A2(G36), .ZN(G176) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n814), .ZN(G217) );
  NAND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n815) );
  XNOR2_X1 U912 ( .A(KEYINPUT103), .B(n815), .ZN(n816) );
  NAND2_X1 U913 ( .A1(n816), .A2(G661), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n817) );
  NAND2_X1 U915 ( .A1(n818), .A2(n817), .ZN(G188) );
  XOR2_X1 U916 ( .A(G108), .B(KEYINPUT114), .Z(G238) );
  INV_X1 U918 ( .A(G120), .ZN(G236) );
  INV_X1 U919 ( .A(G96), .ZN(G221) );
  INV_X1 U920 ( .A(G69), .ZN(G235) );
  NOR2_X1 U921 ( .A1(n820), .A2(n819), .ZN(G325) );
  INV_X1 U922 ( .A(G325), .ZN(G261) );
  XOR2_X1 U923 ( .A(KEYINPUT41), .B(G1971), .Z(n822) );
  XNOR2_X1 U924 ( .A(G1996), .B(G1991), .ZN(n821) );
  XNOR2_X1 U925 ( .A(n822), .B(n821), .ZN(n823) );
  XOR2_X1 U926 ( .A(n823), .B(KEYINPUT108), .Z(n825) );
  XNOR2_X1 U927 ( .A(G1966), .B(G1981), .ZN(n824) );
  XNOR2_X1 U928 ( .A(n825), .B(n824), .ZN(n829) );
  XOR2_X1 U929 ( .A(G1976), .B(G1961), .Z(n827) );
  XNOR2_X1 U930 ( .A(G1986), .B(G1956), .ZN(n826) );
  XNOR2_X1 U931 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U932 ( .A(n829), .B(n828), .Z(n831) );
  XNOR2_X1 U933 ( .A(KEYINPUT107), .B(G2474), .ZN(n830) );
  XNOR2_X1 U934 ( .A(n831), .B(n830), .ZN(G229) );
  XOR2_X1 U935 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n833) );
  XNOR2_X1 U936 ( .A(KEYINPUT104), .B(G2096), .ZN(n832) );
  XNOR2_X1 U937 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U938 ( .A(n834), .B(KEYINPUT105), .Z(n836) );
  XNOR2_X1 U939 ( .A(G2067), .B(G2072), .ZN(n835) );
  XNOR2_X1 U940 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U941 ( .A(G2100), .B(G2090), .Z(n838) );
  XNOR2_X1 U942 ( .A(G2084), .B(G2078), .ZN(n837) );
  XNOR2_X1 U943 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U944 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U945 ( .A(G2678), .B(KEYINPUT42), .ZN(n841) );
  XNOR2_X1 U946 ( .A(n842), .B(n841), .ZN(G227) );
  NAND2_X1 U947 ( .A1(n861), .A2(G124), .ZN(n843) );
  XNOR2_X1 U948 ( .A(n843), .B(KEYINPUT44), .ZN(n845) );
  NAND2_X1 U949 ( .A1(G136), .A2(n865), .ZN(n844) );
  NAND2_X1 U950 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U951 ( .A(n846), .B(KEYINPUT109), .ZN(n848) );
  NAND2_X1 U952 ( .A1(G100), .A2(n866), .ZN(n847) );
  NAND2_X1 U953 ( .A1(n848), .A2(n847), .ZN(n851) );
  NAND2_X1 U954 ( .A1(n862), .A2(G112), .ZN(n849) );
  XOR2_X1 U955 ( .A(KEYINPUT110), .B(n849), .Z(n850) );
  NOR2_X1 U956 ( .A1(n851), .A2(n850), .ZN(n852) );
  XOR2_X1 U957 ( .A(KEYINPUT111), .B(n852), .Z(G162) );
  NAND2_X1 U958 ( .A1(G139), .A2(n865), .ZN(n854) );
  NAND2_X1 U959 ( .A1(G103), .A2(n866), .ZN(n853) );
  NAND2_X1 U960 ( .A1(n854), .A2(n853), .ZN(n860) );
  NAND2_X1 U961 ( .A1(n862), .A2(G115), .ZN(n855) );
  XNOR2_X1 U962 ( .A(n855), .B(KEYINPUT112), .ZN(n857) );
  NAND2_X1 U963 ( .A1(G127), .A2(n861), .ZN(n856) );
  NAND2_X1 U964 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U965 ( .A(KEYINPUT47), .B(n858), .Z(n859) );
  NOR2_X1 U966 ( .A1(n860), .A2(n859), .ZN(n973) );
  NAND2_X1 U967 ( .A1(G130), .A2(n861), .ZN(n864) );
  NAND2_X1 U968 ( .A1(G118), .A2(n862), .ZN(n863) );
  NAND2_X1 U969 ( .A1(n864), .A2(n863), .ZN(n871) );
  NAND2_X1 U970 ( .A1(G142), .A2(n865), .ZN(n868) );
  NAND2_X1 U971 ( .A1(G106), .A2(n866), .ZN(n867) );
  NAND2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U973 ( .A(KEYINPUT45), .B(n869), .Z(n870) );
  NOR2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n973), .B(n872), .ZN(n883) );
  XNOR2_X1 U976 ( .A(G164), .B(G162), .ZN(n881) );
  XOR2_X1 U977 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n875) );
  XNOR2_X1 U978 ( .A(n873), .B(KEYINPUT46), .ZN(n874) );
  XNOR2_X1 U979 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U980 ( .A(n876), .B(n959), .Z(n879) );
  XOR2_X1 U981 ( .A(G160), .B(n877), .Z(n878) );
  XNOR2_X1 U982 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U983 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U984 ( .A(n883), .B(n882), .ZN(n885) );
  XOR2_X1 U985 ( .A(n885), .B(n884), .Z(n886) );
  NOR2_X1 U986 ( .A1(G37), .A2(n886), .ZN(G395) );
  XOR2_X1 U987 ( .A(n887), .B(G286), .Z(n890) );
  XNOR2_X1 U988 ( .A(n888), .B(G171), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U990 ( .A1(G37), .A2(n891), .ZN(G397) );
  XOR2_X1 U991 ( .A(KEYINPUT102), .B(G2446), .Z(n893) );
  XNOR2_X1 U992 ( .A(G2443), .B(G2454), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U994 ( .A(n894), .B(G2451), .Z(n896) );
  XNOR2_X1 U995 ( .A(G1341), .B(G1348), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n900) );
  XOR2_X1 U997 ( .A(G2435), .B(G2427), .Z(n898) );
  XNOR2_X1 U998 ( .A(G2430), .B(G2438), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U1000 ( .A(n900), .B(n899), .Z(n901) );
  NAND2_X1 U1001 ( .A1(G14), .A2(n901), .ZN(n907) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n907), .ZN(n904) );
  NOR2_X1 U1003 ( .A1(G229), .A2(G227), .ZN(n902) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n902), .ZN(n903) );
  NOR2_X1 U1005 ( .A1(n904), .A2(n903), .ZN(n906) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n905) );
  NAND2_X1 U1007 ( .A1(n906), .A2(n905), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(n907), .ZN(G401) );
  XOR2_X1 U1010 ( .A(G2072), .B(G33), .Z(n908) );
  NAND2_X1 U1011 ( .A1(G28), .A2(n908), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(n909), .B(G32), .ZN(n912) );
  XNOR2_X1 U1013 ( .A(n910), .B(G27), .ZN(n911) );
  NOR2_X1 U1014 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1015 ( .A(KEYINPUT118), .B(n913), .Z(n914) );
  NOR2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n920) );
  XOR2_X1 U1017 ( .A(n916), .B(G25), .Z(n918) );
  XNOR2_X1 U1018 ( .A(G2067), .B(G26), .ZN(n917) );
  NOR2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(n921), .B(KEYINPUT53), .ZN(n924) );
  XOR2_X1 U1022 ( .A(G2084), .B(G34), .Z(n922) );
  XNOR2_X1 U1023 ( .A(KEYINPUT54), .B(n922), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n927) );
  XOR2_X1 U1025 ( .A(KEYINPUT117), .B(G2090), .Z(n925) );
  XNOR2_X1 U1026 ( .A(G35), .B(n925), .ZN(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1028 ( .A(KEYINPUT119), .B(n928), .Z(n929) );
  NOR2_X1 U1029 ( .A1(G29), .A2(n929), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(KEYINPUT55), .B(n930), .ZN(n1014) );
  XOR2_X1 U1031 ( .A(G1966), .B(G21), .Z(n942) );
  XNOR2_X1 U1032 ( .A(G1348), .B(KEYINPUT59), .ZN(n931) );
  XNOR2_X1 U1033 ( .A(n931), .B(G4), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(G1341), .B(G19), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(G1981), .B(G6), .ZN(n932) );
  NOR2_X1 U1036 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n939) );
  XOR2_X1 U1038 ( .A(G20), .B(n936), .Z(n937) );
  XNOR2_X1 U1039 ( .A(KEYINPUT124), .B(n937), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1041 ( .A(n940), .B(KEYINPUT60), .ZN(n941) );
  NAND2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1043 ( .A(n943), .B(KEYINPUT125), .ZN(n951) );
  XOR2_X1 U1044 ( .A(G1986), .B(KEYINPUT126), .Z(n944) );
  XNOR2_X1 U1045 ( .A(G24), .B(n944), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(G1971), .B(G22), .ZN(n946) );
  XNOR2_X1 U1047 ( .A(G23), .B(G1976), .ZN(n945) );
  NOR2_X1 U1048 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1050 ( .A(KEYINPUT58), .B(n949), .Z(n950) );
  NAND2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1052 ( .A(G5), .B(G1961), .ZN(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1054 ( .A(n954), .B(KEYINPUT61), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(G16), .B(KEYINPUT123), .ZN(n955) );
  NAND2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n957), .ZN(n1012) );
  XOR2_X1 U1058 ( .A(G2084), .B(G160), .Z(n958) );
  NOR2_X1 U1059 ( .A1(n959), .A2(n958), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1062 ( .A(KEYINPUT115), .B(n964), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n971) );
  XOR2_X1 U1064 ( .A(G2090), .B(G162), .Z(n967) );
  NOR2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(n969), .B(KEYINPUT51), .ZN(n970) );
  NOR2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1068 ( .A(KEYINPUT116), .B(n972), .Z(n978) );
  XOR2_X1 U1069 ( .A(G2072), .B(n973), .Z(n975) );
  XOR2_X1 U1070 ( .A(G164), .B(G2078), .Z(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1072 ( .A(KEYINPUT50), .B(n976), .Z(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(n981), .B(KEYINPUT52), .ZN(n982) );
  NAND2_X1 U1076 ( .A1(n982), .A2(G29), .ZN(n1010) );
  XNOR2_X1 U1077 ( .A(G16), .B(KEYINPUT56), .ZN(n1008) );
  XNOR2_X1 U1078 ( .A(G1966), .B(G168), .ZN(n984) );
  NAND2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(n985), .B(KEYINPUT57), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(G1961), .B(KEYINPUT120), .ZN(n986) );
  XNOR2_X1 U1082 ( .A(n986), .B(G301), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(G1348), .B(n987), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(n992), .B(G1341), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n1006) );
  XNOR2_X1 U1088 ( .A(G166), .B(G1971), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(n995), .B(KEYINPUT122), .ZN(n998) );
  XNOR2_X1 U1090 ( .A(G1956), .B(KEYINPUT121), .ZN(n996) );
  XNOR2_X1 U1091 ( .A(n996), .B(G299), .ZN(n997) );
  NAND2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(n1015), .B(KEYINPUT62), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1016), .ZN(G311) );
  INV_X1 U1103 ( .A(G311), .ZN(G150) );
endmodule

