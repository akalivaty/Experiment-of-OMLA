//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G116), .B2(G270), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G58), .A2(G232), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G50), .A2(G226), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n207), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n210), .B(new_n224), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G1), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n246), .B1(G41), .B2(G45), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT65), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G41), .ZN(new_n251));
  OAI211_X1 g0051(.A(G1), .B(G13), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n246), .B(KEYINPUT65), .C1(G41), .C2(G45), .ZN(new_n253));
  AND3_X1   g0053(.A1(new_n249), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G226), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G222), .A2(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G223), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n256), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n252), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n260), .B(new_n261), .C1(G77), .C2(new_n256), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n247), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n255), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  OR3_X1    g0066(.A1(new_n266), .A2(KEYINPUT68), .A3(G179), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n225), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n246), .B2(G20), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G50), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n246), .A2(G13), .A3(G20), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G50), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n226), .B1(new_n201), .B2(new_n202), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n226), .A2(new_n250), .ZN(new_n276));
  INV_X1    g0076(.A(G150), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G58), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT67), .B1(new_n279), .B2(KEYINPUT8), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT67), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT8), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(new_n282), .A3(G58), .ZN(new_n283));
  AND3_X1   g0083(.A1(new_n279), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT66), .B1(new_n279), .B2(KEYINPUT8), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n280), .B(new_n283), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n250), .A2(G20), .ZN(new_n287));
  AOI211_X1 g0087(.A(new_n275), .B(new_n278), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n269), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n271), .B(new_n274), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G169), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n266), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT68), .B1(new_n266), .B2(G179), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n267), .A2(new_n290), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT9), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n278), .B1(new_n286), .B2(new_n287), .ZN(new_n297));
  INV_X1    g0097(.A(new_n275), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n269), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n300), .A2(KEYINPUT9), .A3(new_n271), .A4(new_n274), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n266), .A2(G200), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n266), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n296), .A2(new_n301), .A3(new_n302), .A4(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n294), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT16), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT3), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n310), .A2(KEYINPUT73), .A3(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT73), .B1(new_n310), .B2(G33), .ZN(new_n314));
  OAI211_X1 g0114(.A(KEYINPUT7), .B(new_n226), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT7), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(new_n256), .B2(G20), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n220), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n279), .A2(new_n220), .ZN(new_n319));
  OAI21_X1  g0119(.A(G20), .B1(new_n319), .B2(new_n201), .ZN(new_n320));
  NOR2_X1   g0120(.A1(G20), .A2(G33), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G159), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n309), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n310), .A2(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n312), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n317), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G68), .ZN(new_n329));
  INV_X1    g0129(.A(new_n323), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(KEYINPUT16), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n324), .A2(new_n331), .A3(new_n269), .ZN(new_n332));
  OR2_X1    g0132(.A1(G223), .A2(G1698), .ZN(new_n333));
  INV_X1    g0133(.A(G226), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G1698), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n256), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G87), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n261), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n254), .A2(G232), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n339), .A2(new_n340), .A3(G190), .A4(new_n265), .ZN(new_n341));
  INV_X1    g0141(.A(new_n272), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n286), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n270), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n343), .B1(new_n286), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n249), .A2(new_n252), .A3(new_n253), .ZN(new_n347));
  INV_X1    g0147(.A(G232), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n265), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n252), .B1(new_n336), .B2(new_n337), .ZN(new_n350));
  OAI21_X1  g0150(.A(G200), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n332), .A2(new_n341), .A3(new_n346), .A4(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT17), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n323), .B1(new_n328), .B2(G68), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n289), .B1(new_n355), .B2(KEYINPUT16), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n345), .B1(new_n356), .B2(new_n324), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n357), .A2(KEYINPUT17), .A3(new_n341), .A4(new_n351), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n332), .A2(new_n346), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n339), .A2(new_n340), .A3(G179), .A4(new_n265), .ZN(new_n361));
  OAI21_X1  g0161(.A(G169), .B1(new_n349), .B2(new_n350), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT18), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT18), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n357), .A2(new_n366), .A3(new_n363), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n308), .A2(new_n359), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n256), .A2(G238), .A3(G1698), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n256), .A2(G232), .A3(new_n258), .ZN(new_n371));
  INV_X1    g0171(.A(G107), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n370), .B(new_n371), .C1(new_n372), .C2(new_n256), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n261), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n254), .A2(G244), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n265), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT69), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n264), .B1(new_n373), .B2(new_n261), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(KEYINPUT69), .A3(new_n375), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(G200), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n279), .A2(KEYINPUT8), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n282), .A2(G58), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(new_n321), .B1(G20), .B2(G77), .ZN(new_n386));
  INV_X1    g0186(.A(new_n287), .ZN(new_n387));
  XOR2_X1   g0187(.A(KEYINPUT15), .B(G87), .Z(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n386), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G77), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n390), .A2(new_n269), .B1(new_n391), .B2(new_n342), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n270), .A2(G77), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n380), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT69), .B1(new_n379), .B2(new_n375), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n381), .B(new_n395), .C1(new_n398), .C2(new_n303), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n264), .B1(new_n254), .B2(G238), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT13), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n334), .A2(new_n258), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n348), .A2(G1698), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n256), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G97), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n261), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n400), .A2(new_n401), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n265), .B1(new_n347), .B2(new_n221), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n252), .B1(new_n404), .B2(new_n405), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT13), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G179), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT72), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT14), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n412), .A2(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n415), .ZN(new_n418));
  INV_X1    g0218(.A(new_n412), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n418), .B1(new_n419), .B2(new_n291), .ZN(new_n420));
  AOI211_X1 g0220(.A(new_n291), .B(new_n418), .C1(new_n408), .C2(new_n411), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n417), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT70), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n276), .B2(new_n202), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n220), .A2(G20), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n287), .A2(G77), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n321), .A2(KEYINPUT70), .A3(G50), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n425), .A2(new_n426), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n269), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT11), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n430), .A2(new_n431), .B1(G68), .B2(new_n270), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(KEYINPUT11), .A3(new_n269), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n342), .A2(new_n220), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(KEYINPUT71), .B2(KEYINPUT12), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(KEYINPUT71), .B2(KEYINPUT12), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n432), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n423), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n378), .A2(new_n291), .A3(new_n380), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n394), .B(new_n442), .C1(new_n398), .C2(G179), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n412), .A2(G200), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n408), .A2(G190), .A3(new_n411), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(new_n437), .A3(new_n439), .A4(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n369), .A2(new_n399), .A3(new_n445), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n312), .A2(new_n325), .A3(G257), .A4(G1698), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n312), .A2(new_n325), .A3(G250), .A4(new_n258), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G294), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT87), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT87), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n451), .A2(new_n452), .A3(new_n456), .A4(new_n453), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n261), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT5), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT78), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(G41), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n251), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n462));
  INV_X1    g0262(.A(G45), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(G1), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n461), .A2(new_n462), .A3(new_n464), .A4(G274), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n461), .A2(new_n464), .A3(new_n462), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(G264), .A3(new_n252), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n458), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n291), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n458), .A2(new_n467), .A3(new_n413), .A4(new_n465), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT86), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT24), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G116), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G20), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n312), .A2(new_n325), .A3(new_n226), .A4(G87), .ZN(new_n477));
  NAND2_X1  g0277(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n256), .A2(new_n226), .A3(G87), .A4(new_n478), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n476), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT23), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n226), .B2(G107), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n372), .A2(KEYINPUT23), .A3(G20), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI211_X1 g0287(.A(new_n473), .B(new_n474), .C1(new_n482), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n480), .A2(new_n481), .ZN(new_n489));
  INV_X1    g0289(.A(new_n476), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(new_n487), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT86), .B1(new_n491), .B2(KEYINPUT24), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n489), .A2(new_n474), .A3(new_n490), .A4(new_n487), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT85), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n482), .A2(KEYINPUT85), .A3(new_n474), .A4(new_n487), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n289), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n342), .A2(KEYINPUT25), .A3(new_n372), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT25), .B1(new_n342), .B2(new_n372), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n246), .A2(G33), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n272), .A2(new_n503), .A3(new_n225), .A4(new_n268), .ZN(new_n504));
  OAI22_X1  g0304(.A1(new_n501), .A2(new_n502), .B1(new_n372), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(KEYINPUT88), .B(new_n472), .C1(new_n499), .C2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT88), .ZN(new_n507));
  AOI211_X1 g0307(.A(new_n476), .B(new_n486), .C1(new_n480), .C2(new_n481), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n473), .B1(new_n508), .B2(new_n474), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n491), .A2(KEYINPUT86), .A3(KEYINPUT24), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n509), .A2(new_n496), .A3(new_n497), .A4(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n505), .B1(new_n511), .B2(new_n269), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n507), .B1(new_n512), .B2(new_n471), .ZN(new_n513));
  INV_X1    g0313(.A(new_n468), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G190), .ZN(new_n515));
  AOI221_X4 g0315(.A(new_n505), .B1(G200), .B2(new_n468), .C1(new_n511), .C2(new_n269), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n506), .A2(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n312), .A2(new_n325), .A3(G244), .A4(new_n258), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT4), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .A4(new_n258), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n256), .A2(G250), .A3(G1698), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n261), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n466), .A2(G257), .A3(new_n252), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n526), .A2(new_n465), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(new_n303), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n524), .A2(KEYINPUT77), .A3(new_n261), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT77), .B1(new_n524), .B2(new_n261), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n529), .B1(G200), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(G97), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n342), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n504), .B2(new_n534), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n315), .A2(new_n317), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G107), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT76), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n537), .A2(KEYINPUT76), .A3(G107), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT75), .ZN(new_n542));
  OR2_X1    g0342(.A1(KEYINPUT74), .A2(G97), .ZN(new_n543));
  NAND2_X1  g0343(.A1(KEYINPUT74), .A2(G97), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n543), .A2(KEYINPUT6), .A3(new_n372), .A4(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT6), .ZN(new_n546));
  AND2_X1   g0346(.A1(G97), .A2(G107), .ZN(new_n547));
  NOR2_X1   g0347(.A1(G97), .A2(G107), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n226), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n276), .A2(new_n391), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n542), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n545), .A2(new_n549), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n551), .B1(new_n553), .B2(G20), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT75), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n540), .A2(new_n541), .A3(new_n552), .A4(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n536), .B1(new_n556), .B2(new_n269), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n533), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n413), .B(new_n527), .C1(new_n530), .C2(new_n531), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n528), .A2(new_n291), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT76), .B1(new_n537), .B2(G107), .ZN(new_n561));
  AOI211_X1 g0361(.A(new_n539), .B(new_n372), .C1(new_n315), .C2(new_n317), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n555), .A2(new_n552), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n289), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n559), .B(new_n560), .C1(new_n565), .C2(new_n536), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n466), .A2(G270), .A3(new_n252), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n465), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n312), .A2(new_n325), .A3(G257), .A4(new_n258), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n312), .A2(new_n325), .A3(G264), .A4(G1698), .ZN(new_n571));
  INV_X1    g0371(.A(G303), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n570), .B(new_n571), .C1(new_n572), .C2(new_n256), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n261), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n291), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n504), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G116), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n272), .A2(G116), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n269), .B1(new_n226), .B2(G116), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n543), .A2(new_n250), .A3(new_n544), .ZN(new_n581));
  AOI21_X1  g0381(.A(G20), .B1(G33), .B2(G283), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT82), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT82), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n581), .A2(new_n585), .A3(new_n582), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n580), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT20), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n577), .B(new_n579), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n580), .ZN(new_n590));
  INV_X1    g0390(.A(new_n586), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n585), .B1(new_n581), .B2(new_n582), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n593), .A2(KEYINPUT20), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n575), .B1(new_n589), .B2(new_n594), .ZN(new_n595));
  XOR2_X1   g0395(.A(KEYINPUT83), .B(KEYINPUT21), .Z(new_n596));
  AND2_X1   g0396(.A1(new_n573), .A2(new_n261), .ZN(new_n597));
  OAI211_X1 g0397(.A(KEYINPUT21), .B(G169), .C1(new_n597), .C2(new_n568), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n569), .A2(G179), .A3(new_n574), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n593), .A2(KEYINPUT20), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n587), .A2(new_n588), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(new_n577), .A4(new_n579), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n595), .A2(new_n596), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n603), .ZN(new_n605));
  OAI21_X1  g0405(.A(G200), .B1(new_n597), .B2(new_n568), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n597), .A2(new_n568), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G190), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n558), .A2(new_n566), .A3(new_n604), .A4(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n388), .A2(new_n272), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n504), .A2(new_n212), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT19), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n226), .B1(new_n405), .B2(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(KEYINPUT74), .A2(G97), .ZN(new_n615));
  NOR2_X1   g0415(.A1(KEYINPUT74), .A2(G97), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n372), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(KEYINPUT80), .A2(G87), .ZN(new_n618));
  NOR2_X1   g0418(.A1(KEYINPUT80), .A2(G87), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n614), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n543), .A2(new_n544), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n613), .B1(new_n622), .B2(new_n387), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n256), .A2(new_n226), .A3(G68), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AOI211_X1 g0425(.A(new_n611), .B(new_n612), .C1(new_n625), .C2(new_n269), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n312), .A2(new_n325), .A3(G244), .A4(G1698), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT79), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT79), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n256), .A2(new_n629), .A3(G244), .A4(G1698), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n256), .A2(G238), .A3(new_n258), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n628), .A2(new_n630), .A3(new_n475), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n261), .ZN(new_n633));
  INV_X1    g0433(.A(new_n464), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n252), .A2(new_n634), .A3(G250), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n263), .B2(new_n634), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n633), .A2(G190), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(G200), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n636), .B1(new_n632), .B2(new_n261), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n626), .B(new_n638), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n633), .A2(new_n413), .A3(new_n637), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n625), .A2(new_n269), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n576), .A2(new_n388), .ZN(new_n644));
  INV_X1    g0444(.A(new_n611), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n642), .B(new_n646), .C1(G169), .C2(new_n640), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT81), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n641), .A2(new_n647), .A3(KEYINPUT81), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n610), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n450), .A2(new_n517), .A3(new_n653), .ZN(G372));
  NAND2_X1  g0454(.A1(new_n559), .A2(new_n560), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n557), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n650), .A2(new_n656), .A3(new_n651), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(KEYINPUT26), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n647), .B(KEYINPUT89), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n648), .A2(new_n557), .A3(new_n655), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n511), .A2(new_n269), .ZN(new_n664));
  INV_X1    g0464(.A(new_n505), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n468), .A2(G200), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n664), .A2(new_n665), .A3(new_n515), .A4(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n648), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(new_n566), .A4(new_n558), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n595), .A2(new_n596), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n600), .A2(new_n603), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n512), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n672), .B1(new_n673), .B2(new_n472), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n663), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n450), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n359), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n444), .A2(new_n678), .A3(new_n448), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n365), .A2(new_n367), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(KEYINPUT90), .A3(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n296), .A2(new_n301), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT10), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n302), .A4(new_n304), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT90), .B1(new_n679), .B2(new_n680), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n294), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n677), .A2(new_n689), .ZN(G369));
  NAND2_X1  g0490(.A1(new_n506), .A2(new_n513), .ZN(new_n691));
  INV_X1    g0491(.A(G13), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G20), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n246), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g0497(.A(KEYINPUT91), .B(G343), .Z(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n673), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n691), .A2(new_n667), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT94), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT94), .B1(new_n517), .B2(new_n701), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n673), .A2(new_n472), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n700), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n603), .A2(new_n700), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n672), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n604), .A2(new_n609), .A3(new_n712), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT92), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n714), .B2(new_n715), .ZN(new_n718));
  OAI21_X1  g0518(.A(G330), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT93), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n711), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT95), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n700), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n709), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n702), .A2(new_n703), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n517), .A2(KEYINPUT94), .A3(new_n701), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n604), .A2(new_n700), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n722), .A2(new_n725), .A3(new_n729), .ZN(G399));
  INV_X1    g0530(.A(new_n208), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G41), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G1), .ZN(new_n734));
  OR3_X1    g0534(.A1(new_n617), .A2(new_n620), .A3(G116), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n734), .A2(new_n735), .B1(new_n228), .B2(new_n733), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT28), .ZN(new_n737));
  INV_X1    g0537(.A(new_n700), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n669), .B1(new_n691), .B2(new_n604), .ZN(new_n739));
  INV_X1    g0539(.A(new_n659), .ZN(new_n740));
  OAI21_X1  g0540(.A(KEYINPUT26), .B1(new_n566), .B2(new_n648), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n740), .B(new_n741), .C1(new_n657), .C2(KEYINPUT26), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n738), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(KEYINPUT29), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT29), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n745), .B(new_n724), .C1(new_n663), .C2(new_n675), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n653), .A2(new_n517), .A3(new_n724), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n607), .A2(G179), .A3(new_n640), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n458), .A2(new_n525), .A3(new_n467), .A4(new_n527), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT30), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n750), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n633), .A2(new_n637), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n599), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT30), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n640), .B(KEYINPUT96), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n607), .A2(G179), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n758), .A2(new_n468), .A3(new_n532), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(KEYINPUT31), .B1(new_n761), .B2(new_n700), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT31), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n763), .B(new_n724), .C1(new_n757), .C2(new_n760), .ZN(new_n764));
  OAI21_X1  g0564(.A(KEYINPUT97), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n532), .A2(new_n759), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n640), .A2(KEYINPUT96), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n640), .A2(KEYINPUT96), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n514), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n766), .A2(new_n769), .B1(new_n751), .B2(new_n756), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n763), .B1(new_n770), .B2(new_n738), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT97), .ZN(new_n772));
  INV_X1    g0572(.A(new_n724), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n761), .A2(KEYINPUT31), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n748), .A2(new_n765), .A3(new_n775), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n776), .A2(G330), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n747), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n737), .B1(new_n778), .B2(G1), .ZN(G364));
  XNOR2_X1  g0579(.A(new_n719), .B(KEYINPUT93), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n734), .B1(G45), .B2(new_n693), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n717), .A2(new_n718), .ZN(new_n782));
  INV_X1    g0582(.A(G330), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n781), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n229), .A2(new_n463), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n731), .A2(new_n256), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n787), .B(new_n788), .C1(new_n244), .C2(new_n463), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n731), .A2(new_n326), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G355), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n789), .B(new_n791), .C1(G116), .C2(new_n208), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n225), .B1(G20), .B2(new_n291), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT98), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(KEYINPUT98), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G13), .A2(G33), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(G20), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n786), .B1(new_n792), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n226), .A2(new_n303), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n413), .A2(new_n639), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G326), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G179), .A2(G200), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n226), .B1(new_n806), .B2(G190), .ZN(new_n807));
  INV_X1    g0607(.A(G294), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n804), .A2(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT99), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  INV_X1    g0612(.A(G311), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n226), .A2(G190), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n413), .A2(G200), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n811), .B(new_n812), .C1(new_n813), .C2(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT100), .Z(new_n818));
  NAND2_X1  g0618(.A1(new_n802), .A2(new_n815), .ZN(new_n819));
  INV_X1    g0619(.A(G322), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n814), .A2(new_n806), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n256), .B1(new_n823), .B2(G329), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n803), .A2(new_n814), .ZN(new_n825));
  XOR2_X1   g0625(.A(KEYINPUT33), .B(G317), .Z(new_n826));
  OAI21_X1  g0626(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n818), .A2(new_n821), .A3(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G283), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n639), .A2(G179), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n814), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n802), .A2(new_n830), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n828), .B1(new_n829), .B2(new_n831), .C1(new_n572), .C2(new_n832), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n804), .A2(new_n202), .B1(new_n819), .B2(new_n279), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n823), .A2(G159), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n326), .B(new_n834), .C1(KEYINPUT32), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n807), .A2(new_n534), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n825), .A2(new_n220), .B1(new_n831), .B2(new_n372), .ZN(new_n838));
  INV_X1    g0638(.A(new_n816), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n837), .B(new_n838), .C1(G77), .C2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n832), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n620), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n835), .A2(KEYINPUT32), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n836), .A2(new_n840), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n833), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT101), .ZN(new_n846));
  INV_X1    g0646(.A(new_n796), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n801), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT102), .Z(new_n849));
  INV_X1    g0649(.A(new_n799), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n717), .A2(new_n718), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n785), .B1(new_n849), .B2(new_n851), .ZN(G396));
  NAND2_X1  g0652(.A1(new_n676), .A2(new_n724), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n394), .A2(new_n700), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n399), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n443), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n443), .A2(new_n700), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT106), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n443), .A2(new_n700), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n443), .B2(new_n855), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n724), .B(new_n862), .C1(new_n663), .C2(new_n675), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n859), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n853), .A2(KEYINPUT106), .A3(new_n858), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n866), .A2(new_n777), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n777), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n786), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n796), .A2(new_n797), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n819), .ZN(new_n872));
  XNOR2_X1  g0672(.A(KEYINPUT103), .B(G143), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n872), .A2(new_n873), .B1(new_n839), .B2(G159), .ZN(new_n874));
  INV_X1    g0674(.A(G137), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n874), .B1(new_n875), .B2(new_n804), .C1(new_n277), .C2(new_n825), .ZN(new_n876));
  XOR2_X1   g0676(.A(KEYINPUT104), .B(KEYINPUT34), .Z(new_n877));
  XNOR2_X1  g0677(.A(new_n876), .B(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n807), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(G58), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n326), .B1(new_n823), .B2(G132), .ZN(new_n881));
  INV_X1    g0681(.A(new_n831), .ZN(new_n882));
  AOI22_X1  g0682(.A1(G50), .A2(new_n841), .B1(new_n882), .B2(G68), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n878), .A2(new_n880), .A3(new_n881), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(G87), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n885), .B1(new_n572), .B2(new_n804), .C1(new_n813), .C2(new_n822), .ZN(new_n886));
  INV_X1    g0686(.A(new_n825), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n256), .B(new_n886), .C1(G283), .C2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(G116), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n816), .A2(new_n889), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n837), .B(new_n890), .C1(G107), .C2(new_n841), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n888), .B(new_n891), .C1(new_n808), .C2(new_n819), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  OAI221_X1 g0693(.A(new_n781), .B1(G77), .B2(new_n871), .C1(new_n893), .C2(new_n847), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT105), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n798), .B2(new_n862), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n869), .A2(new_n896), .ZN(G384));
  INV_X1    g0697(.A(new_n697), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n331), .A2(new_n269), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n355), .A2(KEYINPUT16), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n346), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n898), .B(new_n901), .C1(new_n368), .C2(new_n359), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n360), .B1(new_n364), .B2(new_n898), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT37), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(new_n904), .A3(new_n352), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n901), .B1(new_n364), .B2(new_n898), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n906), .A2(new_n352), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n905), .B1(new_n907), .B2(new_n904), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n902), .A2(new_n908), .A3(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n440), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n448), .B1(new_n914), .B2(new_n738), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n412), .A2(G169), .B1(new_n414), .B2(new_n415), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n916), .A2(new_n416), .A3(new_n421), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n915), .B1(new_n917), .B2(new_n914), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n423), .A2(new_n440), .A3(new_n738), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n856), .A2(new_n857), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n770), .A2(new_n763), .A3(new_n738), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n762), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n920), .B1(new_n748), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n913), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n360), .A2(new_n898), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n680), .B2(new_n678), .ZN(new_n927));
  INV_X1    g0727(.A(new_n905), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n904), .B1(new_n903), .B2(new_n352), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n910), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n925), .B1(new_n931), .B2(new_n912), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n924), .A2(new_n925), .B1(new_n923), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n748), .A2(new_n922), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n933), .A2(new_n450), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n924), .A2(new_n925), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n923), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(G330), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n934), .A2(G330), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n940), .A2(new_n449), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n935), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n449), .B1(new_n744), .B2(new_n746), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(new_n689), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n942), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n863), .A2(new_n857), .ZN(new_n946));
  INV_X1    g0746(.A(new_n918), .ZN(new_n947));
  INV_X1    g0747(.A(new_n919), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n946), .A2(new_n913), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n368), .A2(new_n697), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n902), .A2(new_n908), .A3(KEYINPUT38), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT38), .B1(new_n902), .B2(new_n908), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT39), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT39), .B1(new_n931), .B2(new_n912), .ZN(new_n958));
  OR3_X1    g0758(.A1(new_n957), .A2(new_n919), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT107), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n950), .A2(new_n960), .A3(new_n951), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n953), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n945), .B(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n246), .B2(new_n693), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n889), .B1(new_n553), .B2(KEYINPUT35), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n965), .B(new_n227), .C1(KEYINPUT35), .C2(new_n553), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT36), .ZN(new_n967));
  OAI21_X1  g0767(.A(G77), .B1(new_n279), .B2(new_n220), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n968), .A2(new_n228), .B1(G50), .B2(new_n220), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(G1), .A3(new_n692), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n964), .A2(new_n967), .A3(new_n970), .ZN(G367));
  OAI211_X1 g0771(.A(new_n558), .B(new_n566), .C1(new_n557), .C2(new_n724), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n656), .A2(new_n773), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n722), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n626), .A2(new_n738), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT108), .B1(new_n740), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n668), .A2(new_n977), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n668), .A2(KEYINPUT108), .A3(new_n977), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OR3_X1    g0784(.A1(new_n729), .A2(KEYINPUT42), .A3(new_n975), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n566), .B1(new_n691), .B2(new_n972), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n724), .ZN(new_n987));
  OAI21_X1  g0787(.A(KEYINPUT42), .B1(new_n729), .B2(new_n975), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n984), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n984), .A3(new_n990), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n976), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n993), .ZN(new_n995));
  INV_X1    g0795(.A(new_n976), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n995), .A2(new_n996), .A3(new_n991), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n732), .B(new_n999), .Z(new_n1000));
  NAND3_X1  g0800(.A1(new_n729), .A2(new_n725), .A3(new_n974), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT45), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n729), .A2(KEYINPUT45), .A3(new_n725), .A4(new_n974), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n729), .A2(new_n725), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT44), .B1(new_n1006), .B2(new_n975), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT44), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1008), .B(new_n974), .C1(new_n729), .C2(new_n725), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n1003), .A2(new_n1005), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n722), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n728), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n710), .B(new_n1013), .C1(new_n704), .C2(new_n705), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n729), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n780), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n721), .A2(new_n1014), .A3(new_n729), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT110), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n778), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n778), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT110), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n1004), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1023), .B(new_n722), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1012), .A2(new_n1019), .A3(new_n1021), .A4(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1000), .B1(new_n1025), .B2(new_n778), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n246), .B1(new_n693), .B2(G45), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n998), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n982), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n786), .B1(new_n1030), .B2(new_n799), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n788), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n800), .B1(new_n208), .B2(new_n389), .C1(new_n237), .C2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G159), .A2(new_n887), .B1(new_n839), .B2(G50), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n804), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n873), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1034), .B(new_n1036), .C1(new_n875), .C2(new_n822), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n819), .A2(new_n277), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n256), .B1(new_n807), .B2(new_n220), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n832), .A2(new_n279), .B1(new_n831), .B2(new_n391), .ZN(new_n1040));
  NOR4_X1   g0840(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n256), .B1(new_n823), .B2(G317), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n829), .B2(new_n816), .C1(new_n808), .C2(new_n825), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G311), .A2(new_n1035), .B1(new_n872), .B2(G303), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n832), .A2(new_n889), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1044), .B1(KEYINPUT46), .B2(new_n1045), .C1(new_n622), .C2(new_n831), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1043), .B(new_n1046), .C1(KEYINPUT46), .C2(new_n1045), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n879), .A2(G107), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1041), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT47), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1031), .B(new_n1033), .C1(new_n847), .C2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1029), .A2(new_n1051), .ZN(G387));
  NAND2_X1  g0852(.A1(new_n1021), .A2(new_n1019), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n732), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(KEYINPUT113), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n778), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT114), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT113), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1053), .A2(new_n1061), .A3(new_n732), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1055), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n841), .A2(G77), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n277), .B2(new_n822), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT112), .Z(new_n1066));
  NAND2_X1  g0866(.A1(new_n879), .A2(new_n388), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n286), .A2(new_n887), .B1(new_n882), .B2(G97), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G50), .A2(new_n872), .B1(new_n839), .B2(G68), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n326), .B(new_n1070), .C1(G159), .C2(new_n1035), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G322), .A2(new_n1035), .B1(new_n887), .B2(G311), .ZN(new_n1072));
  INV_X1    g0872(.A(G317), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1072), .B1(new_n572), .B2(new_n816), .C1(new_n1073), .C2(new_n819), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT48), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n829), .B2(new_n807), .C1(new_n808), .C2(new_n832), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT49), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n326), .B1(new_n822), .B2(new_n805), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G116), .B2(new_n882), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1071), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1080), .A2(new_n847), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n735), .A2(new_n790), .B1(new_n372), .B2(new_n731), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT111), .Z(new_n1083));
  NOR3_X1   g0883(.A1(new_n384), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n735), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(G68), .A2(G77), .ZN(new_n1086));
  OAI21_X1  g0886(.A(KEYINPUT50), .B1(new_n384), .B2(G50), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1085), .A2(new_n463), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1088), .B(new_n788), .C1(new_n234), .C2(new_n463), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1083), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1081), .B1(new_n800), .B2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1091), .B(new_n781), .C1(new_n711), .C2(new_n850), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n1027), .B2(new_n1056), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1063), .A2(new_n1094), .ZN(G393));
  NAND3_X1  g0895(.A1(new_n1012), .A2(new_n1028), .A3(new_n1024), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n832), .A2(new_n829), .B1(new_n822), .B2(new_n820), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n804), .A2(new_n1073), .B1(new_n819), .B2(new_n813), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT52), .Z(new_n1099));
  AOI211_X1 g0899(.A(new_n1097), .B(new_n1099), .C1(G116), .C2(new_n879), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n808), .B2(new_n816), .C1(new_n572), .C2(new_n825), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n256), .B(new_n1101), .C1(G107), .C2(new_n882), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n326), .B1(new_n841), .B2(G68), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n887), .A2(G50), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n823), .A2(new_n873), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1103), .A2(new_n885), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G150), .A2(new_n1035), .B1(new_n872), .B2(G159), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT51), .Z(new_n1108));
  NAND2_X1  g0908(.A1(new_n879), .A2(G77), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1106), .B(new_n1110), .C1(new_n385), .C2(new_n839), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n796), .B1(new_n1102), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n975), .A2(new_n799), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n800), .B1(new_n208), .B2(new_n622), .C1(new_n241), .C2(new_n1032), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1112), .A2(new_n781), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1096), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1012), .A2(new_n1024), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n733), .B1(new_n1117), .B2(new_n1053), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1116), .B1(new_n1118), .B2(new_n1025), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(G390));
  NOR2_X1   g0920(.A1(new_n871), .A2(new_n286), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n957), .A2(new_n958), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1121), .B1(new_n1122), .B2(new_n797), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n832), .A2(new_n277), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT53), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1125), .B(new_n256), .C1(new_n875), .C2(new_n825), .ZN(new_n1126));
  INV_X1    g0926(.A(G128), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n804), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(G125), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n822), .A2(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G50), .A2(new_n882), .B1(new_n879), .B2(G159), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n872), .A2(G132), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT54), .B(G143), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(new_n1132), .C1(new_n816), .C2(new_n1133), .ZN(new_n1134));
  NOR4_X1   g0934(.A1(new_n1126), .A2(new_n1128), .A3(new_n1130), .A4(new_n1134), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1109), .B1(new_n889), .B2(new_n819), .C1(new_n622), .C2(new_n816), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n326), .B1(new_n822), .B2(new_n808), .C1(new_n372), .C2(new_n825), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n804), .A2(new_n829), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n832), .A2(new_n212), .B1(new_n831), .B2(new_n220), .ZN(new_n1139));
  NOR4_X1   g0939(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n796), .B1(new_n1135), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1123), .A2(new_n781), .A3(new_n1141), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT115), .Z(new_n1143));
  INV_X1    g0943(.A(new_n929), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n905), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n360), .B(new_n898), .C1(new_n368), .C2(new_n359), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT38), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n919), .B1(new_n954), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n738), .B(new_n856), .C1(new_n739), .C2(new_n742), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1150), .A2(new_n857), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1149), .B1(new_n1151), .B2(new_n947), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n949), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n863), .B2(new_n857), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n1154), .A2(new_n948), .B1(new_n957), .B2(new_n958), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n923), .A2(G330), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n776), .A2(G330), .A3(new_n862), .A4(new_n949), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1152), .A2(new_n1155), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1028), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1150), .A2(new_n857), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1148), .B1(new_n1163), .B2(new_n918), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n946), .A2(new_n949), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n919), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1164), .B1(new_n1166), .B2(new_n1122), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1161), .B1(new_n1167), .B2(new_n1157), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n943), .A2(new_n689), .A3(new_n941), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n783), .B(new_n858), .C1(new_n748), .C2(new_n922), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1151), .B(new_n1160), .C1(new_n949), .C2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n946), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n776), .A2(G330), .A3(new_n862), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n1153), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1173), .B1(new_n1175), .B2(new_n1157), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1169), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1168), .A2(new_n1177), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1174), .A2(new_n1153), .B1(G330), .B2(new_n923), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1171), .B1(new_n1179), .B2(new_n1173), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1159), .A2(new_n1161), .A3(new_n1169), .A4(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1178), .A2(new_n732), .A3(new_n1181), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1143), .A2(new_n1162), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(G378));
  INV_X1    g0984(.A(KEYINPUT121), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n953), .A2(new_n1185), .A3(new_n959), .A4(new_n961), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n290), .A2(new_n898), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT55), .B1(new_n686), .B2(new_n294), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT55), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n294), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(new_n684), .C2(new_n685), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1189), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  XOR2_X1   g0994(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1195));
  NAND2_X1  g0995(.A1(new_n308), .A2(new_n1191), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n686), .A2(KEYINPUT55), .A3(new_n294), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n1188), .A3(new_n1197), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1194), .A2(new_n1195), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1195), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AND4_X1   g1001(.A1(G330), .A2(new_n936), .A3(new_n1201), .A4(new_n937), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1201), .B1(new_n933), .B2(G330), .ZN(new_n1203));
  OAI21_X1  g1003(.A(KEYINPUT120), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1187), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1201), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n938), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n933), .A2(G330), .A3(new_n1201), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(KEYINPUT121), .B1(new_n1209), .B2(new_n962), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(new_n1186), .A3(KEYINPUT120), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1205), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1028), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n1127), .A2(new_n819), .B1(new_n832), .B2(new_n1133), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT116), .Z(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n1129), .B2(new_n804), .C1(new_n277), .C2(new_n807), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G132), .B2(new_n887), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n875), .B2(new_n816), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1218), .B(new_n1219), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G33), .B(new_n1220), .C1(G159), .C2(new_n882), .ZN(new_n1221));
  AOI21_X1  g1021(.A(G41), .B1(new_n823), .B2(G124), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n251), .B1(new_n310), .B2(new_n250), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1221), .A2(new_n1222), .B1(new_n202), .B2(new_n1223), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1064), .B1(new_n822), .B2(new_n829), .C1(new_n889), .C2(new_n804), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n256), .B(new_n1225), .C1(G68), .C2(new_n879), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n389), .A2(new_n816), .B1(new_n534), .B2(new_n825), .ZN(new_n1227));
  AOI211_X1 g1027(.A(G41), .B(new_n1227), .C1(G58), .C2(new_n882), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(new_n372), .C2(new_n819), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT58), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1224), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n796), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1206), .A2(new_n797), .B1(new_n202), .B2(new_n870), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1233), .A3(new_n781), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT119), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1213), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT57), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n953), .A2(new_n961), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1238), .A2(new_n959), .A3(new_n1208), .A4(new_n1207), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1209), .A2(new_n962), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1237), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1181), .A2(KEYINPUT122), .A3(new_n1169), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT122), .B1(new_n1181), .B2(new_n1169), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1241), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n732), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1169), .B1(new_n1168), .B2(new_n1177), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT122), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1181), .A2(KEYINPUT122), .A3(new_n1169), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT57), .B1(new_n1250), .B2(new_n1212), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1236), .B1(new_n1245), .B2(new_n1251), .ZN(G375));
  INV_X1    g1052(.A(new_n1180), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1169), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1000), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n1256), .A3(new_n1177), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n949), .A2(new_n798), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n889), .A2(new_n825), .B1(new_n819), .B2(new_n829), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1067), .B1(new_n808), .B2(new_n804), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1259), .B(new_n1260), .C1(G107), .C2(new_n839), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n823), .A2(G303), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n326), .B1(new_n831), .B2(new_n391), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1263), .B(KEYINPUT123), .Z(new_n1264));
  NAND2_X1  g1064(.A1(new_n841), .A2(G97), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1261), .A2(new_n1262), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n825), .A2(new_n1133), .B1(new_n822), .B2(new_n1127), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n326), .B(new_n1267), .C1(G150), .C2(new_n839), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1035), .A2(G132), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n879), .A2(G50), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n819), .A2(new_n875), .B1(new_n831), .B2(new_n279), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(G159), .B2(new_n841), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .A4(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n847), .B1(new_n1266), .B2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n871), .A2(G68), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(new_n1258), .A2(new_n786), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1180), .B2(new_n1028), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1257), .A2(new_n1277), .ZN(G381));
  OAI211_X1 g1078(.A(new_n1236), .B(new_n1183), .C1(new_n1245), .C2(new_n1251), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1061), .B1(new_n1053), .B2(new_n732), .ZN(new_n1281));
  AOI211_X1 g1081(.A(KEYINPUT113), .B(new_n733), .C1(new_n1021), .C2(new_n1019), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1281), .A2(new_n1282), .A3(new_n1059), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1283), .A2(G396), .A3(new_n1093), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1029), .A2(new_n1051), .A3(new_n1119), .ZN(new_n1286));
  OR4_X1    g1086(.A1(G384), .A2(new_n1285), .A3(G381), .A4(new_n1286), .ZN(G407));
  OAI211_X1 g1087(.A(G407), .B(G213), .C1(new_n698), .C2(new_n1279), .ZN(G409));
  NAND3_X1  g1088(.A1(new_n1250), .A2(new_n1256), .A3(new_n1212), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1290));
  OAI211_X1 g1090(.A(KEYINPUT124), .B(new_n1234), .C1(new_n1290), .C2(new_n1027), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT124), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1027), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1234), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1292), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1289), .A2(new_n1291), .A3(new_n1183), .A4(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n699), .A2(G213), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G375), .A2(G378), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT60), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1255), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1253), .A2(KEYINPUT60), .A3(new_n1254), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1301), .A2(new_n732), .A3(new_n1177), .A4(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(G384), .A3(new_n1277), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G384), .B1(new_n1303), .B2(new_n1277), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1298), .A2(new_n1299), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1297), .ZN(new_n1309));
  OAI211_X1 g1109(.A(G2897), .B(new_n1309), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1306), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1309), .A2(G2897), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1311), .A2(new_n1304), .A3(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1310), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1314), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT63), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1308), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT126), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1318), .B1(new_n1308), .B2(new_n1316), .ZN(new_n1319));
  INV_X1    g1119(.A(G396), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1320), .B1(new_n1063), .B2(new_n1094), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1284), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT125), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1286), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1119), .B1(new_n1029), .B2(new_n1051), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1322), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(G396), .B1(new_n1283), .B2(new_n1093), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1063), .A2(new_n1320), .A3(new_n1094), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G387), .A2(G390), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1329), .A2(new_n1330), .A3(new_n1323), .A4(new_n1286), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1326), .A2(new_n1331), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1332), .A2(KEYINPUT61), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1212), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1237), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n733), .B1(new_n1250), .B2(new_n1241), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1183), .B1(new_n1337), .B2(new_n1236), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1340), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(new_n1307), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1317), .A2(new_n1319), .A3(new_n1333), .A4(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT62), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1340), .A2(new_n1344), .A3(new_n1307), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1213), .A2(new_n1235), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1346), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1347));
  OAI211_X1 g1147(.A(new_n1297), .B(new_n1296), .C1(new_n1347), .C2(new_n1183), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1310), .A2(new_n1313), .ZN(new_n1349));
  AOI21_X1  g1149(.A(KEYINPUT61), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1343), .A2(new_n1345), .A3(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(new_n1332), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1342), .A2(new_n1352), .ZN(G405));
  INV_X1    g1153(.A(new_n1307), .ZN(new_n1354));
  OAI21_X1  g1154(.A(KEYINPUT127), .B1(new_n1280), .B2(new_n1338), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT127), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1299), .A2(new_n1356), .A3(new_n1279), .ZN(new_n1357));
  AND3_X1   g1157(.A1(new_n1355), .A2(new_n1332), .A3(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1332), .B1(new_n1355), .B2(new_n1357), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1354), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1332), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1357), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1356), .B1(new_n1299), .B2(new_n1279), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1361), .B1(new_n1362), .B2(new_n1363), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1355), .A2(new_n1332), .A3(new_n1357), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1364), .A2(new_n1307), .A3(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1360), .A2(new_n1366), .ZN(G402));
endmodule


