//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n549, new_n551, new_n552, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n588,
    new_n591, new_n592, new_n594, new_n595, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT66), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  OR4_X1    g028(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n461), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n461), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(G160));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  OR2_X1    g047(.A1(G100), .A2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI221_X1 g050(.A(new_n475), .B1(new_n474), .B2(new_n473), .C1(G112), .C2(new_n461), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n476), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(G102), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n466), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(G126), .B1(new_n462), .B2(new_n463), .ZN(new_n489));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n488), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n477), .A2(new_n495), .A3(G138), .A4(new_n461), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT68), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n492), .A2(new_n500), .A3(new_n497), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n504), .A2(new_n506), .A3(new_n511), .A4(new_n513), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n510), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND3_X1  g096(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n515), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT69), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n507), .A2(new_n514), .A3(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND2_X1  g105(.A1(new_n507), .A2(G64), .ZN(new_n531));
  INV_X1    g106(.A(G77), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n532), .B2(new_n503), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G651), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n515), .A2(new_n536), .B1(new_n537), .B2(new_n518), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n535), .A2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n515), .A2(new_n541), .B1(new_n542), .B2(new_n518), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT70), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n509), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  NAND3_X1  g128(.A1(new_n514), .A2(G53), .A3(G543), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT9), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n509), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n507), .A2(new_n514), .A3(G91), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(G299));
  AND2_X1   g134(.A1(new_n514), .A2(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G49), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n507), .A2(new_n514), .A3(G87), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(G288));
  NAND4_X1  g139(.A1(new_n511), .A2(new_n513), .A3(G48), .A4(G543), .ZN(new_n565));
  INV_X1    g140(.A(G86), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n518), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n504), .A2(new_n506), .A3(G61), .ZN(new_n568));
  NAND2_X1  g143(.A1(G73), .A2(G543), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n509), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G305));
  NAND2_X1  g147(.A1(new_n560), .A2(G47), .ZN(new_n573));
  INV_X1    g148(.A(G85), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  OAI221_X1 g150(.A(new_n573), .B1(new_n574), .B2(new_n518), .C1(new_n509), .C2(new_n575), .ZN(G290));
  INV_X1    g151(.A(G92), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n518), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT10), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n560), .A2(G54), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n509), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n585), .B1(G171), .B2(new_n584), .ZN(G321));
  XNOR2_X1  g161(.A(G321), .B(KEYINPUT71), .ZN(G284));
  NAND2_X1  g162(.A1(G299), .A2(new_n584), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n588), .B1(G168), .B2(new_n584), .ZN(G297));
  OAI21_X1  g164(.A(new_n588), .B1(G168), .B2(new_n584), .ZN(G280));
  INV_X1    g165(.A(new_n583), .ZN(new_n591));
  INV_X1    g166(.A(G559), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(G860), .ZN(G148));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G868), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g171(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g172(.A(new_n466), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n477), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g174(.A(KEYINPUT72), .B(KEYINPUT12), .Z(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT13), .ZN(new_n602));
  XNOR2_X1  g177(.A(KEYINPUT73), .B(G2100), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(KEYINPUT74), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n603), .A2(KEYINPUT74), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n483), .A2(G135), .ZN(new_n607));
  NOR2_X1   g182(.A1(G99), .A2(G2105), .ZN(new_n608));
  OAI21_X1  g183(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n609));
  INV_X1    g184(.A(G123), .ZN(new_n610));
  OAI221_X1 g185(.A(new_n607), .B1(new_n608), .B2(new_n609), .C1(new_n610), .C2(new_n478), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(G2096), .Z(new_n612));
  OAI211_X1 g187(.A(new_n606), .B(new_n612), .C1(new_n604), .C2(new_n602), .ZN(G156));
  XNOR2_X1  g188(.A(KEYINPUT15), .B(G2430), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2435), .ZN(new_n615));
  XOR2_X1   g190(.A(G2427), .B(G2438), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT14), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2443), .ZN(new_n619));
  XOR2_X1   g194(.A(G1341), .B(G1348), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2446), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT16), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n619), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2451), .B(G2454), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT75), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n623), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G14), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT76), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(G401));
  XOR2_X1   g204(.A(G2084), .B(G2090), .Z(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2067), .B(G2678), .Z(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT17), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT18), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2072), .B(G2078), .Z(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(new_n633), .B2(KEYINPUT18), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2096), .B(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(G227));
  XNOR2_X1  g217(.A(G1971), .B(G1976), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT19), .ZN(new_n644));
  XOR2_X1   g219(.A(G1956), .B(G2474), .Z(new_n645));
  XOR2_X1   g220(.A(G1961), .B(G1966), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n644), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n645), .A2(new_n646), .ZN(new_n650));
  AOI22_X1  g225(.A1(new_n648), .A2(KEYINPUT20), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n652), .A2(new_n644), .A3(new_n647), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n651), .B(new_n653), .C1(KEYINPUT20), .C2(new_n648), .ZN(new_n654));
  XOR2_X1   g229(.A(G1991), .B(G1996), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT78), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G1981), .B(G1986), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT77), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n659), .B(new_n661), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G229));
  INV_X1    g238(.A(G29), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(G35), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(G162), .B2(new_n664), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT29), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n479), .A2(G129), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n598), .A2(G105), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n483), .A2(G141), .ZN(new_n671));
  NAND3_X1  g246(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT26), .Z(new_n673));
  NAND4_X1  g248(.A1(new_n669), .A2(new_n670), .A3(new_n671), .A4(new_n673), .ZN(new_n674));
  MUX2_X1   g249(.A(G32), .B(new_n674), .S(G29), .Z(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT86), .Z(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT27), .B(G1996), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT87), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n598), .A2(G103), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT25), .Z(new_n681));
  NAND2_X1  g256(.A1(new_n483), .A2(G139), .ZN(new_n682));
  AOI22_X1  g257(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n681), .B(new_n682), .C1(new_n461), .C2(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(G33), .B(new_n684), .S(G29), .Z(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(G2072), .Z(new_n686));
  AND2_X1   g261(.A1(KEYINPUT24), .A2(G34), .ZN(new_n687));
  NOR2_X1   g262(.A1(KEYINPUT24), .A2(G34), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n687), .A2(new_n688), .A3(G29), .ZN(new_n689));
  INV_X1    g264(.A(G160), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(G29), .ZN(new_n691));
  INV_X1    g266(.A(G2084), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT85), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n679), .A2(new_n686), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT88), .ZN(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n547), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n697), .B2(G19), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT82), .B(G1341), .Z(new_n700));
  OAI22_X1  g275(.A1(new_n699), .A2(new_n700), .B1(new_n677), .B2(new_n676), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n591), .A2(new_n697), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G4), .B2(new_n697), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT81), .B(G1348), .Z(new_n705));
  OAI21_X1  g280(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AOI211_X1 g281(.A(new_n701), .B(new_n706), .C1(new_n705), .C2(new_n704), .ZN(new_n707));
  NAND2_X1  g282(.A1(G299), .A2(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(KEYINPUT23), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n697), .A2(G20), .ZN(new_n710));
  MUX2_X1   g285(.A(KEYINPUT23), .B(new_n709), .S(new_n710), .Z(new_n711));
  AND2_X1   g286(.A1(new_n711), .A2(G1956), .ZN(new_n712));
  NOR2_X1   g287(.A1(G168), .A2(new_n697), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n697), .B2(G21), .ZN(new_n714));
  INV_X1    g289(.A(G1966), .ZN(new_n715));
  OAI22_X1  g290(.A1(new_n714), .A2(new_n715), .B1(G1956), .B2(new_n711), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n712), .B(new_n716), .C1(new_n715), .C2(new_n714), .ZN(new_n717));
  NOR2_X1   g292(.A1(G27), .A2(G29), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G164), .B2(G29), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(G2078), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT31), .B(G11), .ZN(new_n721));
  OAI21_X1  g296(.A(KEYINPUT89), .B1(G5), .B2(G16), .ZN(new_n722));
  OR3_X1    g297(.A1(KEYINPUT89), .A2(G5), .A3(G16), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n722), .B(new_n723), .C1(G301), .C2(new_n697), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1961), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n479), .A2(G128), .B1(G140), .B2(new_n483), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n461), .A2(G116), .ZN(new_n727));
  OR3_X1    g302(.A1(KEYINPUT83), .A2(G104), .A3(G2105), .ZN(new_n728));
  OAI21_X1  g303(.A(KEYINPUT83), .B1(G104), .B2(G2105), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n728), .A2(G2104), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n726), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n664), .A2(G26), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT84), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT28), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G2067), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G28), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n739), .B2(KEYINPUT30), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(KEYINPUT30), .B2(new_n739), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n611), .B2(new_n664), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n691), .B2(new_n692), .ZN(new_n743));
  AND4_X1   g318(.A1(new_n721), .A2(new_n725), .A3(new_n738), .A4(new_n743), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n707), .A2(new_n717), .A3(new_n720), .A4(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n696), .A2(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G24), .B(G290), .S(G16), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G1986), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n483), .A2(G131), .ZN(new_n749));
  NOR2_X1   g324(.A1(G95), .A2(G2105), .ZN(new_n750));
  OAI21_X1  g325(.A(G2104), .B1(new_n461), .B2(G107), .ZN(new_n751));
  INV_X1    g326(.A(G119), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n749), .B1(new_n750), .B2(new_n751), .C1(new_n752), .C2(new_n478), .ZN(new_n753));
  MUX2_X1   g328(.A(G25), .B(new_n753), .S(G29), .Z(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT79), .Z(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT35), .B(G1991), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n747), .A2(G1986), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n697), .A2(G22), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G166), .B2(new_n697), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1971), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n697), .A2(G23), .ZN(new_n764));
  INV_X1    g339(.A(G288), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(new_n697), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT33), .Z(new_n767));
  AOI21_X1  g342(.A(new_n763), .B1(G1976), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n697), .A2(G6), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n571), .B2(new_n697), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT32), .B(G1981), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n768), .B(new_n772), .C1(G1976), .C2(new_n767), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n748), .B(new_n760), .C1(new_n773), .C2(KEYINPUT34), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT80), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT36), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n773), .A2(KEYINPUT34), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n777), .B1(new_n776), .B2(new_n778), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n668), .B(new_n746), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(G311));
  NAND2_X1  g358(.A1(new_n782), .A2(KEYINPUT90), .ZN(new_n784));
  INV_X1    g359(.A(new_n781), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(new_n779), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT90), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n786), .A2(new_n787), .A3(new_n668), .A4(new_n746), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n784), .A2(new_n788), .ZN(G150));
  AOI22_X1  g364(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(new_n509), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT91), .B(G55), .Z(new_n792));
  INV_X1    g367(.A(G93), .ZN(new_n793));
  OAI22_X1  g368(.A1(new_n515), .A2(new_n792), .B1(new_n793), .B2(new_n518), .ZN(new_n794));
  OAI21_X1  g369(.A(G860), .B1(new_n791), .B2(new_n794), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT37), .Z(new_n796));
  INV_X1    g371(.A(KEYINPUT92), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n544), .A2(new_n797), .A3(new_n546), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n791), .A2(new_n794), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n797), .B1(new_n544), .B2(new_n546), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n547), .A2(new_n797), .A3(new_n799), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n583), .A2(new_n592), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n804), .B(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n796), .B1(new_n808), .B2(G860), .ZN(G145));
  XNOR2_X1  g384(.A(new_n485), .B(new_n690), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(new_n611), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n674), .B(new_n498), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(new_n731), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(new_n684), .ZN(new_n814));
  INV_X1    g389(.A(G130), .ZN(new_n815));
  NOR2_X1   g390(.A1(G106), .A2(G2105), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n478), .A2(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G142), .B2(new_n483), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(new_n753), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(new_n601), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n814), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n822), .A2(KEYINPUT93), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n814), .A2(new_n821), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n822), .B2(KEYINPUT93), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n811), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(G37), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n822), .A2(new_n811), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n828), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g406(.A(G290), .B(G288), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT95), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(G303), .B(new_n571), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n832), .A2(new_n833), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n832), .A2(new_n835), .A3(new_n833), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(KEYINPUT96), .A2(KEYINPUT42), .ZN(new_n842));
  NAND2_X1  g417(.A1(KEYINPUT96), .A2(KEYINPUT42), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n843), .B2(new_n841), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n804), .B(new_n594), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n583), .A2(new_n557), .A3(new_n558), .A4(new_n555), .ZN(new_n848));
  NAND4_X1  g423(.A1(G299), .A2(new_n580), .A3(new_n579), .A4(new_n582), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n848), .A2(KEYINPUT41), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT41), .B1(new_n848), .B2(new_n849), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n847), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n847), .B2(new_n850), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n848), .A2(new_n849), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n857), .B2(new_n846), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n845), .B(new_n858), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G868), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(G868), .B2(new_n799), .ZN(G331));
  XNOR2_X1  g436(.A(G331), .B(KEYINPUT97), .ZN(G295));
  NAND4_X1  g437(.A1(G301), .A2(new_n525), .A3(new_n526), .A4(new_n528), .ZN(new_n863));
  NAND2_X1  g438(.A1(G171), .A2(G286), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n863), .B(new_n864), .C1(new_n802), .C2(new_n803), .ZN(new_n865));
  INV_X1    g440(.A(new_n801), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n866), .A2(new_n799), .A3(new_n798), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n863), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n800), .A2(new_n801), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n865), .A2(new_n870), .A3(KEYINPUT98), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n804), .A2(new_n872), .A3(new_n868), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n853), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT99), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n865), .A2(new_n870), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n804), .A2(KEYINPUT100), .A3(new_n868), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n857), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n871), .A2(new_n853), .A3(new_n881), .A4(new_n873), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n875), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n840), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT101), .B1(new_n884), .B2(new_n827), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n886));
  AOI211_X1 g461(.A(new_n886), .B(G37), .C1(new_n883), .C2(new_n840), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n883), .A2(new_n840), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT43), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n850), .A2(new_n851), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n879), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n856), .B1(new_n871), .B2(new_n873), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n840), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AND4_X1   g469(.A1(KEYINPUT43), .A2(new_n889), .A3(new_n827), .A4(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT44), .B1(new_n890), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(new_n888), .B2(new_n889), .ZN(new_n899));
  AND4_X1   g474(.A1(new_n898), .A2(new_n889), .A3(new_n827), .A4(new_n894), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n896), .A2(new_n901), .ZN(G397));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n903));
  NAND3_X1  g478(.A1(G160), .A2(new_n903), .A3(G40), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n483), .A2(G137), .B1(G101), .B2(new_n598), .ZN(new_n905));
  INV_X1    g480(.A(G125), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(new_n481), .B2(new_n482), .ZN(new_n907));
  INV_X1    g482(.A(new_n469), .ZN(new_n908));
  OAI21_X1  g483(.A(G2105), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n909), .A3(G40), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT103), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(KEYINPUT102), .B(G1384), .Z(new_n913));
  AOI21_X1  g488(.A(KEYINPUT45), .B1(new_n498), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n731), .B(G2067), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT104), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n753), .A2(new_n756), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n753), .A2(new_n756), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n674), .B(G1996), .ZN(new_n921));
  NOR4_X1   g496(.A1(new_n918), .A2(new_n919), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(G290), .B(G1986), .Z(new_n923));
  AOI21_X1  g498(.A(new_n915), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(KEYINPUT120), .B(KEYINPUT51), .Z(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G8), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n492), .A2(new_n500), .A3(new_n497), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n500), .B1(new_n492), .B2(new_n497), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n928), .A2(new_n929), .A3(G1384), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT50), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT105), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G1384), .B1(new_n492), .B2(new_n497), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n911), .A2(new_n904), .B1(new_n933), .B2(new_n931), .ZN(new_n934));
  INV_X1    g509(.A(G1384), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n499), .A2(new_n935), .A3(new_n501), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT50), .ZN(new_n938));
  XOR2_X1   g513(.A(KEYINPUT113), .B(G2084), .Z(new_n939));
  NAND4_X1  g514(.A1(new_n932), .A2(new_n934), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n933), .A2(KEYINPUT45), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n912), .B(new_n941), .C1(new_n936), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n715), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n927), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(KEYINPUT107), .B(G8), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(G168), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n926), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT121), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI211_X1 g526(.A(KEYINPUT121), .B(new_n926), .C1(new_n945), .C2(new_n948), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n947), .B1(new_n940), .B2(new_n944), .ZN(new_n953));
  OAI22_X1  g528(.A1(new_n953), .A2(KEYINPUT122), .B1(G168), .B2(new_n947), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n940), .A2(new_n944), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n946), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT122), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n951), .B(new_n952), .C1(new_n954), .C2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT62), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n956), .A2(new_n948), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n961), .B1(new_n960), .B2(new_n962), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n947), .B1(new_n912), .B2(new_n933), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n966));
  INV_X1    g541(.A(G1976), .ZN(new_n967));
  NAND2_X1  g542(.A1(G288), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n765), .A2(G1976), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n965), .A2(new_n966), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n966), .B1(new_n965), .B2(new_n969), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1981), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT109), .B1(new_n571), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  NOR4_X1   g551(.A1(new_n567), .A2(new_n570), .A3(new_n976), .A4(G1981), .ZN(new_n977));
  OAI22_X1  g552(.A1(new_n975), .A2(new_n977), .B1(new_n974), .B2(new_n571), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT49), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI221_X1 g555(.A(KEYINPUT49), .B1(new_n974), .B2(new_n571), .C1(new_n975), .C2(new_n977), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n965), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n903), .B1(G160), .B2(G40), .ZN(new_n983));
  AND4_X1   g558(.A1(new_n903), .A2(new_n905), .A3(new_n909), .A4(G40), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n933), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(new_n969), .A3(new_n946), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n987), .A2(KEYINPUT108), .A3(new_n966), .A4(new_n968), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n973), .A2(new_n982), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n936), .A2(new_n942), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n913), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n912), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1971), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G2090), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n932), .A2(new_n995), .A3(new_n934), .A4(new_n938), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n927), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(G303), .A2(G8), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT106), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT106), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1000), .A2(new_n1004), .A3(new_n1001), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n989), .B1(new_n997), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n912), .B1(new_n931), .B2(new_n933), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT111), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n930), .A2(new_n931), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n912), .B(new_n1011), .C1(new_n931), .C2(new_n933), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1009), .A2(new_n995), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n947), .B1(new_n1013), .B2(new_n994), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1002), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(KEYINPUT112), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n1014), .B2(new_n1002), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1007), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n992), .A2(G2078), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1022));
  INV_X1    g597(.A(G1961), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n932), .A2(new_n934), .A3(new_n938), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1021), .A2(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(G2078), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1025), .B1(new_n1027), .B2(new_n943), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1020), .A2(G171), .A3(new_n1028), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n963), .A2(new_n964), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n972), .B1(new_n986), .B2(KEYINPUT52), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n985), .A2(new_n969), .A3(new_n966), .A4(new_n946), .ZN(new_n1032));
  INV_X1    g607(.A(new_n968), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n982), .B1(new_n970), .B2(new_n972), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT110), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n973), .A2(new_n1038), .A3(new_n988), .A4(new_n982), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(new_n997), .A3(new_n1006), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n982), .A2(new_n967), .A3(new_n765), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(new_n975), .B2(new_n977), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1043), .A2(new_n965), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT63), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n997), .B2(new_n1006), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n994), .A2(new_n996), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1002), .B1(new_n1048), .B2(G8), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n953), .A2(G168), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1040), .A2(new_n1047), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1048), .A2(G8), .A3(new_n1006), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1037), .A2(new_n1054), .A3(KEYINPUT63), .A4(new_n1039), .ZN(new_n1055));
  OAI211_X1 g630(.A(G168), .B(new_n953), .C1(new_n997), .C2(new_n1002), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT114), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1050), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1007), .A2(new_n1017), .A3(new_n1019), .A4(new_n1059), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1060), .A2(new_n1046), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1041), .B(new_n1045), .C1(new_n1058), .C2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1030), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1024), .A2(new_n705), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n912), .A2(new_n737), .A3(new_n933), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1066), .ZN(new_n1068));
  AOI211_X1 g643(.A(KEYINPUT116), .B(new_n1068), .C1(new_n1024), .C2(new_n705), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT60), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT119), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1072), .B(KEYINPUT60), .C1(new_n1067), .C2(new_n1069), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(new_n591), .A3(new_n1073), .ZN(new_n1074));
  OR3_X1    g649(.A1(new_n1067), .A2(new_n1069), .A3(KEYINPUT60), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1070), .A2(KEYINPUT119), .A3(new_n583), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1078));
  INV_X1    g653(.A(G1956), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(G299), .B(KEYINPUT57), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT56), .B(G2072), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n990), .A2(new_n912), .A3(new_n991), .A4(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1080), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT115), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n1081), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1080), .A2(new_n1089), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1086), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT61), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1088), .A2(KEYINPUT61), .A3(new_n1085), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT58), .B(G1341), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n985), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n992), .B2(G1996), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(KEYINPUT117), .B(new_n1096), .C1(new_n992), .C2(G1996), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1099), .A2(new_n547), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1101), .A2(KEYINPUT118), .A3(KEYINPUT59), .ZN(new_n1102));
  NAND2_X1  g677(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1099), .A2(new_n547), .A3(new_n1103), .A4(new_n1100), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1093), .A2(new_n1094), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1077), .A2(new_n1106), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1067), .A2(new_n1069), .A3(new_n583), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1088), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1086), .B(new_n1090), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(G301), .B(KEYINPUT54), .ZN(new_n1112));
  INV_X1    g687(.A(new_n991), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1113), .A2(new_n1027), .A3(new_n914), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n910), .B(KEYINPUT124), .Z(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1025), .A2(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1020), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1028), .A2(new_n1112), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n960), .A2(new_n962), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1111), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n924), .B1(new_n1063), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n915), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n918), .B2(new_n674), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT46), .ZN(new_n1127));
  OR3_X1    g702(.A1(new_n915), .A2(new_n1127), .A3(G1996), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(new_n915), .B2(G1996), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT47), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n915), .A2(G1986), .A3(G290), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1132), .B(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n922), .B2(new_n915), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n918), .A2(new_n921), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n919), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(G2067), .B2(new_n731), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1125), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1131), .A2(new_n1135), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT126), .B1(new_n1124), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1140), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1053), .A2(new_n1057), .B1(new_n1060), .B2(new_n1046), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(new_n1044), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1120), .A2(KEYINPUT62), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1041), .B(new_n1145), .C1(new_n1148), .C2(new_n1029), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1121), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1142), .B(new_n1143), .C1(new_n1151), .C2(new_n924), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1141), .A2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g728(.A1(new_n884), .A2(new_n827), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n1155), .A2(new_n886), .ZN(new_n1156));
  NAND3_X1  g730(.A1(new_n884), .A2(KEYINPUT101), .A3(new_n827), .ZN(new_n1157));
  NAND3_X1  g731(.A1(new_n1156), .A2(new_n889), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g732(.A(new_n900), .B1(new_n1158), .B2(KEYINPUT43), .ZN(new_n1159));
  NOR2_X1   g733(.A1(G227), .A2(new_n459), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n628), .A2(new_n662), .A3(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g735(.A(new_n1161), .B(KEYINPUT127), .ZN(new_n1162));
  NOR3_X1   g736(.A1(new_n1159), .A2(new_n1162), .A3(new_n830), .ZN(G308));
  OR3_X1    g737(.A1(new_n1159), .A2(new_n1162), .A3(new_n830), .ZN(G225));
endmodule


