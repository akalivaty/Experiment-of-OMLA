

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U557 ( .A1(n676), .A2(n668), .ZN(n669) );
  NOR2_X1 U558 ( .A1(n657), .A2(n939), .ZN(n676) );
  INV_X1 U559 ( .A(KEYINPUT31), .ZN(n696) );
  INV_X1 U560 ( .A(n644), .ZN(n700) );
  NOR2_X2 U561 ( .A1(n597), .A2(n528), .ZN(n786) );
  NOR2_X2 U562 ( .A1(G2105), .A2(n537), .ZN(n990) );
  NOR2_X1 U563 ( .A1(G651), .A2(n597), .ZN(n790) );
  AND2_X1 U564 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U565 ( .A(G543), .B(KEYINPUT0), .ZN(n524) );
  XNOR2_X1 U566 ( .A(n524), .B(KEYINPUT69), .ZN(n597) );
  INV_X1 U567 ( .A(G651), .ZN(n528) );
  NAND2_X1 U568 ( .A1(n786), .A2(G72), .ZN(n527) );
  NOR2_X1 U569 ( .A1(G651), .A2(G543), .ZN(n525) );
  XNOR2_X1 U570 ( .A(n525), .B(KEYINPUT64), .ZN(n787) );
  NAND2_X1 U571 ( .A1(G85), .A2(n787), .ZN(n526) );
  NAND2_X1 U572 ( .A1(n527), .A2(n526), .ZN(n533) );
  NAND2_X1 U573 ( .A1(G47), .A2(n790), .ZN(n531) );
  NOR2_X1 U574 ( .A1(G543), .A2(n528), .ZN(n529) );
  XOR2_X1 U575 ( .A(KEYINPUT1), .B(n529), .Z(n791) );
  NAND2_X1 U576 ( .A1(G60), .A2(n791), .ZN(n530) );
  NAND2_X1 U577 ( .A1(n531), .A2(n530), .ZN(n532) );
  OR2_X1 U578 ( .A1(n533), .A2(n532), .ZN(G290) );
  NOR2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n534) );
  XOR2_X2 U580 ( .A(KEYINPUT17), .B(n534), .Z(n989) );
  NAND2_X1 U581 ( .A1(G138), .A2(n989), .ZN(n536) );
  INV_X1 U582 ( .A(G2104), .ZN(n537) );
  NAND2_X1 U583 ( .A1(G102), .A2(n990), .ZN(n535) );
  NAND2_X1 U584 ( .A1(n536), .A2(n535), .ZN(n542) );
  INV_X1 U585 ( .A(G2105), .ZN(n538) );
  NOR2_X1 U586 ( .A1(G2104), .A2(n538), .ZN(n985) );
  NAND2_X1 U587 ( .A1(G126), .A2(n985), .ZN(n540) );
  NOR2_X1 U588 ( .A1(n538), .A2(n537), .ZN(n986) );
  NAND2_X1 U589 ( .A1(G114), .A2(n986), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U591 ( .A1(n542), .A2(n541), .ZN(G164) );
  NAND2_X1 U592 ( .A1(n989), .A2(G137), .ZN(n543) );
  XNOR2_X1 U593 ( .A(KEYINPUT68), .B(n543), .ZN(n552) );
  NAND2_X1 U594 ( .A1(G125), .A2(n985), .ZN(n544) );
  XNOR2_X1 U595 ( .A(n544), .B(KEYINPUT66), .ZN(n550) );
  NAND2_X1 U596 ( .A1(G101), .A2(n990), .ZN(n545) );
  XNOR2_X1 U597 ( .A(n545), .B(KEYINPUT67), .ZN(n546) );
  XNOR2_X1 U598 ( .A(n546), .B(KEYINPUT23), .ZN(n548) );
  NAND2_X1 U599 ( .A1(G113), .A2(n986), .ZN(n547) );
  AND2_X1 U600 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U601 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X2 U602 ( .A(n553), .B(KEYINPUT65), .ZN(G160) );
  XOR2_X1 U603 ( .A(KEYINPUT81), .B(KEYINPUT2), .Z(n555) );
  NAND2_X1 U604 ( .A1(G73), .A2(n786), .ZN(n554) );
  XNOR2_X1 U605 ( .A(n555), .B(n554), .ZN(n562) );
  NAND2_X1 U606 ( .A1(n790), .A2(G48), .ZN(n557) );
  NAND2_X1 U607 ( .A1(G86), .A2(n787), .ZN(n556) );
  NAND2_X1 U608 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U609 ( .A1(n791), .A2(G61), .ZN(n558) );
  XOR2_X1 U610 ( .A(KEYINPUT80), .B(n558), .Z(n559) );
  NOR2_X1 U611 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U612 ( .A1(n562), .A2(n561), .ZN(G305) );
  NAND2_X1 U613 ( .A1(n791), .A2(G64), .ZN(n564) );
  NAND2_X1 U614 ( .A1(n790), .A2(G52), .ZN(n563) );
  NAND2_X1 U615 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U616 ( .A(KEYINPUT70), .B(n565), .ZN(n570) );
  NAND2_X1 U617 ( .A1(n786), .A2(G77), .ZN(n567) );
  NAND2_X1 U618 ( .A1(G90), .A2(n787), .ZN(n566) );
  NAND2_X1 U619 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U620 ( .A(KEYINPUT9), .B(n568), .Z(n569) );
  NOR2_X1 U621 ( .A1(n570), .A2(n569), .ZN(G171) );
  INV_X1 U622 ( .A(G171), .ZN(G301) );
  NAND2_X1 U623 ( .A1(n786), .A2(G78), .ZN(n572) );
  NAND2_X1 U624 ( .A1(G91), .A2(n787), .ZN(n571) );
  NAND2_X1 U625 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U626 ( .A1(G65), .A2(n791), .ZN(n573) );
  XNOR2_X1 U627 ( .A(KEYINPUT71), .B(n573), .ZN(n574) );
  NOR2_X1 U628 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U629 ( .A1(n790), .A2(G53), .ZN(n576) );
  NAND2_X1 U630 ( .A1(n577), .A2(n576), .ZN(G299) );
  NAND2_X1 U631 ( .A1(G51), .A2(n790), .ZN(n579) );
  NAND2_X1 U632 ( .A1(G63), .A2(n791), .ZN(n578) );
  NAND2_X1 U633 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U634 ( .A(KEYINPUT6), .B(n580), .ZN(n587) );
  NAND2_X1 U635 ( .A1(G89), .A2(n787), .ZN(n581) );
  XNOR2_X1 U636 ( .A(n581), .B(KEYINPUT4), .ZN(n583) );
  NAND2_X1 U637 ( .A1(G76), .A2(n786), .ZN(n582) );
  NAND2_X1 U638 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U639 ( .A(KEYINPUT77), .B(n584), .ZN(n585) );
  XNOR2_X1 U640 ( .A(KEYINPUT5), .B(n585), .ZN(n586) );
  NOR2_X1 U641 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U642 ( .A(KEYINPUT7), .B(n588), .Z(G168) );
  XOR2_X1 U643 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U644 ( .A1(n786), .A2(G75), .ZN(n590) );
  NAND2_X1 U645 ( .A1(G88), .A2(n787), .ZN(n589) );
  NAND2_X1 U646 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U647 ( .A(KEYINPUT83), .B(n591), .ZN(n596) );
  NAND2_X1 U648 ( .A1(G50), .A2(n790), .ZN(n593) );
  NAND2_X1 U649 ( .A1(G62), .A2(n791), .ZN(n592) );
  NAND2_X1 U650 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U651 ( .A(KEYINPUT82), .B(n594), .Z(n595) );
  NAND2_X1 U652 ( .A1(n596), .A2(n595), .ZN(G303) );
  INV_X1 U653 ( .A(G303), .ZN(G166) );
  NAND2_X1 U654 ( .A1(G49), .A2(n790), .ZN(n599) );
  NAND2_X1 U655 ( .A1(G87), .A2(n597), .ZN(n598) );
  NAND2_X1 U656 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U657 ( .A1(n791), .A2(n600), .ZN(n602) );
  NAND2_X1 U658 ( .A1(G651), .A2(G74), .ZN(n601) );
  NAND2_X1 U659 ( .A1(n602), .A2(n601), .ZN(G288) );
  NAND2_X1 U660 ( .A1(G105), .A2(n990), .ZN(n603) );
  XNOR2_X1 U661 ( .A(n603), .B(KEYINPUT38), .ZN(n610) );
  NAND2_X1 U662 ( .A1(G129), .A2(n985), .ZN(n605) );
  NAND2_X1 U663 ( .A1(G141), .A2(n989), .ZN(n604) );
  NAND2_X1 U664 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U665 ( .A1(n986), .A2(G117), .ZN(n606) );
  XOR2_X1 U666 ( .A(KEYINPUT92), .B(n606), .Z(n607) );
  NOR2_X1 U667 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U668 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U669 ( .A(KEYINPUT93), .B(n611), .Z(n983) );
  NAND2_X1 U670 ( .A1(G1996), .A2(n983), .ZN(n612) );
  XNOR2_X1 U671 ( .A(n612), .B(KEYINPUT94), .ZN(n621) );
  XOR2_X1 U672 ( .A(G1991), .B(KEYINPUT91), .Z(n878) );
  NAND2_X1 U673 ( .A1(G119), .A2(n985), .ZN(n614) );
  NAND2_X1 U674 ( .A1(G131), .A2(n989), .ZN(n613) );
  NAND2_X1 U675 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U676 ( .A1(n990), .A2(G95), .ZN(n615) );
  XOR2_X1 U677 ( .A(KEYINPUT90), .B(n615), .Z(n616) );
  NOR2_X1 U678 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U679 ( .A1(n986), .A2(G107), .ZN(n618) );
  NAND2_X1 U680 ( .A1(n619), .A2(n618), .ZN(n981) );
  NAND2_X1 U681 ( .A1(n878), .A2(n981), .ZN(n620) );
  NAND2_X1 U682 ( .A1(n621), .A2(n620), .ZN(n746) );
  INV_X1 U683 ( .A(n746), .ZN(n851) );
  XOR2_X1 U684 ( .A(G1986), .B(G290), .Z(n924) );
  NAND2_X1 U685 ( .A1(n851), .A2(n924), .ZN(n623) );
  NOR2_X1 U686 ( .A1(G164), .A2(G1384), .ZN(n636) );
  NAND2_X1 U687 ( .A1(G160), .A2(G40), .ZN(n622) );
  NOR2_X1 U688 ( .A1(n636), .A2(n622), .ZN(n755) );
  NAND2_X1 U689 ( .A1(n623), .A2(n755), .ZN(n635) );
  XNOR2_X1 U690 ( .A(KEYINPUT89), .B(KEYINPUT36), .ZN(n634) );
  NAND2_X1 U691 ( .A1(G128), .A2(n985), .ZN(n625) );
  NAND2_X1 U692 ( .A1(G116), .A2(n986), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U694 ( .A(KEYINPUT35), .B(n626), .ZN(n632) );
  NAND2_X1 U695 ( .A1(G140), .A2(n989), .ZN(n628) );
  NAND2_X1 U696 ( .A1(G104), .A2(n990), .ZN(n627) );
  NAND2_X1 U697 ( .A1(n628), .A2(n627), .ZN(n630) );
  XOR2_X1 U698 ( .A(KEYINPUT34), .B(KEYINPUT88), .Z(n629) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(n631) );
  NAND2_X1 U700 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U701 ( .A(n634), .B(n633), .ZN(n1001) );
  XNOR2_X1 U702 ( .A(G2067), .B(KEYINPUT37), .ZN(n753) );
  NOR2_X1 U703 ( .A1(n1001), .A2(n753), .ZN(n842) );
  NAND2_X1 U704 ( .A1(n842), .A2(n755), .ZN(n752) );
  NAND2_X1 U705 ( .A1(n635), .A2(n752), .ZN(n744) );
  XNOR2_X1 U706 ( .A(G1981), .B(G305), .ZN(n931) );
  AND2_X1 U707 ( .A1(G40), .A2(n636), .ZN(n637) );
  AND2_X1 U708 ( .A1(G160), .A2(n637), .ZN(n644) );
  NAND2_X1 U709 ( .A1(n700), .A2(G8), .ZN(n734) );
  XOR2_X1 U710 ( .A(G2078), .B(KEYINPUT25), .Z(n877) );
  NOR2_X1 U711 ( .A1(n877), .A2(n700), .ZN(n639) );
  INV_X1 U712 ( .A(n700), .ZN(n670) );
  XNOR2_X1 U713 ( .A(G1961), .B(KEYINPUT96), .ZN(n896) );
  NOR2_X1 U714 ( .A1(n670), .A2(n896), .ZN(n638) );
  NOR2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n689) );
  OR2_X1 U716 ( .A1(n689), .A2(G301), .ZN(n688) );
  INV_X1 U717 ( .A(G299), .ZN(n923) );
  NAND2_X1 U718 ( .A1(n670), .A2(G2072), .ZN(n640) );
  XNOR2_X1 U719 ( .A(n640), .B(KEYINPUT27), .ZN(n642) );
  AND2_X1 U720 ( .A1(G1956), .A2(n700), .ZN(n641) );
  NOR2_X1 U721 ( .A1(n642), .A2(n641), .ZN(n680) );
  NOR2_X1 U722 ( .A1(n923), .A2(n680), .ZN(n643) );
  XOR2_X1 U723 ( .A(n643), .B(KEYINPUT28), .Z(n684) );
  NAND2_X1 U724 ( .A1(n644), .A2(G1996), .ZN(n645) );
  XOR2_X1 U725 ( .A(KEYINPUT26), .B(n645), .Z(n657) );
  NAND2_X1 U726 ( .A1(n787), .A2(G81), .ZN(n646) );
  XNOR2_X1 U727 ( .A(n646), .B(KEYINPUT12), .ZN(n647) );
  XNOR2_X1 U728 ( .A(n647), .B(KEYINPUT72), .ZN(n649) );
  NAND2_X1 U729 ( .A1(G68), .A2(n786), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U731 ( .A(n650), .B(KEYINPUT13), .ZN(n652) );
  NAND2_X1 U732 ( .A1(G43), .A2(n790), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n791), .A2(G56), .ZN(n653) );
  XOR2_X1 U735 ( .A(KEYINPUT14), .B(n653), .Z(n654) );
  NOR2_X1 U736 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U737 ( .A(KEYINPUT73), .B(n656), .ZN(n939) );
  XNOR2_X1 U738 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n667) );
  NAND2_X1 U739 ( .A1(G66), .A2(n791), .ZN(n664) );
  NAND2_X1 U740 ( .A1(n790), .A2(G54), .ZN(n659) );
  NAND2_X1 U741 ( .A1(G92), .A2(n787), .ZN(n658) );
  NAND2_X1 U742 ( .A1(n659), .A2(n658), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n786), .A2(G79), .ZN(n660) );
  XOR2_X1 U744 ( .A(KEYINPUT74), .B(n660), .Z(n661) );
  NOR2_X1 U745 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U746 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U747 ( .A(n665), .B(KEYINPUT15), .ZN(n666) );
  XNOR2_X2 U748 ( .A(n667), .B(n666), .ZN(n1010) );
  INV_X1 U749 ( .A(n1010), .ZN(n784) );
  NAND2_X1 U750 ( .A1(G1341), .A2(n700), .ZN(n675) );
  AND2_X1 U751 ( .A1(n784), .A2(n675), .ZN(n668) );
  XNOR2_X1 U752 ( .A(n669), .B(KEYINPUT97), .ZN(n674) );
  NOR2_X1 U753 ( .A1(n670), .A2(G1348), .ZN(n672) );
  NOR2_X1 U754 ( .A1(G2067), .A2(n700), .ZN(n671) );
  NOR2_X1 U755 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U756 ( .A1(n674), .A2(n673), .ZN(n679) );
  NAND2_X1 U757 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U758 ( .A1(n1010), .A2(n677), .ZN(n678) );
  NAND2_X1 U759 ( .A1(n679), .A2(n678), .ZN(n682) );
  NAND2_X1 U760 ( .A1(n923), .A2(n680), .ZN(n681) );
  NAND2_X1 U761 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U762 ( .A1(n684), .A2(n683), .ZN(n686) );
  XOR2_X1 U763 ( .A(KEYINPUT29), .B(KEYINPUT98), .Z(n685) );
  XNOR2_X1 U764 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U765 ( .A1(n688), .A2(n687), .ZN(n699) );
  NAND2_X1 U766 ( .A1(n689), .A2(G301), .ZN(n690) );
  XNOR2_X1 U767 ( .A(n690), .B(KEYINPUT99), .ZN(n695) );
  NOR2_X1 U768 ( .A1(G1966), .A2(n734), .ZN(n711) );
  NOR2_X1 U769 ( .A1(G2084), .A2(n700), .ZN(n708) );
  NOR2_X1 U770 ( .A1(n711), .A2(n708), .ZN(n691) );
  NAND2_X1 U771 ( .A1(G8), .A2(n691), .ZN(n692) );
  XNOR2_X1 U772 ( .A(KEYINPUT30), .B(n692), .ZN(n693) );
  NOR2_X1 U773 ( .A1(n693), .A2(G168), .ZN(n694) );
  NOR2_X1 U774 ( .A1(n695), .A2(n694), .ZN(n697) );
  XNOR2_X1 U775 ( .A(n697), .B(n696), .ZN(n698) );
  NAND2_X1 U776 ( .A1(n699), .A2(n698), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n709), .A2(G286), .ZN(n705) );
  NOR2_X1 U778 ( .A1(G1971), .A2(n734), .ZN(n702) );
  NOR2_X1 U779 ( .A1(G2090), .A2(n700), .ZN(n701) );
  NOR2_X1 U780 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U781 ( .A1(n703), .A2(G303), .ZN(n704) );
  NAND2_X1 U782 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U783 ( .A1(n706), .A2(G8), .ZN(n707) );
  XNOR2_X1 U784 ( .A(n707), .B(KEYINPUT32), .ZN(n715) );
  NAND2_X1 U785 ( .A1(G8), .A2(n708), .ZN(n713) );
  INV_X1 U786 ( .A(n709), .ZN(n710) );
  NOR2_X1 U787 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U788 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U789 ( .A1(n715), .A2(n714), .ZN(n731) );
  INV_X1 U790 ( .A(n731), .ZN(n718) );
  INV_X1 U791 ( .A(G1971), .ZN(n933) );
  NAND2_X1 U792 ( .A1(G166), .A2(n933), .ZN(n717) );
  NOR2_X1 U793 ( .A1(G1976), .A2(G288), .ZN(n722) );
  INV_X1 U794 ( .A(n722), .ZN(n716) );
  NAND2_X1 U795 ( .A1(n717), .A2(n716), .ZN(n927) );
  NOR2_X1 U796 ( .A1(n718), .A2(n927), .ZN(n719) );
  NOR2_X1 U797 ( .A1(n734), .A2(n719), .ZN(n720) );
  NAND2_X1 U798 ( .A1(G1976), .A2(G288), .ZN(n928) );
  NAND2_X1 U799 ( .A1(n720), .A2(n928), .ZN(n721) );
  INV_X1 U800 ( .A(KEYINPUT33), .ZN(n724) );
  NAND2_X1 U801 ( .A1(n721), .A2(n724), .ZN(n727) );
  INV_X1 U802 ( .A(n734), .ZN(n738) );
  NAND2_X1 U803 ( .A1(n738), .A2(n722), .ZN(n723) );
  NOR2_X1 U804 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U805 ( .A(n725), .B(KEYINPUT100), .Z(n726) );
  NAND2_X1 U806 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U807 ( .A1(n931), .A2(n728), .ZN(n742) );
  NOR2_X1 U808 ( .A1(G2090), .A2(G303), .ZN(n729) );
  XOR2_X1 U809 ( .A(KEYINPUT101), .B(n729), .Z(n730) );
  NAND2_X1 U810 ( .A1(G8), .A2(n730), .ZN(n732) );
  NAND2_X1 U811 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U812 ( .A1(n734), .A2(n733), .ZN(n740) );
  NOR2_X1 U813 ( .A1(G1981), .A2(G305), .ZN(n735) );
  XOR2_X1 U814 ( .A(n735), .B(KEYINPUT24), .Z(n736) );
  XNOR2_X1 U815 ( .A(KEYINPUT95), .B(n736), .ZN(n737) );
  NAND2_X1 U816 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U817 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U818 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U819 ( .A1(n744), .A2(n743), .ZN(n759) );
  NOR2_X1 U820 ( .A1(G1996), .A2(n983), .ZN(n843) );
  NOR2_X1 U821 ( .A1(G1986), .A2(G290), .ZN(n745) );
  NOR2_X1 U822 ( .A1(n878), .A2(n981), .ZN(n839) );
  NOR2_X1 U823 ( .A1(n745), .A2(n839), .ZN(n747) );
  NOR2_X1 U824 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U825 ( .A1(n843), .A2(n748), .ZN(n749) );
  XNOR2_X1 U826 ( .A(n749), .B(KEYINPUT39), .ZN(n750) );
  XNOR2_X1 U827 ( .A(n750), .B(KEYINPUT102), .ZN(n751) );
  NAND2_X1 U828 ( .A1(n752), .A2(n751), .ZN(n754) );
  NAND2_X1 U829 ( .A1(n1001), .A2(n753), .ZN(n853) );
  NAND2_X1 U830 ( .A1(n754), .A2(n853), .ZN(n756) );
  NAND2_X1 U831 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U832 ( .A(n757), .B(KEYINPUT103), .ZN(n758) );
  OR2_X1 U833 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U834 ( .A(n760), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U835 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U836 ( .A(G132), .ZN(G219) );
  INV_X1 U837 ( .A(G82), .ZN(G220) );
  INV_X1 U838 ( .A(G120), .ZN(G236) );
  INV_X1 U839 ( .A(G69), .ZN(G235) );
  INV_X1 U840 ( .A(G108), .ZN(G238) );
  NAND2_X1 U841 ( .A1(G7), .A2(G661), .ZN(n761) );
  XNOR2_X1 U842 ( .A(n761), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U843 ( .A(G223), .ZN(n826) );
  NAND2_X1 U844 ( .A1(n826), .A2(G567), .ZN(n762) );
  XOR2_X1 U845 ( .A(KEYINPUT11), .B(n762), .Z(G234) );
  INV_X1 U846 ( .A(n939), .ZN(n763) );
  NAND2_X1 U847 ( .A1(n763), .A2(G860), .ZN(G153) );
  NOR2_X1 U848 ( .A1(n1010), .A2(G868), .ZN(n765) );
  INV_X1 U849 ( .A(G868), .ZN(n808) );
  NOR2_X1 U850 ( .A1(n808), .A2(G301), .ZN(n764) );
  NOR2_X1 U851 ( .A1(n765), .A2(n764), .ZN(G284) );
  NOR2_X1 U852 ( .A1(G286), .A2(n808), .ZN(n767) );
  NOR2_X1 U853 ( .A1(G868), .A2(G299), .ZN(n766) );
  NOR2_X1 U854 ( .A1(n767), .A2(n766), .ZN(G297) );
  INV_X1 U855 ( .A(G559), .ZN(n770) );
  NOR2_X1 U856 ( .A1(G860), .A2(n770), .ZN(n768) );
  NOR2_X1 U857 ( .A1(n1010), .A2(n768), .ZN(n769) );
  XOR2_X1 U858 ( .A(KEYINPUT16), .B(n769), .Z(G148) );
  NAND2_X1 U859 ( .A1(n770), .A2(n784), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n771), .A2(G868), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n939), .A2(n808), .ZN(n772) );
  NAND2_X1 U862 ( .A1(n773), .A2(n772), .ZN(G282) );
  NAND2_X1 U863 ( .A1(n985), .A2(G123), .ZN(n774) );
  XNOR2_X1 U864 ( .A(n774), .B(KEYINPUT18), .ZN(n776) );
  NAND2_X1 U865 ( .A1(G99), .A2(n990), .ZN(n775) );
  NAND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G111), .A2(n986), .ZN(n778) );
  NAND2_X1 U868 ( .A1(G135), .A2(n989), .ZN(n777) );
  NAND2_X1 U869 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n982) );
  XNOR2_X1 U871 ( .A(n982), .B(G2096), .ZN(n781) );
  XNOR2_X1 U872 ( .A(n781), .B(KEYINPUT78), .ZN(n783) );
  INV_X1 U873 ( .A(G2100), .ZN(n782) );
  NAND2_X1 U874 ( .A1(n783), .A2(n782), .ZN(G156) );
  NAND2_X1 U875 ( .A1(G559), .A2(n784), .ZN(n806) );
  XNOR2_X1 U876 ( .A(n939), .B(n806), .ZN(n785) );
  NOR2_X1 U877 ( .A1(n785), .A2(G860), .ZN(n797) );
  NAND2_X1 U878 ( .A1(n786), .A2(G80), .ZN(n789) );
  NAND2_X1 U879 ( .A1(G93), .A2(n787), .ZN(n788) );
  NAND2_X1 U880 ( .A1(n789), .A2(n788), .ZN(n796) );
  NAND2_X1 U881 ( .A1(G55), .A2(n790), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G67), .A2(n791), .ZN(n792) );
  NAND2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U884 ( .A(KEYINPUT79), .B(n794), .Z(n795) );
  OR2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n809) );
  XOR2_X1 U886 ( .A(n797), .B(n809), .Z(G145) );
  XNOR2_X1 U887 ( .A(n923), .B(G166), .ZN(n798) );
  XNOR2_X1 U888 ( .A(n798), .B(G290), .ZN(n805) );
  XNOR2_X1 U889 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n800) );
  XNOR2_X1 U890 ( .A(G288), .B(KEYINPUT19), .ZN(n799) );
  XNOR2_X1 U891 ( .A(n800), .B(n799), .ZN(n801) );
  XNOR2_X1 U892 ( .A(n809), .B(n801), .ZN(n802) );
  XNOR2_X1 U893 ( .A(G305), .B(n802), .ZN(n803) );
  XOR2_X1 U894 ( .A(n803), .B(n939), .Z(n804) );
  XNOR2_X1 U895 ( .A(n805), .B(n804), .ZN(n1011) );
  XOR2_X1 U896 ( .A(n1011), .B(n806), .Z(n807) );
  NOR2_X1 U897 ( .A1(n808), .A2(n807), .ZN(n811) );
  NOR2_X1 U898 ( .A1(G868), .A2(n809), .ZN(n810) );
  NOR2_X1 U899 ( .A1(n811), .A2(n810), .ZN(G295) );
  NAND2_X1 U900 ( .A1(G2078), .A2(G2084), .ZN(n812) );
  XOR2_X1 U901 ( .A(KEYINPUT20), .B(n812), .Z(n813) );
  NAND2_X1 U902 ( .A1(G2090), .A2(n813), .ZN(n814) );
  XNOR2_X1 U903 ( .A(KEYINPUT21), .B(n814), .ZN(n815) );
  NAND2_X1 U904 ( .A1(n815), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U905 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U906 ( .A1(G235), .A2(G236), .ZN(n816) );
  XOR2_X1 U907 ( .A(KEYINPUT86), .B(n816), .Z(n817) );
  NOR2_X1 U908 ( .A1(G238), .A2(n817), .ZN(n818) );
  NAND2_X1 U909 ( .A1(G57), .A2(n818), .ZN(n955) );
  NAND2_X1 U910 ( .A1(n955), .A2(G567), .ZN(n823) );
  NOR2_X1 U911 ( .A1(G220), .A2(G219), .ZN(n819) );
  XOR2_X1 U912 ( .A(KEYINPUT22), .B(n819), .Z(n820) );
  NOR2_X1 U913 ( .A1(G218), .A2(n820), .ZN(n821) );
  NAND2_X1 U914 ( .A1(G96), .A2(n821), .ZN(n956) );
  NAND2_X1 U915 ( .A1(n956), .A2(G2106), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n957) );
  NAND2_X1 U917 ( .A1(G661), .A2(G483), .ZN(n824) );
  XOR2_X1 U918 ( .A(KEYINPUT87), .B(n824), .Z(n825) );
  NOR2_X1 U919 ( .A1(n957), .A2(n825), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n828), .A2(G36), .ZN(G176) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U923 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G1), .A2(G3), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U926 ( .A(n830), .B(KEYINPUT104), .ZN(G188) );
  XNOR2_X1 U927 ( .A(G96), .B(KEYINPUT105), .ZN(G221) );
  NAND2_X1 U929 ( .A1(n986), .A2(G112), .ZN(n837) );
  NAND2_X1 U930 ( .A1(G136), .A2(n989), .ZN(n832) );
  NAND2_X1 U931 ( .A1(G100), .A2(n990), .ZN(n831) );
  NAND2_X1 U932 ( .A1(n832), .A2(n831), .ZN(n835) );
  NAND2_X1 U933 ( .A1(n985), .A2(G124), .ZN(n833) );
  XOR2_X1 U934 ( .A(KEYINPUT44), .B(n833), .Z(n834) );
  NOR2_X1 U935 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U936 ( .A1(n837), .A2(n836), .ZN(n838) );
  XOR2_X1 U937 ( .A(KEYINPUT112), .B(n838), .Z(G162) );
  NOR2_X1 U938 ( .A1(n839), .A2(n982), .ZN(n840) );
  XOR2_X1 U939 ( .A(KEYINPUT118), .B(n840), .Z(n841) );
  NOR2_X1 U940 ( .A1(n842), .A2(n841), .ZN(n847) );
  XOR2_X1 U941 ( .A(G2090), .B(G162), .Z(n844) );
  NOR2_X1 U942 ( .A1(n844), .A2(n843), .ZN(n845) );
  XOR2_X1 U943 ( .A(KEYINPUT51), .B(n845), .Z(n846) );
  NAND2_X1 U944 ( .A1(n847), .A2(n846), .ZN(n849) );
  XOR2_X1 U945 ( .A(G160), .B(G2084), .Z(n848) );
  NOR2_X1 U946 ( .A1(n849), .A2(n848), .ZN(n850) );
  NAND2_X1 U947 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U948 ( .A(n852), .B(KEYINPUT119), .ZN(n854) );
  NAND2_X1 U949 ( .A1(n854), .A2(n853), .ZN(n869) );
  NAND2_X1 U950 ( .A1(n986), .A2(G115), .ZN(n855) );
  XNOR2_X1 U951 ( .A(n855), .B(KEYINPUT114), .ZN(n857) );
  NAND2_X1 U952 ( .A1(G127), .A2(n985), .ZN(n856) );
  NAND2_X1 U953 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U954 ( .A(n858), .B(KEYINPUT47), .ZN(n860) );
  NAND2_X1 U955 ( .A1(G139), .A2(n989), .ZN(n859) );
  NAND2_X1 U956 ( .A1(n860), .A2(n859), .ZN(n863) );
  NAND2_X1 U957 ( .A1(G103), .A2(n990), .ZN(n861) );
  XNOR2_X1 U958 ( .A(KEYINPUT113), .B(n861), .ZN(n862) );
  NOR2_X1 U959 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U960 ( .A(KEYINPUT115), .B(n864), .Z(n998) );
  XOR2_X1 U961 ( .A(G2072), .B(n998), .Z(n866) );
  XOR2_X1 U962 ( .A(G164), .B(G2078), .Z(n865) );
  NOR2_X1 U963 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U964 ( .A(KEYINPUT50), .B(n867), .Z(n868) );
  NOR2_X1 U965 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U966 ( .A(KEYINPUT52), .B(n870), .ZN(n872) );
  INV_X1 U967 ( .A(KEYINPUT55), .ZN(n871) );
  NAND2_X1 U968 ( .A1(n872), .A2(n871), .ZN(n873) );
  NAND2_X1 U969 ( .A1(n873), .A2(G29), .ZN(n953) );
  XOR2_X1 U970 ( .A(G2072), .B(G33), .Z(n874) );
  NAND2_X1 U971 ( .A1(n874), .A2(G28), .ZN(n884) );
  XNOR2_X1 U972 ( .A(G2067), .B(G26), .ZN(n876) );
  XNOR2_X1 U973 ( .A(G1996), .B(G32), .ZN(n875) );
  NOR2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n882) );
  XNOR2_X1 U975 ( .A(n877), .B(G27), .ZN(n880) );
  XNOR2_X1 U976 ( .A(n878), .B(G25), .ZN(n879) );
  NOR2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n881) );
  NAND2_X1 U978 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U979 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U980 ( .A(KEYINPUT53), .B(n885), .Z(n888) );
  XOR2_X1 U981 ( .A(G34), .B(KEYINPUT54), .Z(n886) );
  XNOR2_X1 U982 ( .A(G2084), .B(n886), .ZN(n887) );
  NAND2_X1 U983 ( .A1(n888), .A2(n887), .ZN(n890) );
  XNOR2_X1 U984 ( .A(G35), .B(G2090), .ZN(n889) );
  NOR2_X1 U985 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U986 ( .A(KEYINPUT55), .B(n891), .ZN(n893) );
  INV_X1 U987 ( .A(G29), .ZN(n892) );
  NAND2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n894) );
  NAND2_X1 U989 ( .A1(n894), .A2(G11), .ZN(n895) );
  XNOR2_X1 U990 ( .A(n895), .B(KEYINPUT120), .ZN(n922) );
  XNOR2_X1 U991 ( .A(n896), .B(G5), .ZN(n910) );
  XOR2_X1 U992 ( .A(G1966), .B(G21), .Z(n907) );
  XNOR2_X1 U993 ( .A(G1348), .B(KEYINPUT59), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n897), .B(G4), .ZN(n901) );
  XNOR2_X1 U995 ( .A(G1956), .B(G20), .ZN(n899) );
  XNOR2_X1 U996 ( .A(G6), .B(G1981), .ZN(n898) );
  NOR2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n900) );
  NAND2_X1 U998 ( .A1(n901), .A2(n900), .ZN(n904) );
  XOR2_X1 U999 ( .A(G19), .B(G1341), .Z(n902) );
  XNOR2_X1 U1000 ( .A(KEYINPUT123), .B(n902), .ZN(n903) );
  NOR2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n905), .B(KEYINPUT60), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n908), .B(KEYINPUT124), .ZN(n909) );
  NOR2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1006 ( .A(KEYINPUT125), .B(n911), .Z(n918) );
  XNOR2_X1 U1007 ( .A(G22), .B(n933), .ZN(n913) );
  XOR2_X1 U1008 ( .A(G1976), .B(G23), .Z(n912) );
  NAND2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(n915) );
  XNOR2_X1 U1010 ( .A(G24), .B(G1986), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(KEYINPUT58), .B(n916), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(KEYINPUT61), .B(n919), .ZN(n920) );
  NOR2_X1 U1015 ( .A1(n920), .A2(G16), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(n950) );
  XNOR2_X1 U1017 ( .A(n923), .B(G1956), .ZN(n925) );
  NAND2_X1 U1018 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1019 ( .A1(n927), .A2(n926), .ZN(n929) );
  NAND2_X1 U1020 ( .A1(n929), .A2(n928), .ZN(n945) );
  XOR2_X1 U1021 ( .A(G168), .B(G1966), .Z(n930) );
  NOR2_X1 U1022 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1023 ( .A(KEYINPUT57), .B(n932), .Z(n943) );
  XNOR2_X1 U1024 ( .A(n1010), .B(G1348), .ZN(n935) );
  NOR2_X1 U1025 ( .A1(n933), .A2(G166), .ZN(n934) );
  NOR2_X1 U1026 ( .A1(n935), .A2(n934), .ZN(n938) );
  XNOR2_X1 U1027 ( .A(G1961), .B(KEYINPUT121), .ZN(n936) );
  XNOR2_X1 U1028 ( .A(n936), .B(G301), .ZN(n937) );
  NAND2_X1 U1029 ( .A1(n938), .A2(n937), .ZN(n941) );
  XNOR2_X1 U1030 ( .A(G1341), .B(n939), .ZN(n940) );
  NOR2_X1 U1031 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1032 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1033 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1034 ( .A(KEYINPUT122), .B(n946), .Z(n948) );
  XNOR2_X1 U1035 ( .A(G16), .B(KEYINPUT56), .ZN(n947) );
  NAND2_X1 U1036 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1037 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1038 ( .A(KEYINPUT126), .B(n951), .Z(n952) );
  NAND2_X1 U1039 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1040 ( .A(KEYINPUT62), .B(n954), .Z(G311) );
  XNOR2_X1 U1041 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  NOR2_X1 U1042 ( .A1(n956), .A2(n955), .ZN(G325) );
  INV_X1 U1043 ( .A(G325), .ZN(G261) );
  INV_X1 U1044 ( .A(n957), .ZN(G319) );
  XOR2_X1 U1045 ( .A(KEYINPUT41), .B(KEYINPUT111), .Z(n959) );
  XNOR2_X1 U1046 ( .A(G1996), .B(G1991), .ZN(n958) );
  XNOR2_X1 U1047 ( .A(n959), .B(n958), .ZN(n969) );
  XOR2_X1 U1048 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n961) );
  XNOR2_X1 U1049 ( .A(G1956), .B(G1976), .ZN(n960) );
  XNOR2_X1 U1050 ( .A(n961), .B(n960), .ZN(n965) );
  XOR2_X1 U1051 ( .A(G1986), .B(G1981), .Z(n963) );
  XNOR2_X1 U1052 ( .A(G1961), .B(G1971), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(n963), .B(n962), .ZN(n964) );
  XOR2_X1 U1054 ( .A(n965), .B(n964), .Z(n967) );
  XNOR2_X1 U1055 ( .A(G1966), .B(G2474), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(n967), .B(n966), .ZN(n968) );
  XOR2_X1 U1057 ( .A(n969), .B(n968), .Z(G229) );
  XOR2_X1 U1058 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n971) );
  XNOR2_X1 U1059 ( .A(KEYINPUT108), .B(G2678), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(n971), .B(n970), .ZN(n972) );
  XOR2_X1 U1061 ( .A(n972), .B(G2100), .Z(n974) );
  XNOR2_X1 U1062 ( .A(G2078), .B(G2072), .ZN(n973) );
  XNOR2_X1 U1063 ( .A(n974), .B(n973), .ZN(n978) );
  XOR2_X1 U1064 ( .A(KEYINPUT42), .B(G2096), .Z(n976) );
  XNOR2_X1 U1065 ( .A(G2090), .B(KEYINPUT106), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(n976), .B(n975), .ZN(n977) );
  XOR2_X1 U1067 ( .A(n978), .B(n977), .Z(n980) );
  XNOR2_X1 U1068 ( .A(G2067), .B(G2084), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(n980), .B(n979), .ZN(G227) );
  XNOR2_X1 U1070 ( .A(n982), .B(n981), .ZN(n984) );
  XNOR2_X1 U1071 ( .A(n984), .B(n983), .ZN(n997) );
  NAND2_X1 U1072 ( .A1(G130), .A2(n985), .ZN(n988) );
  NAND2_X1 U1073 ( .A1(G118), .A2(n986), .ZN(n987) );
  NAND2_X1 U1074 ( .A1(n988), .A2(n987), .ZN(n995) );
  NAND2_X1 U1075 ( .A1(G142), .A2(n989), .ZN(n992) );
  NAND2_X1 U1076 ( .A1(G106), .A2(n990), .ZN(n991) );
  NAND2_X1 U1077 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1078 ( .A(KEYINPUT45), .B(n993), .Z(n994) );
  NOR2_X1 U1079 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1080 ( .A(n997), .B(n996), .Z(n1000) );
  XNOR2_X1 U1081 ( .A(G160), .B(n998), .ZN(n999) );
  XNOR2_X1 U1082 ( .A(n1000), .B(n999), .ZN(n1006) );
  XNOR2_X1 U1083 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n1003) );
  XNOR2_X1 U1084 ( .A(n1001), .B(G164), .ZN(n1002) );
  XNOR2_X1 U1085 ( .A(n1003), .B(n1002), .ZN(n1004) );
  XOR2_X1 U1086 ( .A(G162), .B(n1004), .Z(n1005) );
  XNOR2_X1 U1087 ( .A(n1006), .B(n1005), .ZN(n1007) );
  NOR2_X1 U1088 ( .A1(G37), .A2(n1007), .ZN(G395) );
  XOR2_X1 U1089 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n1009) );
  XNOR2_X1 U1090 ( .A(G171), .B(G286), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(n1009), .B(n1008), .ZN(n1013) );
  XOR2_X1 U1092 ( .A(n1011), .B(n1010), .Z(n1012) );
  XNOR2_X1 U1093 ( .A(n1013), .B(n1012), .ZN(n1014) );
  NOR2_X1 U1094 ( .A1(G37), .A2(n1014), .ZN(G397) );
  XOR2_X1 U1095 ( .A(G2446), .B(G2451), .Z(n1016) );
  XNOR2_X1 U1096 ( .A(G1348), .B(G2430), .ZN(n1015) );
  XNOR2_X1 U1097 ( .A(n1016), .B(n1015), .ZN(n1022) );
  XOR2_X1 U1098 ( .A(G2443), .B(G2438), .Z(n1018) );
  XNOR2_X1 U1099 ( .A(G2454), .B(G2435), .ZN(n1017) );
  XNOR2_X1 U1100 ( .A(n1018), .B(n1017), .ZN(n1020) );
  XOR2_X1 U1101 ( .A(G1341), .B(G2427), .Z(n1019) );
  XNOR2_X1 U1102 ( .A(n1020), .B(n1019), .ZN(n1021) );
  XOR2_X1 U1103 ( .A(n1022), .B(n1021), .Z(n1023) );
  NAND2_X1 U1104 ( .A1(G14), .A2(n1023), .ZN(n1029) );
  NAND2_X1 U1105 ( .A1(G319), .A2(n1029), .ZN(n1026) );
  NOR2_X1 U1106 ( .A1(G229), .A2(G227), .ZN(n1024) );
  XNOR2_X1 U1107 ( .A(KEYINPUT49), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1108 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  NOR2_X1 U1109 ( .A1(G395), .A2(G397), .ZN(n1027) );
  NAND2_X1 U1110 ( .A1(n1028), .A2(n1027), .ZN(G225) );
  INV_X1 U1111 ( .A(G225), .ZN(G308) );
  INV_X1 U1112 ( .A(G57), .ZN(G237) );
  INV_X1 U1113 ( .A(n1029), .ZN(G401) );
endmodule

