//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G125), .ZN(new_n461));
  INV_X1    g036(.A(G113), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI22_X1  g038(.A1(new_n460), .A2(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(G2105), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n464), .A2(G2105), .B1(G101), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n460), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n471), .A2(KEYINPUT66), .A3(G137), .A4(new_n468), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n468), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT68), .Z(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OR3_X1    g058(.A1(new_n460), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT67), .B1(new_n460), .B2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n483), .B1(G136), .B2(new_n487), .ZN(G162));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n458), .C2(new_n459), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT69), .A2(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n468), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n489), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n489), .B(KEYINPUT70), .C1(new_n494), .C2(new_n495), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(G138), .B(new_n468), .C1(new_n458), .C2(new_n459), .ZN(new_n501));
  XOR2_X1   g076(.A(KEYINPUT71), .B(KEYINPUT4), .Z(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n471), .A2(G138), .A3(new_n468), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n510), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n519), .A2(G651), .B1(new_n526), .B2(G88), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n513), .B1(new_n522), .B2(new_n523), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G50), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT72), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n516), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n514), .A2(KEYINPUT74), .A3(new_n515), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G63), .ZN(new_n537));
  NOR3_X1   g112(.A1(new_n536), .A2(new_n537), .A3(new_n521), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n528), .A2(G51), .ZN(new_n541));
  INV_X1    g116(.A(G89), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n540), .B(new_n541), .C1(new_n525), .C2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n538), .A2(new_n543), .ZN(G168));
  NAND3_X1  g119(.A1(new_n534), .A2(G64), .A3(new_n535), .ZN(new_n545));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n521), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n528), .A2(G52), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n525), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(G171));
  XNOR2_X1  g126(.A(KEYINPUT75), .B(G81), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n525), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n528), .A2(G43), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n536), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n555), .B1(new_n558), .B2(G651), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n528), .A2(G53), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n526), .A2(G91), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n516), .A2(G65), .ZN(new_n568));
  AND2_X1   g143(.A1(G78), .A2(G543), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  INV_X1    g148(.A(G74), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n521), .B1(new_n536), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n528), .A2(new_n576), .A3(G49), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n576), .B1(new_n528), .B2(G49), .ZN(new_n578));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n577), .A2(new_n578), .B1(new_n579), .B2(new_n525), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT77), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(G288));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n514), .B2(new_n515), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n528), .A2(G48), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n592), .B(new_n593), .C1(new_n594), .C2(new_n525), .ZN(G305));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G60), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n536), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n526), .A2(G85), .B1(G47), .B2(new_n528), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND3_X1  g179(.A1(new_n526), .A2(KEYINPUT10), .A3(G92), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n525), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n517), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G54), .B2(new_n528), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G171), .B2(new_n615), .ZN(G284));
  OAI21_X1  g192(.A(new_n616), .B1(G171), .B2(new_n615), .ZN(G321));
  NAND2_X1  g193(.A1(G299), .A2(new_n615), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n615), .B2(G168), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(new_n615), .B2(G168), .ZN(G280));
  INV_X1    g196(.A(new_n614), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n558), .A2(G651), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n625), .A2(new_n554), .A3(new_n553), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(new_n615), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n614), .A2(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n615), .B2(new_n628), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n478), .A2(G123), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT80), .ZN(new_n632));
  INV_X1    g207(.A(G135), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n468), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n632), .B1(new_n486), .B2(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT81), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(G2096), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n471), .A2(new_n465), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n642), .B(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n639), .A2(new_n640), .A3(new_n645), .ZN(G156));
  XOR2_X1   g221(.A(KEYINPUT15), .B(G2435), .Z(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT82), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2427), .B(G2430), .Z(new_n650));
  OAI21_X1  g225(.A(KEYINPUT14), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT83), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n660), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(G401));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT17), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT84), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n665), .A2(new_n668), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n671), .B(new_n667), .C1(new_n664), .C2(new_n668), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n666), .A2(new_n664), .A3(new_n668), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2096), .B(G2100), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n679), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n679), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT85), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n693), .B(new_n694), .Z(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G23), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n581), .B2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT33), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT86), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NAND2_X1  g279(.A1(G166), .A2(G16), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G16), .B2(G22), .ZN(new_n706));
  INV_X1    g281(.A(G1971), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  NOR2_X1   g284(.A1(G6), .A2(G16), .ZN(new_n710));
  INV_X1    g285(.A(G305), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT32), .B(G1981), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n703), .A2(new_n704), .A3(new_n708), .A4(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(KEYINPUT34), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(KEYINPUT34), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G25), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n487), .A2(G131), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n722));
  INV_X1    g297(.A(G107), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(G2105), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G119), .B2(new_n478), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n720), .B1(new_n727), .B2(new_n719), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT35), .B(G1991), .Z(new_n729));
  XOR2_X1   g304(.A(new_n728), .B(new_n729), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n697), .A2(G24), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n603), .B2(new_n697), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(G1986), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n732), .A2(G1986), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n730), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n717), .A2(new_n718), .A3(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT36), .Z(new_n737));
  XOR2_X1   g312(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n738));
  NAND3_X1  g313(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n468), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G139), .B2(new_n487), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT90), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(new_n719), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n719), .B2(G33), .ZN(new_n746));
  INV_X1    g321(.A(G2072), .ZN(new_n747));
  NOR2_X1   g322(.A1(G16), .A2(G19), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n559), .B2(G16), .ZN(new_n749));
  OAI22_X1  g324(.A1(new_n746), .A2(new_n747), .B1(G1341), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n719), .A2(G35), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G162), .B2(new_n719), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G2090), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n750), .B(new_n755), .C1(G1341), .C2(new_n749), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n746), .A2(new_n747), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n697), .A2(G20), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT23), .Z(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G299), .B2(G16), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1956), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n697), .A2(G5), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G171), .B2(new_n697), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G1961), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(G1961), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n757), .A2(new_n761), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT93), .B(KEYINPUT31), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G11), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n769), .A2(G28), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n719), .B1(new_n769), .B2(G28), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT24), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n719), .B1(new_n772), .B2(G34), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n773), .A2(KEYINPUT91), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(G34), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n773), .B2(KEYINPUT91), .ZN(new_n776));
  OAI22_X1  g351(.A1(new_n474), .A2(new_n719), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G2084), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n768), .B1(new_n770), .B2(new_n771), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n622), .A2(new_n697), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G4), .B2(new_n697), .ZN(new_n781));
  INV_X1    g356(.A(G1348), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n783), .B1(new_n719), .B2(new_n638), .C1(new_n782), .C2(new_n781), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n719), .A2(G27), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G164), .B2(new_n719), .ZN(new_n786));
  INV_X1    g361(.A(G2078), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n777), .A2(new_n778), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n697), .A2(G21), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G168), .B2(new_n697), .ZN(new_n791));
  INV_X1    g366(.A(G1966), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n788), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n766), .A2(new_n784), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n796));
  INV_X1    g371(.A(G116), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G2105), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G128), .B2(new_n478), .ZN(new_n799));
  INV_X1    g374(.A(G140), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n486), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT87), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G29), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT88), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n719), .A2(G26), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT28), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G2067), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n719), .A2(G32), .ZN(new_n810));
  NAND3_X1  g385(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT26), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n478), .A2(G129), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n465), .A2(G105), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n487), .B2(G141), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n810), .B1(new_n816), .B2(new_n719), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT92), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT27), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G1996), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n756), .A2(new_n795), .A3(new_n809), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n737), .A2(new_n821), .ZN(G311));
  INV_X1    g397(.A(G311), .ZN(G150));
  NAND2_X1  g398(.A1(new_n622), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n534), .A2(G67), .A3(new_n535), .ZN(new_n826));
  NAND2_X1  g401(.A1(G80), .A2(G543), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n521), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n528), .A2(G55), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT95), .B(G93), .Z(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n525), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n626), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n559), .A2(new_n832), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n825), .B(new_n836), .Z(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  INV_X1    g413(.A(G860), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n832), .A2(new_n839), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(G145));
  AND2_X1   g419(.A1(KEYINPUT69), .A2(G114), .ZN(new_n845));
  NOR2_X1   g420(.A1(KEYINPUT69), .A2(G114), .ZN(new_n846));
  OAI21_X1  g421(.A(G2105), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n495), .ZN(new_n848));
  AOI22_X1  g423(.A1(G126), .A2(new_n478), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n507), .A2(KEYINPUT96), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT96), .B1(new_n507), .B2(new_n849), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n802), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n816), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n802), .B(new_n852), .ZN(new_n856));
  INV_X1    g431(.A(new_n816), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n744), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n855), .A2(new_n858), .ZN(new_n861));
  INV_X1    g436(.A(new_n743), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n478), .A2(G130), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n468), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n487), .B2(G142), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(new_n642), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n727), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n870), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n637), .B(new_n474), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(G162), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT97), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n872), .A2(new_n873), .A3(new_n878), .A4(new_n875), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n875), .B1(new_n872), .B2(new_n873), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n881), .A2(G37), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n880), .A2(KEYINPUT40), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT40), .B1(new_n880), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(G395));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n836), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n628), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n889));
  NAND2_X1  g464(.A1(G299), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT99), .A4(new_n570), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n622), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n614), .A2(new_n889), .A3(G299), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT41), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n896), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n888), .A2(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n887), .A2(new_n628), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n887), .A2(new_n628), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n894), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(G303), .B(G305), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT100), .B1(new_n599), .B2(new_n601), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n599), .A2(KEYINPUT100), .A3(new_n601), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n582), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n582), .A3(new_n908), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n911), .ZN(new_n913));
  INV_X1    g488(.A(new_n905), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n913), .A2(new_n909), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n904), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n918));
  INV_X1    g493(.A(new_n916), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n900), .A2(new_n919), .A3(new_n903), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n918), .B1(new_n917), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(G868), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(G868), .B2(new_n832), .ZN(G295));
  OAI21_X1  g499(.A(new_n923), .B1(G868), .B2(new_n832), .ZN(G331));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n834), .A2(G301), .A3(new_n835), .ZN(new_n928));
  AOI21_X1  g503(.A(G301), .B1(new_n834), .B2(new_n835), .ZN(new_n929));
  OAI21_X1  g504(.A(G286), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n836), .A2(G171), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n834), .A2(G301), .A3(new_n835), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(G168), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n897), .B(KEYINPUT102), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT103), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n894), .B2(KEYINPUT41), .ZN(new_n937));
  AOI211_X1 g512(.A(KEYINPUT103), .B(new_n896), .C1(new_n892), .C2(new_n893), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n934), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n894), .B1(new_n930), .B2(new_n933), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n919), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G37), .ZN(new_n943));
  INV_X1    g518(.A(new_n894), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n928), .A2(new_n929), .A3(G286), .ZN(new_n945));
  AOI21_X1  g520(.A(G168), .B1(new_n931), .B2(new_n932), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n898), .A2(new_n930), .A3(new_n933), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(new_n948), .A3(new_n916), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n942), .A2(KEYINPUT43), .A3(new_n943), .A4(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n943), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n916), .B1(new_n947), .B2(new_n948), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n927), .B1(new_n950), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n942), .A2(new_n951), .A3(new_n943), .A4(new_n949), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT43), .B1(new_n952), .B2(new_n953), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n927), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n926), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT44), .B1(new_n957), .B2(new_n958), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n955), .A2(new_n962), .A3(KEYINPUT104), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(G397));
  XNOR2_X1  g539(.A(new_n802), .B(new_n808), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT45), .B1(new_n852), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n461), .B1(new_n476), .B2(new_n477), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n462), .A2(new_n463), .ZN(new_n969));
  OAI21_X1  g544(.A(G2105), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n465), .A2(G101), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n473), .A2(G40), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT105), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n466), .A2(KEYINPUT105), .A3(G40), .A4(new_n473), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n967), .A2(new_n977), .ZN(new_n978));
  OR3_X1    g553(.A1(new_n965), .A2(KEYINPUT108), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT108), .B1(new_n965), .B2(new_n978), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n978), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n983));
  INV_X1    g558(.A(G1996), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT107), .B1(new_n978), .B2(G1996), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n816), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n982), .A2(G1996), .A3(new_n857), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n981), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  XOR2_X1   g565(.A(new_n726), .B(new_n729), .Z(new_n991));
  AOI21_X1  g566(.A(new_n990), .B1(new_n982), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g567(.A1(G290), .A2(G1986), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT106), .ZN(new_n994));
  NAND2_X1  g569(.A1(G290), .A2(G1986), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n996), .B(new_n982), .C1(new_n994), .C2(new_n995), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT112), .B(G1981), .Z(new_n999));
  NAND2_X1  g574(.A1(new_n711), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n1001));
  OR3_X1    g576(.A1(G288), .A2(new_n1001), .A3(G1976), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1001), .B1(G288), .B2(G1976), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n1005));
  INV_X1    g580(.A(new_n592), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n593), .B1(new_n525), .B2(new_n594), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1005), .B(G1981), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1005), .B1(G305), .B2(G1981), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1000), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT49), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(KEYINPUT49), .B(new_n1000), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1000), .B1(new_n1004), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n496), .B1(new_n503), .B2(new_n506), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G1384), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n974), .A2(new_n1018), .A3(new_n975), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G8), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(KEYINPUT110), .A2(KEYINPUT55), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(KEYINPUT110), .A2(KEYINPUT55), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g602(.A1(G166), .A2(new_n1021), .A3(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(G166), .A2(new_n1021), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(new_n1025), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n500), .B2(new_n507), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n974), .B(new_n975), .C1(new_n1031), .C2(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n507), .A2(new_n849), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT96), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n507), .A2(KEYINPUT96), .A3(new_n849), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1035), .A2(KEYINPUT45), .A3(new_n966), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT109), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n852), .A2(KEYINPUT109), .A3(KEYINPUT45), .A4(new_n966), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1032), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(G1971), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1033), .A2(new_n966), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(KEYINPUT50), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n976), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n508), .A2(new_n966), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT50), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(G2090), .ZN(new_n1049));
  OAI221_X1 g624(.A(G8), .B1(new_n1028), .B2(new_n1030), .C1(new_n1042), .C2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n583), .A2(new_n585), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n581), .A2(G1976), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1022), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1013), .A2(new_n1022), .A3(new_n1014), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1019), .A2(new_n1054), .A3(G8), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1058), .A2(KEYINPUT111), .A3(KEYINPUT52), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT111), .B1(new_n1058), .B2(KEYINPUT52), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1057), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1023), .B1(new_n1050), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT45), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1043), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1065), .B1(new_n977), .B2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1067), .A2(new_n1065), .A3(new_n974), .A4(new_n975), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1031), .A2(KEYINPUT45), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n792), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT50), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1031), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n974), .B(new_n975), .C1(KEYINPUT50), .C2(new_n1043), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1074), .A2(new_n1075), .A3(G2084), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1021), .B1(new_n1072), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G168), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT63), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(G8), .B1(new_n1042), .B2(new_n1049), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1030), .A2(new_n1028), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1081), .A2(new_n1084), .A3(new_n1050), .A4(new_n1062), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT50), .B1(new_n1017), .B2(G1384), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1086), .A2(new_n974), .A3(new_n975), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1031), .A2(new_n1073), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1088), .A2(new_n1090), .A3(G2090), .ZN(new_n1091));
  OAI21_X1  g666(.A(G8), .B1(new_n1042), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1083), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1093), .A2(new_n1050), .A3(new_n1062), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1080), .B1(new_n1094), .B2(new_n1079), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1064), .B1(new_n1085), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1040), .A2(new_n1039), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1032), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT56), .B(G2072), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(G1956), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT57), .B1(new_n566), .B2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n1105), .B(G299), .Z(new_n1106));
  NOR2_X1   g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1101), .B1(new_n1041), .B2(new_n1099), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1106), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT117), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1103), .A2(new_n1111), .A3(new_n1106), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(G1348), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1019), .A2(G2067), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n622), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1107), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT60), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT60), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1120), .B1(new_n1122), .B2(new_n622), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n782), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1020), .A2(new_n808), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT60), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1126), .A2(KEYINPUT119), .A3(new_n614), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1119), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1122), .A2(new_n1120), .A3(new_n622), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT119), .B1(new_n1126), .B2(new_n614), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1129), .A2(new_n1130), .A3(KEYINPUT60), .A4(new_n1118), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1110), .A2(new_n1134), .A3(new_n1112), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1109), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1133), .B1(new_n1107), .B2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT58), .B(G1341), .Z(new_n1138));
  AOI22_X1  g713(.A1(new_n1041), .A2(new_n984), .B1(new_n1019), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT59), .B1(new_n1139), .B2(new_n626), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1097), .A2(new_n1098), .A3(new_n984), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1019), .A2(new_n1138), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(new_n559), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1140), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1135), .A2(new_n1137), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1132), .B1(new_n1147), .B2(KEYINPUT118), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1135), .A2(new_n1137), .A3(new_n1146), .A4(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1117), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT53), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1152), .A2(G2078), .ZN(new_n1153));
  NAND3_X1  g728(.A1(G160), .A2(G40), .A3(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n967), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT122), .B1(new_n1155), .B2(new_n1097), .ZN(new_n1156));
  AOI21_X1  g731(.A(G1961), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1041), .A2(new_n787), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n1152), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1155), .A2(new_n1097), .A3(KEYINPUT122), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1158), .A2(new_n1160), .A3(G301), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT123), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1161), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1164), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1165), .A2(new_n1166), .A3(G301), .A4(new_n1160), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1157), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1018), .A2(KEYINPUT45), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT115), .B1(new_n1169), .B2(new_n976), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1170), .A2(new_n1070), .A3(new_n1069), .A4(new_n1153), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(G301), .B1(new_n1172), .B2(new_n1160), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1163), .A2(new_n1167), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT54), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1165), .A2(new_n1160), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(G171), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1180));
  AOI21_X1  g755(.A(KEYINPUT53), .B1(new_n1041), .B2(new_n787), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1176), .B1(new_n1182), .B2(G301), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1094), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(G168), .A2(new_n1021), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT121), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT51), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1170), .A2(new_n1070), .A3(new_n1069), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1076), .B1(new_n1189), .B2(new_n792), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1188), .B1(new_n1190), .B2(new_n1021), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1072), .A2(new_n1077), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT120), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1192), .A2(new_n1185), .B1(new_n1193), .B2(KEYINPUT51), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1185), .B1(new_n1078), .B2(new_n1186), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1193), .A2(KEYINPUT51), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1196), .ZN(new_n1197));
  OAI211_X1 g772(.A(new_n1191), .B(new_n1194), .C1(new_n1195), .C2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1177), .A2(new_n1184), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1096), .B1(new_n1151), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT124), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1093), .A2(new_n1173), .A3(new_n1050), .A4(new_n1062), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1202), .B1(new_n1198), .B2(KEYINPUT62), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1185), .ZN(new_n1204));
  OAI22_X1  g779(.A1(new_n1190), .A2(new_n1204), .B1(KEYINPUT120), .B2(new_n1187), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1078), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1205), .B1(new_n1206), .B2(new_n1188), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1190), .A2(KEYINPUT121), .A3(new_n1021), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1196), .B1(new_n1208), .B2(new_n1185), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1207), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1201), .B1(new_n1203), .B2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1192), .A2(new_n1186), .A3(G8), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1197), .B1(new_n1213), .B2(new_n1204), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1194), .A2(new_n1191), .ZN(new_n1215));
  OAI21_X1  g790(.A(KEYINPUT62), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1202), .ZN(new_n1217));
  AND4_X1   g792(.A1(new_n1201), .A2(new_n1216), .A3(new_n1211), .A4(new_n1217), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1212), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n998), .B1(new_n1200), .B2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g795(.A1(new_n993), .A2(new_n978), .ZN(new_n1221));
  XOR2_X1   g796(.A(new_n1221), .B(KEYINPUT48), .Z(new_n1222));
  NAND2_X1  g797(.A1(new_n727), .A2(new_n729), .ZN(new_n1223));
  OAI22_X1  g798(.A1(new_n990), .A2(new_n1223), .B1(G2067), .B2(new_n802), .ZN(new_n1224));
  AOI22_X1  g799(.A1(new_n992), .A2(new_n1222), .B1(new_n1224), .B2(new_n982), .ZN(new_n1225));
  INV_X1    g800(.A(KEYINPUT46), .ZN(new_n1226));
  NAND3_X1  g801(.A1(new_n985), .A2(new_n1226), .A3(new_n986), .ZN(new_n1227));
  XOR2_X1   g802(.A(new_n1227), .B(KEYINPUT125), .Z(new_n1228));
  AOI21_X1  g803(.A(new_n978), .B1(new_n965), .B2(new_n816), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1229), .B1(new_n987), .B2(KEYINPUT46), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g806(.A(KEYINPUT47), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1228), .A2(new_n1230), .A3(KEYINPUT47), .ZN(new_n1234));
  NAND3_X1  g809(.A1(new_n1233), .A2(KEYINPUT126), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1225), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g811(.A(KEYINPUT126), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1237));
  NOR2_X1   g812(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1220), .A2(new_n1238), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g814(.A1(new_n880), .A2(new_n882), .ZN(new_n1241));
  INV_X1    g815(.A(G319), .ZN(new_n1242));
  NOR2_X1   g816(.A1(G227), .A2(new_n1242), .ZN(new_n1243));
  XOR2_X1   g817(.A(new_n1243), .B(KEYINPUT127), .Z(new_n1244));
  NOR3_X1   g818(.A1(G401), .A2(G229), .A3(new_n1244), .ZN(new_n1245));
  NAND3_X1  g819(.A1(new_n1241), .A2(new_n1245), .A3(new_n959), .ZN(G225));
  INV_X1    g820(.A(G225), .ZN(G308));
endmodule


