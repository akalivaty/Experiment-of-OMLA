//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  INV_X1    g001(.A(G228gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n209), .B2(KEYINPUT2), .ZN(new_n210));
  INV_X1    g009(.A(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT74), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT74), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G148gat), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT75), .A4(G141gat), .ZN(new_n215));
  INV_X1    g014(.A(G141gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT73), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT73), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G141gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n219), .A3(G148gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT74), .B(G148gat), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT75), .B1(new_n222), .B2(G141gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n210), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT2), .B1(new_n216), .B2(new_n211), .ZN(new_n225));
  NAND2_X1  g024(.A1(G141gat), .A2(G148gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(new_n206), .A3(new_n209), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G211gat), .B(G218gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT70), .B(G211gat), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT22), .B1(new_n232), .B2(G218gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(G197gat), .B(G204gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n231), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G218gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(KEYINPUT70), .A2(G211gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(KEYINPUT70), .A2(G211gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n234), .B(new_n230), .C1(new_n241), .C2(KEYINPUT22), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT29), .B1(new_n236), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n229), .B1(new_n243), .B2(KEYINPUT3), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n236), .A2(new_n242), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n224), .A2(new_n246), .A3(new_n228), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT29), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n205), .B(new_n244), .C1(new_n249), .C2(KEYINPUT82), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n227), .A2(new_n206), .A3(new_n209), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n212), .A2(new_n214), .A3(G141gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT75), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n220), .A3(new_n215), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n251), .B1(new_n255), .B2(new_n210), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT29), .B1(new_n256), .B2(new_n246), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT82), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n257), .A2(new_n258), .A3(new_n245), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n202), .B1(new_n250), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n205), .ZN(new_n261));
  INV_X1    g060(.A(new_n242), .ZN(new_n262));
  INV_X1    g061(.A(new_n240), .ZN(new_n263));
  OAI21_X1  g062(.A(G218gat), .B1(new_n263), .B2(new_n238), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT22), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n230), .B1(new_n266), .B2(new_n234), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n248), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n246), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n261), .B1(new_n269), .B2(new_n229), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n258), .B1(new_n257), .B2(new_n245), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n249), .A2(KEYINPUT82), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT83), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n260), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G22gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n249), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n205), .B1(new_n276), .B2(new_n244), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n274), .A2(KEYINPUT84), .A3(new_n275), .A4(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G78gat), .B(G106gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(G50gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n277), .B1(new_n260), .B2(new_n273), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n275), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n274), .A2(new_n278), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT84), .B1(new_n287), .B2(G22gat), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n284), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(KEYINPUT85), .A3(G22gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT85), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(new_n285), .B2(new_n275), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n283), .B1(new_n285), .B2(new_n275), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT86), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n290), .A2(new_n292), .A3(new_n293), .A4(KEYINPUT86), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n289), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n245), .ZN(new_n299));
  INV_X1    g098(.A(G226gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(new_n204), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT27), .B(G183gat), .ZN(new_n303));
  INV_X1    g102(.A(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT28), .ZN(new_n306));
  NAND2_X1  g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT26), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NOR3_X1   g109(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n311));
  INV_X1    g110(.A(G183gat), .ZN(new_n312));
  OAI22_X1  g111(.A1(new_n310), .A2(new_n311), .B1(new_n312), .B2(new_n304), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  OR2_X1    g113(.A1(new_n308), .A2(KEYINPUT23), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n316), .B1(new_n308), .B2(KEYINPUT23), .ZN(new_n317));
  NAND3_X1  g116(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT66), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n307), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n315), .A2(new_n317), .A3(new_n318), .A4(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT24), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(G183gat), .A3(G190gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(G183gat), .B(G190gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(new_n322), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n308), .A2(KEYINPUT23), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT64), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n308), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n329), .A2(new_n315), .A3(new_n307), .A4(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n316), .B1(new_n331), .B2(new_n325), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n326), .B1(new_n332), .B2(KEYINPUT65), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT65), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n334), .B(new_n316), .C1(new_n331), .C2(new_n325), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n314), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n302), .B1(new_n336), .B2(KEYINPUT29), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n336), .A2(new_n302), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n299), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n332), .A2(KEYINPUT65), .ZN(new_n341));
  INV_X1    g140(.A(new_n326), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n335), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n314), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT71), .B1(new_n345), .B2(new_n301), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n336), .A2(new_n347), .A3(new_n302), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n337), .B(new_n245), .C1(new_n346), .C2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  NAND3_X1  g151(.A1(new_n340), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT30), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n353), .A2(KEYINPUT72), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n353), .B2(KEYINPUT72), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n352), .B1(new_n340), .B2(new_n349), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(G1gat), .B(G29gat), .Z(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT78), .ZN(new_n360));
  XNOR2_X1  g159(.A(G57gat), .B(G85gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT79), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n360), .B(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G127gat), .B(G134gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT67), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G127gat), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT67), .B1(new_n370), .B2(G134gat), .ZN(new_n371));
  INV_X1    g170(.A(G120gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G113gat), .ZN(new_n373));
  INV_X1    g172(.A(G113gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G120gat), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  OAI22_X1  g175(.A1(new_n369), .A2(new_n371), .B1(KEYINPUT1), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(KEYINPUT1), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n367), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n256), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n381), .A2(KEYINPUT4), .A3(new_n256), .ZN(new_n385));
  INV_X1    g184(.A(new_n247), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n380), .B1(new_n256), .B2(new_n246), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n384), .B(new_n385), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT76), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n229), .A2(new_n380), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n382), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n390), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n229), .A2(KEYINPUT76), .A3(new_n380), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n389), .A2(new_n390), .B1(KEYINPUT5), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT5), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n388), .A2(new_n398), .A3(new_n394), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n366), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n399), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(KEYINPUT5), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(new_n394), .B2(new_n388), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n403), .A3(new_n365), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT6), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n400), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n401), .A2(new_n403), .A3(KEYINPUT6), .A4(new_n365), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n358), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n345), .A2(new_n381), .ZN(new_n410));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n336), .A2(new_n380), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n410), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT32), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT68), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT68), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(new_n417), .A3(KEYINPUT32), .ZN(new_n418));
  XNOR2_X1  g217(.A(G15gat), .B(G43gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(G71gat), .B(G99gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n421), .B1(new_n414), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n416), .A2(new_n418), .A3(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n414), .B(KEYINPUT32), .C1(new_n422), .C2(new_n421), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n413), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT34), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n411), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n429), .A2(KEYINPUT69), .ZN(new_n430));
  INV_X1    g229(.A(new_n427), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT34), .B1(new_n431), .B2(new_n412), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(KEYINPUT69), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n433), .A2(new_n432), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n436), .A2(new_n425), .A3(new_n424), .A4(new_n430), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NOR4_X1   g237(.A1(new_n298), .A2(new_n409), .A3(KEYINPUT35), .A4(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n296), .A2(new_n297), .ZN(new_n441));
  INV_X1    g240(.A(new_n289), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n438), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(KEYINPUT88), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n298), .B2(new_n438), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n409), .A2(KEYINPUT80), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n358), .A2(new_n449), .A3(new_n408), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n445), .A2(new_n447), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT35), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n440), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n448), .A2(new_n450), .A3(new_n298), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT36), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n438), .B(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n408), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT37), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n352), .A2(new_n458), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n357), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n337), .B1(new_n302), .B2(new_n336), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n458), .B1(new_n461), .B2(new_n245), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n337), .B(new_n299), .C1(new_n346), .C2(new_n348), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT38), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n457), .A2(new_n353), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT38), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n340), .A2(new_n349), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT37), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n467), .B1(new_n460), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n388), .A2(new_n394), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n393), .A2(new_n395), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n471), .B(KEYINPUT39), .C1(new_n394), .C2(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n473), .B(new_n366), .C1(KEYINPUT39), .C2(new_n471), .ZN(new_n474));
  NOR2_X1   g273(.A1(KEYINPUT87), .A2(KEYINPUT40), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n475), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n404), .A3(new_n477), .ZN(new_n478));
  OAI22_X1  g277(.A1(new_n466), .A2(new_n470), .B1(new_n478), .B2(new_n358), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n454), .B(new_n456), .C1(new_n479), .C2(new_n298), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n453), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT16), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n482), .B1(new_n483), .B2(G1gat), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(G1gat), .B2(new_n482), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(G8gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(G29gat), .A2(G36gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT14), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G29gat), .A2(G36gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G43gat), .B(G50gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(KEYINPUT15), .A3(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n490), .B(KEYINPUT90), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n492), .B(KEYINPUT15), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n486), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(KEYINPUT17), .ZN(new_n499));
  INV_X1    g298(.A(new_n486), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G229gat), .A2(G233gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT18), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT91), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n501), .A2(KEYINPUT91), .A3(KEYINPUT18), .A4(new_n502), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT18), .B1(new_n501), .B2(new_n502), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n486), .A2(new_n497), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n498), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n502), .B(KEYINPUT13), .Z(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G113gat), .B(G141gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G169gat), .B(G197gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n519), .B(KEYINPUT12), .Z(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n507), .A2(new_n514), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n521), .B1(new_n507), .B2(new_n514), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n481), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT92), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT92), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n481), .A2(new_n529), .A3(new_n526), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT99), .ZN(new_n532));
  INV_X1    g331(.A(G64gat), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n533), .A2(G57gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(G57gat), .ZN(new_n535));
  AND2_X1   g334(.A1(G71gat), .A2(G78gat), .ZN(new_n536));
  OAI22_X1  g335(.A1(new_n534), .A2(new_n535), .B1(KEYINPUT9), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G71gat), .B(G78gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n486), .B1(KEYINPUT21), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT94), .ZN(new_n541));
  NAND2_X1  g340(.A1(G231gat), .A2(G233gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT93), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n541), .B(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n539), .A2(KEYINPUT21), .ZN(new_n547));
  XNOR2_X1  g346(.A(G127gat), .B(G155gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G183gat), .B(G211gat), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n546), .A2(new_n551), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G85gat), .A2(G92gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT7), .ZN(new_n556));
  NAND2_X1  g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557));
  INV_X1    g356(.A(G85gat), .ZN(new_n558));
  INV_X1    g357(.A(G92gat), .ZN(new_n559));
  AOI22_X1  g358(.A1(KEYINPUT8), .A2(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G99gat), .B(G106gat), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n561), .B(new_n562), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT97), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n497), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n561), .B(new_n562), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n566), .A2(KEYINPUT97), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(KEYINPUT97), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n499), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT41), .ZN(new_n571));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n572), .B(KEYINPUT95), .Z(new_n573));
  OAI211_X1 g372(.A(new_n565), .B(new_n570), .C1(new_n571), .C2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G190gat), .B(G218gat), .Z(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT98), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n574), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n571), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT96), .ZN(new_n579));
  XOR2_X1   g378(.A(G134gat), .B(G162gat), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n577), .B(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n532), .B1(new_n554), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n581), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n577), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n552), .A2(new_n553), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(KEYINPUT99), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n539), .A2(KEYINPUT10), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n564), .A2(KEYINPUT101), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n567), .A2(new_n568), .A3(new_n590), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT101), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n539), .B1(new_n566), .B2(KEYINPUT100), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(KEYINPUT100), .B2(new_n566), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT100), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n563), .A2(new_n598), .A3(new_n539), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT10), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n589), .B1(new_n595), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n589), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n597), .A2(new_n602), .A3(new_n599), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G120gat), .B(G148gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT103), .ZN(new_n606));
  XNOR2_X1  g405(.A(G176gat), .B(G204gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n603), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n608), .B1(new_n610), .B2(KEYINPUT102), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n601), .B(new_n611), .C1(KEYINPUT102), .C2(new_n610), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n588), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n531), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(new_n408), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(G1gat), .Z(G1324gat));
  INV_X1    g416(.A(new_n358), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n531), .A2(new_n618), .A3(new_n614), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT16), .B(G8gat), .Z(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT42), .ZN(new_n621));
  OR3_X1    g420(.A1(new_n619), .A2(KEYINPUT105), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT105), .B1(new_n619), .B2(new_n621), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT42), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n620), .B2(KEYINPUT104), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n626), .B1(KEYINPUT104), .B2(new_n620), .ZN(new_n627));
  OAI22_X1  g426(.A1(new_n619), .A2(new_n627), .B1(new_n625), .B2(G8gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(G1325gat));
  OR2_X1    g428(.A1(new_n456), .A2(KEYINPUT106), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n456), .A2(KEYINPUT106), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(G15gat), .B1(new_n615), .B2(new_n632), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n438), .A2(G15gat), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n615), .B2(new_n634), .ZN(G1326gat));
  NOR2_X1   g434(.A1(new_n615), .A2(new_n443), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT43), .B(G22gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(G1327gat));
  NOR3_X1   g437(.A1(new_n585), .A2(new_n613), .A3(new_n586), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n408), .A2(G29gat), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n531), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT45), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n448), .A2(new_n450), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT88), .B1(new_n443), .B2(new_n444), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n298), .A2(new_n438), .A3(new_n446), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n439), .B1(new_n647), .B2(KEYINPUT35), .ZN(new_n648));
  INV_X1    g447(.A(new_n480), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n582), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n481), .A2(KEYINPUT44), .A3(new_n582), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n613), .B(KEYINPUT107), .Z(new_n655));
  AND3_X1   g454(.A1(new_n655), .A2(new_n526), .A3(new_n554), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(G29gat), .B1(new_n657), .B2(new_n408), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n642), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n643), .A2(new_n658), .A3(new_n659), .ZN(G1328gat));
  NAND2_X1  g459(.A1(new_n531), .A2(new_n639), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n358), .A2(G36gat), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  OR3_X1    g462(.A1(new_n661), .A2(KEYINPUT46), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(G36gat), .B1(new_n657), .B2(new_n358), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT46), .B1(new_n661), .B2(new_n663), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(G1329gat));
  OAI21_X1  g466(.A(G43gat), .B1(new_n657), .B2(new_n456), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n438), .A2(G43gat), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n531), .A2(new_n639), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(KEYINPUT47), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n672));
  INV_X1    g471(.A(new_n632), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n652), .A2(new_n673), .A3(new_n653), .A4(new_n656), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(G43gat), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n672), .B1(new_n670), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI211_X1 g477(.A(KEYINPUT109), .B(new_n672), .C1(new_n670), .C2(new_n675), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n671), .B1(new_n678), .B2(new_n679), .ZN(G1330gat));
  OAI21_X1  g479(.A(G50gat), .B1(new_n657), .B2(new_n443), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n443), .A2(G50gat), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n531), .A2(new_n639), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT48), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n681), .A2(KEYINPUT48), .A3(new_n683), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(G1331gat));
  NOR3_X1   g487(.A1(new_n588), .A2(new_n526), .A3(new_n655), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n481), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n457), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g491(.A1(new_n690), .A2(new_n618), .ZN(new_n693));
  NOR2_X1   g492(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n694));
  AND2_X1   g493(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n693), .B2(new_n694), .ZN(G1333gat));
  NAND2_X1  g496(.A1(new_n690), .A2(new_n673), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n438), .A2(G71gat), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n698), .A2(G71gat), .B1(new_n690), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g500(.A1(new_n690), .A2(new_n298), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g502(.A1(new_n526), .A2(new_n586), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n613), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n654), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G85gat), .B1(new_n708), .B2(new_n408), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n585), .B1(new_n453), .B2(new_n480), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n710), .A2(KEYINPUT51), .A3(new_n704), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT51), .B1(new_n710), .B2(new_n704), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n457), .A2(new_n558), .A3(new_n613), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n709), .B1(new_n713), .B2(new_n714), .ZN(G1336gat));
  NAND4_X1  g514(.A1(new_n652), .A2(new_n618), .A3(new_n653), .A4(new_n707), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G92gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT110), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT52), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n655), .A2(G92gat), .A3(new_n358), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n711), .B2(new_n712), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n717), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n720), .B1(new_n717), .B2(new_n722), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n719), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n717), .A2(new_n722), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT111), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n717), .B2(KEYINPUT110), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n717), .A2(new_n720), .A3(new_n722), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n725), .A2(new_n731), .ZN(G1337gat));
  OAI21_X1  g531(.A(G99gat), .B1(new_n708), .B2(new_n632), .ZN(new_n733));
  OR3_X1    g532(.A1(new_n438), .A2(new_n706), .A3(G99gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n713), .B2(new_n734), .ZN(G1338gat));
  OAI21_X1  g534(.A(G106gat), .B1(new_n708), .B2(new_n443), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n655), .A2(new_n443), .A3(G106gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n711), .B2(new_n712), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT53), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT53), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n736), .A2(new_n741), .A3(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(G1339gat));
  NAND2_X1  g542(.A1(new_n510), .A2(new_n512), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n501), .B2(new_n502), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n745), .A2(KEYINPUT112), .A3(new_n519), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n745), .A2(new_n519), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n747), .A2(KEYINPUT112), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n613), .A2(new_n522), .A3(new_n746), .A4(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750));
  INV_X1    g549(.A(new_n600), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n751), .A2(new_n591), .A3(new_n602), .A4(new_n594), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n601), .A2(KEYINPUT54), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT54), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n754), .B(new_n589), .C1(new_n595), .C2(new_n600), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n608), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n750), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n601), .A2(KEYINPUT54), .A3(new_n752), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n758), .A2(KEYINPUT55), .A3(new_n608), .A4(new_n755), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n612), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n749), .B1(new_n760), .B2(new_n525), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT113), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n763), .B(new_n749), .C1(new_n760), .C2(new_n525), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n585), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n522), .A3(new_n746), .ZN(new_n766));
  OR3_X1    g565(.A1(new_n760), .A2(new_n585), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n554), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n583), .A2(new_n587), .A3(new_n525), .A4(new_n706), .ZN(new_n770));
  AOI211_X1 g569(.A(new_n438), .B(new_n298), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n618), .A2(new_n408), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n773), .A2(new_n374), .A3(new_n525), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n408), .B1(new_n769), .B2(new_n770), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n445), .A2(new_n447), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n775), .A2(new_n358), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(G113gat), .B1(new_n777), .B2(new_n526), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n774), .A2(new_n778), .ZN(G1340gat));
  NOR3_X1   g578(.A1(new_n773), .A2(new_n372), .A3(new_n655), .ZN(new_n780));
  AOI21_X1  g579(.A(G120gat), .B1(new_n777), .B2(new_n613), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(G1341gat));
  NOR3_X1   g581(.A1(new_n773), .A2(new_n370), .A3(new_n554), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n777), .A2(new_n586), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(G127gat), .B1(new_n784), .B2(new_n785), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(G1342gat));
  OAI21_X1  g587(.A(G134gat), .B1(new_n773), .B2(new_n585), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n582), .A2(new_n358), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT115), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(G134gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n776), .A3(new_n792), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n793), .A2(KEYINPUT56), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(KEYINPUT56), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n789), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT116), .ZN(G1343gat));
  NOR2_X1   g596(.A1(new_n673), .A2(new_n443), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n775), .A3(new_n358), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n799), .A2(G141gat), .A3(new_n525), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(KEYINPUT58), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n217), .A2(new_n219), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n456), .A2(new_n772), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n769), .A2(new_n770), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT57), .B1(new_n804), .B2(new_n298), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n443), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n761), .A2(new_n585), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT117), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n767), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n809), .A2(KEYINPUT117), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n554), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n808), .B1(new_n813), .B2(new_n770), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n526), .B(new_n803), .C1(new_n805), .C2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n802), .B1(new_n816), .B2(KEYINPUT119), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n801), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n815), .A2(KEYINPUT118), .A3(new_n802), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT118), .B1(new_n815), .B2(new_n802), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n821), .A2(new_n822), .A3(new_n800), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(G1344gat));
  OAI21_X1  g624(.A(KEYINPUT59), .B1(new_n799), .B2(new_n706), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n222), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n586), .B1(new_n765), .B2(new_n767), .ZN(new_n828));
  INV_X1    g627(.A(new_n770), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n807), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n809), .A2(new_n767), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n829), .B1(new_n831), .B2(new_n554), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n806), .B1(new_n832), .B2(new_n443), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n613), .A3(new_n803), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n805), .A2(new_n814), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n803), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n706), .A2(KEYINPUT59), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n827), .B(new_n836), .C1(new_n838), .C2(new_n839), .ZN(G1345gat));
  OAI21_X1  g639(.A(G155gat), .B1(new_n838), .B2(new_n554), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n586), .A2(new_n207), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n799), .B2(new_n842), .ZN(G1346gat));
  NOR2_X1   g642(.A1(new_n791), .A2(G162gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n798), .A2(new_n775), .A3(new_n844), .ZN(new_n845));
  XOR2_X1   g644(.A(new_n845), .B(KEYINPUT120), .Z(new_n846));
  NAND3_X1  g645(.A1(new_n837), .A2(new_n582), .A3(new_n803), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n846), .B1(new_n848), .B2(new_n208), .ZN(G1347gat));
  OAI21_X1  g648(.A(new_n408), .B1(new_n828), .B2(new_n829), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n776), .A2(new_n618), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(G169gat), .B1(new_n852), .B2(new_n526), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n457), .A2(new_n358), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n771), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n526), .A2(G169gat), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(G1348gat));
  OAI21_X1  g657(.A(G176gat), .B1(new_n855), .B2(new_n655), .ZN(new_n859));
  INV_X1    g658(.A(G176gat), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n852), .A2(new_n860), .A3(new_n613), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1349gat));
  NAND3_X1  g661(.A1(new_n771), .A2(new_n586), .A3(new_n854), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT121), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n771), .A2(new_n865), .A3(new_n586), .A4(new_n854), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(G183gat), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n586), .A2(new_n303), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n852), .A2(new_n870), .B1(KEYINPUT122), .B2(KEYINPUT60), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n867), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n869), .B1(new_n867), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(G1350gat));
  NAND3_X1  g673(.A1(new_n852), .A2(new_n304), .A3(new_n582), .ZN(new_n875));
  OAI21_X1  g674(.A(G190gat), .B1(new_n855), .B2(new_n585), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n876), .A2(KEYINPUT61), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(KEYINPUT61), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(G1351gat));
  NAND4_X1  g678(.A1(new_n630), .A2(new_n618), .A3(new_n298), .A4(new_n631), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(KEYINPUT123), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n850), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(KEYINPUT123), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(G197gat), .B1(new_n884), .B2(new_n526), .ZN(new_n885));
  INV_X1    g684(.A(new_n834), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n632), .A2(new_n854), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n526), .A2(G197gat), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(G1352gat));
  NOR3_X1   g689(.A1(new_n886), .A2(new_n655), .A3(new_n887), .ZN(new_n891));
  INV_X1    g690(.A(G204gat), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n884), .A2(new_n892), .A3(new_n613), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(KEYINPUT62), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(KEYINPUT62), .B2(new_n894), .ZN(G1353gat));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT63), .ZN(new_n898));
  AOI211_X1 g697(.A(new_n554), .B(new_n887), .C1(new_n830), .C2(new_n833), .ZN(new_n899));
  INV_X1    g698(.A(G211gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n834), .A2(new_n586), .A3(new_n632), .A4(new_n854), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n901), .A2(KEYINPUT125), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n554), .A2(new_n232), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n882), .A2(new_n883), .A3(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n882), .A2(KEYINPUT124), .A3(new_n883), .A4(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n911), .B(new_n898), .C1(new_n899), .C2(new_n900), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n897), .B1(new_n904), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n901), .A2(new_n903), .A3(KEYINPUT125), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n915), .A2(KEYINPUT126), .A3(new_n912), .A4(new_n910), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1354gat));
  NAND3_X1  g716(.A1(new_n884), .A2(new_n237), .A3(new_n582), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n886), .A2(new_n585), .A3(new_n887), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n237), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n920), .B(new_n921), .ZN(G1355gat));
endmodule


