//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  INV_X1    g004(.A(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n205), .A2(new_n206), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT23), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(KEYINPUT25), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(KEYINPUT24), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G190gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT24), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  XOR2_X1   g018(.A(new_n219), .B(KEYINPUT66), .Z(new_n220));
  AOI21_X1  g019(.A(new_n212), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(G169gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(KEYINPUT23), .A3(new_n206), .ZN(new_n224));
  INV_X1    g023(.A(new_n218), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n219), .B(KEYINPUT64), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n210), .B(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n221), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n207), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(new_n208), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n216), .B1(new_n207), .B2(new_n229), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT28), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT27), .B(G183gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(KEYINPUT67), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT67), .B1(new_n213), .B2(KEYINPUT27), .ZN(new_n236));
  INV_X1    g035(.A(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n233), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n234), .A2(KEYINPUT28), .A3(new_n237), .ZN(new_n240));
  AOI211_X1 g039(.A(new_n231), .B(new_n232), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n228), .A2(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(G113gat), .B(G120gat), .Z(new_n243));
  XOR2_X1   g042(.A(KEYINPUT70), .B(KEYINPUT1), .Z(new_n244));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G134gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n253), .A2(KEYINPUT69), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(KEYINPUT69), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n246), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n242), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n228), .A2(new_n241), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n255), .ZN(new_n259));
  INV_X1    g058(.A(new_n246), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n257), .A2(G227gat), .A3(G233gat), .A4(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n204), .B1(new_n263), .B2(KEYINPUT32), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT33), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n265), .B1(new_n263), .B2(new_n266), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n204), .A2(new_n266), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n263), .A2(KEYINPUT32), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n263), .A2(KEYINPUT72), .A3(KEYINPUT32), .A4(new_n270), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n262), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT34), .ZN(new_n277));
  NAND2_X1  g076(.A1(G227gat), .A2(G233gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n277), .B1(new_n276), .B2(new_n278), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT73), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n269), .A2(new_n275), .A3(new_n282), .ZN(new_n283));
  OR3_X1    g082(.A1(new_n280), .A2(KEYINPUT73), .A3(new_n281), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n284), .A2(new_n275), .A3(new_n282), .A4(new_n269), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n286), .A2(KEYINPUT36), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT36), .B1(new_n286), .B2(new_n287), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G211gat), .A2(G218gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(G197gat), .A2(G204gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(G197gat), .A2(G204gat), .ZN(new_n294));
  OAI22_X1  g093(.A1(new_n292), .A2(KEYINPUT22), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n295), .A2(KEYINPUT74), .ZN(new_n296));
  NOR2_X1   g095(.A1(G211gat), .A2(G218gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n296), .B(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT29), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n258), .A2(KEYINPUT75), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n258), .A2(KEYINPUT75), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n242), .A2(new_n300), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n299), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n299), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n258), .A2(new_n302), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n303), .A2(new_n304), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n308), .B(new_n309), .C1(new_n310), .C2(new_n300), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G8gat), .B(G36gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(G64gat), .B(G92gat), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n313), .B(new_n314), .Z(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT76), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT30), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n307), .A2(new_n311), .A3(new_n319), .A4(new_n315), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n317), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n315), .B1(new_n307), .B2(new_n311), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n312), .A2(new_n316), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n322), .B1(new_n323), .B2(KEYINPUT30), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT81), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT79), .ZN(new_n327));
  XOR2_X1   g126(.A(G155gat), .B(G162gat), .Z(new_n328));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n329));
  XOR2_X1   g128(.A(G141gat), .B(G148gat), .Z(new_n330));
  AOI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT2), .ZN(new_n332));
  INV_X1    g131(.A(G155gat), .ZN(new_n333));
  INV_X1    g132(.A(G162gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n330), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  OAI221_X1 g136(.A(new_n330), .B1(new_n332), .B2(new_n335), .C1(new_n328), .C2(new_n329), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n340));
  NAND3_X1  g139(.A1(new_n256), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n339), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n261), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n327), .B(new_n341), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n339), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n342), .A2(KEYINPUT3), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n261), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT5), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n343), .A2(KEYINPUT79), .A3(new_n340), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n345), .A2(new_n351), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n340), .B1(new_n261), .B2(new_n342), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n256), .A2(KEYINPUT4), .A3(new_n339), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n355), .A2(new_n349), .A3(new_n356), .A4(new_n350), .ZN(new_n357));
  INV_X1    g156(.A(new_n350), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n256), .A2(new_n339), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n358), .B1(new_n343), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n357), .A2(new_n360), .A3(KEYINPUT5), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G1gat), .B(G29gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT0), .ZN(new_n364));
  XNOR2_X1  g163(.A(G57gat), .B(G85gat), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n364), .B(new_n365), .Z(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT6), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n326), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n366), .B1(new_n354), .B2(new_n361), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n371), .A2(KEYINPUT6), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n354), .A2(new_n366), .A3(new_n361), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n375), .A2(new_n374), .A3(new_n376), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n325), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G78gat), .B(G106gat), .Z(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(G50gat), .ZN(new_n382));
  XOR2_X1   g181(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G228gat), .ZN(new_n385));
  INV_X1    g184(.A(G233gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT29), .B1(new_n339), .B2(new_n346), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT3), .B1(new_n299), .B2(new_n301), .ZN(new_n389));
  OAI221_X1 g188(.A(new_n387), .B1(new_n388), .B2(new_n299), .C1(new_n389), .C2(new_n339), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n299), .B1(new_n347), .B2(new_n301), .ZN(new_n391));
  INV_X1    g190(.A(new_n298), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT29), .B1(new_n392), .B2(new_n295), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n392), .B2(new_n295), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n339), .B1(new_n394), .B2(new_n346), .ZN(new_n395));
  OAI22_X1  g194(.A1(new_n391), .A2(new_n395), .B1(new_n385), .B2(new_n386), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n384), .B1(new_n398), .B2(G22gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(G22gat), .B2(new_n398), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n399), .B(KEYINPUT83), .C1(G22gat), .C2(new_n398), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G22gat), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n398), .B1(KEYINPUT84), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n397), .A2(new_n407), .A3(G22gat), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n384), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT85), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n406), .A2(KEYINPUT85), .A3(new_n384), .A4(new_n408), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n404), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n290), .B(KEYINPUT86), .C1(new_n380), .C2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT86), .ZN(new_n416));
  INV_X1    g215(.A(new_n372), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT81), .B1(new_n371), .B2(KEYINPUT6), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n375), .A2(new_n376), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT80), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n421), .A3(new_n379), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n321), .A2(new_n324), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n414), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT36), .ZN(new_n425));
  INV_X1    g224(.A(new_n281), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n279), .ZN(new_n427));
  AOI211_X1 g226(.A(KEYINPUT73), .B(new_n427), .C1(new_n269), .C2(new_n275), .ZN(new_n428));
  AND4_X1   g227(.A1(new_n284), .A2(new_n269), .A3(new_n275), .A4(new_n282), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n286), .A2(KEYINPUT36), .A3(new_n287), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n416), .B1(new_n424), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n345), .A2(new_n349), .A3(new_n353), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n358), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n343), .A2(new_n359), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n435), .B(KEYINPUT39), .C1(new_n358), .C2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT39), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n434), .A2(new_n438), .A3(new_n358), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT87), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n439), .A2(new_n440), .A3(new_n366), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n440), .B1(new_n439), .B2(new_n366), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n437), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT40), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(KEYINPUT40), .B(new_n437), .C1(new_n441), .C2(new_n442), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n325), .A2(new_n445), .A3(new_n368), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n419), .A2(KEYINPUT89), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT89), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n373), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n450), .A3(new_n420), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n309), .B1(new_n310), .B2(new_n300), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n299), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n453), .A2(KEYINPUT88), .ZN(new_n454));
  OR3_X1    g253(.A1(new_n305), .A2(new_n299), .A3(new_n306), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n455), .B1(new_n453), .B2(KEYINPUT88), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT37), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n316), .B1(new_n312), .B2(KEYINPUT37), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n458), .A2(KEYINPUT38), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n312), .A2(KEYINPUT37), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT38), .B1(new_n461), .B2(new_n458), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n460), .A2(new_n317), .A3(new_n320), .A4(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n414), .B(new_n447), .C1(new_n451), .C2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n415), .A2(new_n433), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n286), .A2(new_n287), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n414), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n467), .A2(new_n468), .A3(new_n325), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n451), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n466), .A2(new_n414), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n380), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT35), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n465), .A2(new_n475), .ZN(new_n476));
  OR2_X1    g275(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n478));
  AOI21_X1  g277(.A(G36gat), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G29gat), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n480), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n481));
  OR3_X1    g280(.A1(new_n479), .A2(KEYINPUT15), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT15), .B1(new_n479), .B2(new_n481), .ZN(new_n483));
  XNOR2_X1  g282(.A(G43gat), .B(G50gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n483), .A2(new_n484), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(KEYINPUT90), .A2(KEYINPUT17), .ZN(new_n488));
  NOR2_X1   g287(.A1(KEYINPUT90), .A2(KEYINPUT17), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT17), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n485), .A2(new_n486), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT94), .ZN(new_n496));
  NAND2_X1  g295(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(G85gat), .A3(G92gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(G85gat), .A2(G92gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(KEYINPUT92), .A3(KEYINPUT7), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G99gat), .A2(G106gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT93), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(KEYINPUT93), .A2(G99gat), .A3(G106gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(KEYINPUT8), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G85gat), .ZN(new_n507));
  INV_X1    g306(.A(G92gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n501), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(G99gat), .B(G106gat), .Z(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n511), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n498), .A2(new_n500), .B1(new_n507), .B2(new_n508), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(new_n506), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n496), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n510), .A2(new_n511), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n514), .A2(new_n513), .A3(new_n506), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(KEYINPUT94), .A3(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n495), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(G232gat), .A2(G233gat), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n520), .A2(new_n487), .B1(KEYINPUT41), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  XOR2_X1   g324(.A(G190gat), .B(G218gat), .Z(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n525), .A2(new_n526), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n523), .A2(KEYINPUT41), .ZN(new_n531));
  XNOR2_X1  g330(.A(G134gat), .B(G162gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n529), .B2(new_n528), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G71gat), .A2(G78gat), .ZN(new_n539));
  INV_X1    g338(.A(G71gat), .ZN(new_n540));
  INV_X1    g339(.A(G78gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT9), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n539), .B(new_n542), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(G57gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(G64gat), .ZN(new_n547));
  INV_X1    g346(.A(G64gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G57gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n542), .A2(new_n539), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n539), .A2(new_n544), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n545), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT21), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G231gat), .A2(G233gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G127gat), .ZN(new_n559));
  INV_X1    g358(.A(G8gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(G15gat), .B(G22gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT16), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(G1gat), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n560), .B1(new_n563), .B2(KEYINPUT91), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(G1gat), .B2(new_n561), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n565), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n555), .B2(new_n554), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n559), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(new_n333), .ZN(new_n573));
  XOR2_X1   g372(.A(G183gat), .B(G211gat), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n576), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n538), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n545), .B(new_n553), .C1(new_n512), .C2(new_n515), .ZN(new_n582));
  NAND2_X1  g381(.A1(G230gat), .A2(G233gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n517), .A2(new_n554), .A3(new_n518), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT95), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G120gat), .B(G148gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(G176gat), .B(G204gat), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n589), .B(new_n590), .Z(new_n591));
  INV_X1    g390(.A(KEYINPUT10), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n554), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n516), .A2(new_n519), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT10), .B1(new_n582), .B2(new_n585), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n583), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n588), .A2(new_n591), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT96), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n591), .B1(new_n588), .B2(new_n597), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n581), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n495), .A2(new_n569), .ZN(new_n603));
  NAND2_X1  g402(.A1(G229gat), .A2(G233gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n568), .A2(new_n487), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT18), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n603), .A2(KEYINPUT18), .A3(new_n604), .A4(new_n605), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n604), .B(KEYINPUT13), .Z(new_n610));
  INV_X1    g409(.A(new_n605), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n568), .A2(new_n487), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G113gat), .B(G141gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G197gat), .ZN(new_n616));
  XOR2_X1   g415(.A(KEYINPUT11), .B(G169gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  NAND2_X1  g418(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n608), .A2(new_n609), .A3(new_n621), .A4(new_n613), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n602), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n476), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n422), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g429(.A(new_n560), .B1(new_n627), .B2(new_n325), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT16), .B(G8gat), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n626), .A2(new_n423), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT42), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(KEYINPUT42), .B2(new_n633), .ZN(G1325gat));
  NOR3_X1   g434(.A1(new_n626), .A2(G15gat), .A3(new_n467), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n627), .A2(new_n432), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(G15gat), .B2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT97), .Z(G1326gat));
  NOR2_X1   g438(.A1(new_n626), .A2(new_n414), .ZN(new_n640));
  XOR2_X1   g439(.A(KEYINPUT43), .B(G22gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(G1327gat));
  INV_X1    g441(.A(new_n601), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n643), .A2(new_n624), .A3(new_n579), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n476), .A2(new_n538), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n646), .A2(new_n480), .A3(new_n628), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT45), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n649), .B1(new_n476), .B2(new_n538), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n537), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n534), .A2(KEYINPUT98), .A3(new_n536), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n424), .A2(new_n432), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n464), .A2(new_n656), .ZN(new_n657));
  AOI211_X1 g456(.A(KEYINPUT44), .B(new_n655), .C1(new_n475), .C2(new_n657), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n650), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n644), .ZN(new_n660));
  OAI21_X1  g459(.A(G29gat), .B1(new_n660), .B2(new_n422), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n648), .A2(new_n661), .ZN(G1328gat));
  OAI21_X1  g461(.A(G36gat), .B1(new_n660), .B2(new_n423), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n645), .A2(G36gat), .A3(new_n423), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT46), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(G1329gat));
  INV_X1    g465(.A(G43gat), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(new_n645), .B2(new_n467), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n432), .A2(G43gat), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n668), .B1(new_n660), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g470(.A(KEYINPUT48), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n645), .A2(G50gat), .A3(new_n414), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n672), .B1(new_n673), .B2(KEYINPUT100), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n468), .B(new_n644), .C1(new_n650), .C2(new_n658), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(G50gat), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n674), .B(new_n676), .C1(KEYINPUT100), .C2(new_n673), .ZN(new_n677));
  INV_X1    g476(.A(new_n673), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT99), .B1(new_n679), .B2(new_n672), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n673), .B1(new_n675), .B2(G50gat), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n681), .A2(new_n682), .A3(KEYINPUT48), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n677), .B1(new_n680), .B2(new_n683), .ZN(G1331gat));
  NAND2_X1  g483(.A1(new_n475), .A2(new_n657), .ZN(new_n685));
  NOR4_X1   g484(.A1(new_n538), .A2(new_n580), .A3(new_n623), .A4(new_n601), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n422), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT101), .B(G57gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1332gat));
  NOR2_X1   g489(.A1(new_n687), .A2(new_n423), .ZN(new_n691));
  NOR2_X1   g490(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n692));
  AND2_X1   g491(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n691), .B2(new_n692), .ZN(G1333gat));
  NOR3_X1   g494(.A1(new_n687), .A2(G71gat), .A3(new_n467), .ZN(new_n696));
  INV_X1    g495(.A(new_n687), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n432), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(G71gat), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g499(.A1(new_n687), .A2(new_n414), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(new_n541), .ZN(G1335gat));
  NAND3_X1  g501(.A1(new_n580), .A2(new_n538), .A3(new_n624), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n475), .B2(new_n657), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT51), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n628), .A2(new_n507), .A3(new_n643), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT103), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n579), .A2(new_n601), .A3(new_n623), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n659), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n711), .B2(new_n422), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G85gat), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n711), .A2(new_n709), .A3(new_n422), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n708), .B1(new_n713), .B2(new_n714), .ZN(G1336gat));
  NAND3_X1  g514(.A1(new_n659), .A2(new_n325), .A3(new_n710), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G92gat), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n423), .A2(G92gat), .A3(new_n601), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT52), .B1(new_n705), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT51), .ZN(new_n721));
  OR3_X1    g520(.A1(new_n704), .A2(KEYINPUT104), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n704), .B2(KEYINPUT104), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n722), .A2(new_n723), .A3(new_n718), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n724), .B1(new_n716), .B2(G92gat), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n720), .B1(new_n725), .B2(new_n726), .ZN(G1337gat));
  OAI21_X1  g526(.A(G99gat), .B1(new_n711), .B2(new_n290), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n467), .A2(G99gat), .A3(new_n601), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n705), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1338gat));
  NAND3_X1  g530(.A1(new_n659), .A2(new_n468), .A3(new_n710), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G106gat), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT107), .B(KEYINPUT53), .Z(new_n734));
  NOR3_X1   g533(.A1(new_n414), .A2(G106gat), .A3(new_n601), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT105), .Z(new_n736));
  AOI21_X1  g535(.A(new_n734), .B1(new_n705), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n736), .B(KEYINPUT106), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n722), .A2(new_n723), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(new_n732), .B2(G106gat), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT53), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n738), .B1(new_n741), .B2(new_n742), .ZN(G1339gat));
  NOR2_X1   g542(.A1(new_n602), .A2(new_n623), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n517), .A2(new_n554), .A3(new_n518), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n554), .B1(new_n517), .B2(new_n518), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n592), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n584), .B1(new_n747), .B2(new_n594), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT54), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n591), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n747), .A2(new_n584), .A3(new_n594), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT108), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n747), .A2(new_n754), .A3(new_n594), .A4(new_n584), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n753), .A2(KEYINPUT54), .A3(new_n597), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT109), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n748), .A2(new_n749), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n758), .A2(new_n753), .A3(new_n759), .A4(new_n755), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n751), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n599), .B1(KEYINPUT55), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n757), .A2(new_n760), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n750), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT110), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n761), .A2(new_n767), .A3(KEYINPUT55), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n623), .B(new_n762), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n604), .B1(new_n603), .B2(new_n605), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT111), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  OR3_X1    g571(.A1(new_n611), .A2(new_n612), .A3(new_n610), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n770), .B2(KEYINPUT111), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n618), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n775), .A2(new_n622), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n643), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n769), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n769), .A2(KEYINPUT112), .A3(new_n777), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n780), .A2(new_n655), .A3(new_n781), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n776), .B(new_n762), .C1(new_n766), .C2(new_n768), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n654), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n744), .B1(new_n786), .B2(new_n580), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n468), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n628), .A2(new_n423), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n467), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(G113gat), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n791), .A2(new_n792), .A3(new_n624), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n787), .A2(new_n422), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n469), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n623), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n793), .B1(new_n792), .B2(new_n797), .ZN(G1340gat));
  INV_X1    g597(.A(G120gat), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n791), .A2(new_n799), .A3(new_n601), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n796), .A2(new_n643), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n799), .B2(new_n801), .ZN(G1341gat));
  OAI21_X1  g601(.A(G127gat), .B1(new_n791), .B2(new_n580), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n580), .A2(G127gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n795), .B2(new_n804), .ZN(G1342gat));
  NAND3_X1  g604(.A1(new_n796), .A2(new_n249), .A3(new_n538), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n806), .A2(KEYINPUT56), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(KEYINPUT56), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n788), .A2(new_n538), .A3(new_n790), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n809), .A2(new_n810), .A3(G134gat), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n809), .B2(G134gat), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n807), .B(new_n808), .C1(new_n811), .C2(new_n812), .ZN(G1343gat));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n414), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n764), .A2(new_n818), .A3(new_n765), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT114), .B1(new_n761), .B2(KEYINPUT55), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n762), .A2(new_n819), .A3(new_n623), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n777), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n537), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n785), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT115), .B1(new_n824), .B2(new_n579), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n579), .B1(new_n785), .B2(new_n823), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n744), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n817), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n579), .B1(new_n782), .B2(new_n785), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n468), .B1(new_n830), .B2(new_n744), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n829), .B1(new_n815), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n789), .A2(new_n432), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n814), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n831), .A2(new_n815), .ZN(new_n836));
  OAI211_X1 g635(.A(KEYINPUT116), .B(new_n833), .C1(new_n836), .C2(new_n829), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n837), .A3(new_n623), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n432), .A2(new_n325), .A3(new_n414), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n794), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n624), .A2(G141gat), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n838), .A2(G141gat), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n794), .A2(new_n839), .A3(new_n842), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n844), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n623), .B(new_n833), .C1(new_n836), .C2(new_n829), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(G141gat), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(KEYINPUT117), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850));
  AOI211_X1 g649(.A(new_n850), .B(new_n846), .C1(new_n847), .C2(G141gat), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n843), .A2(new_n844), .B1(new_n849), .B2(new_n851), .ZN(G1344gat));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853));
  AOI211_X1 g652(.A(new_n853), .B(G148gat), .C1(new_n841), .C2(new_n643), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n835), .A2(new_n837), .A3(new_n643), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n853), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT119), .B1(new_n787), .B2(new_n817), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n858), .B(new_n816), .C1(new_n830), .C2(new_n744), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n823), .B1(new_n537), .B2(new_n783), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n744), .B1(new_n860), .B2(new_n580), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n815), .B1(new_n861), .B2(new_n414), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n857), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n833), .A2(KEYINPUT118), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n833), .A2(KEYINPUT118), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n601), .A2(new_n853), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n856), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n854), .B1(new_n868), .B2(G148gat), .ZN(G1345gat));
  NAND3_X1  g668(.A1(new_n841), .A2(new_n333), .A3(new_n579), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n835), .A2(new_n837), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(new_n579), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n872), .B2(new_n333), .ZN(G1346gat));
  AOI21_X1  g672(.A(G162gat), .B1(new_n841), .B2(new_n538), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n655), .A2(new_n334), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n871), .B2(new_n875), .ZN(G1347gat));
  NOR3_X1   g675(.A1(new_n628), .A2(new_n423), .A3(new_n467), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n788), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G169gat), .B1(new_n878), .B2(new_n624), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n787), .A2(new_n628), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n472), .A2(new_n325), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n623), .A2(new_n223), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n883), .B2(new_n884), .ZN(G1348gat));
  OAI21_X1  g684(.A(G176gat), .B1(new_n878), .B2(new_n601), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n643), .A2(new_n206), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT120), .ZN(G1349gat));
  OAI21_X1  g688(.A(G183gat), .B1(new_n878), .B2(new_n580), .ZN(new_n890));
  AND4_X1   g689(.A1(new_n234), .A2(new_n880), .A3(new_n579), .A4(new_n882), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(KEYINPUT121), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(KEYINPUT121), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(KEYINPUT60), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT60), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n896), .B(new_n890), .C1(new_n892), .C2(new_n893), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1350gat));
  NAND3_X1  g697(.A1(new_n788), .A2(new_n538), .A3(new_n877), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n899), .A2(new_n900), .A3(G190gat), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n899), .B2(G190gat), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n654), .A2(new_n237), .ZN(new_n903));
  OAI22_X1  g702(.A1(new_n901), .A2(new_n902), .B1(new_n883), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n904), .B(new_n905), .ZN(G1351gat));
  NOR3_X1   g705(.A1(new_n432), .A2(new_n423), .A3(new_n414), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n880), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n908), .A2(KEYINPUT123), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(KEYINPUT123), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g710(.A(KEYINPUT124), .B(G197gat), .Z(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n623), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n290), .A2(new_n422), .A3(new_n325), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT125), .Z(new_n915));
  AND2_X1   g714(.A1(new_n863), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n916), .A2(new_n623), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n917), .B2(new_n912), .ZN(G1352gat));
  NOR3_X1   g717(.A1(new_n908), .A2(G204gat), .A3(new_n601), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT62), .ZN(new_n920));
  INV_X1    g719(.A(G204gat), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n916), .A2(new_n643), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(G1353gat));
  INV_X1    g722(.A(G211gat), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n924), .A3(new_n579), .A4(new_n910), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n914), .A2(new_n580), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n863), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT63), .B1(new_n927), .B2(G211gat), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT63), .ZN(new_n929));
  AOI211_X1 g728(.A(new_n929), .B(new_n924), .C1(new_n863), .C2(new_n926), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n925), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT126), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n925), .B(new_n933), .C1(new_n928), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1354gat));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n916), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n538), .B1(new_n916), .B2(new_n936), .ZN(new_n938));
  OAI21_X1  g737(.A(G218gat), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(G218gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n911), .A2(new_n940), .A3(new_n654), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1355gat));
endmodule


