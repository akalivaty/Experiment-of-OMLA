//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT67), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G953), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G237), .ZN(new_n193));
  AND4_X1   g007(.A1(G143), .A2(new_n192), .A3(G214), .A4(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(G237), .B1(new_n189), .B2(new_n191), .ZN(new_n195));
  AOI21_X1  g009(.A(G143), .B1(new_n195), .B2(G214), .ZN(new_n196));
  OAI21_X1  g010(.A(G131), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT89), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n192), .A2(G214), .A3(new_n193), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n195), .A2(G143), .A3(G214), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT89), .A3(G131), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n199), .A2(KEYINPUT17), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT91), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G125), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G140), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT74), .A4(KEYINPUT16), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT16), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n211), .B2(KEYINPUT16), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n209), .B(new_n214), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT16), .ZN(new_n220));
  OR3_X1    g034(.A1(new_n212), .A2(KEYINPUT16), .A3(G140), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(new_n216), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n209), .B1(new_n222), .B2(new_n214), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n204), .ZN(new_n225));
  INV_X1    g039(.A(G131), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT17), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT89), .B1(new_n204), .B2(G131), .ZN(new_n229));
  AOI211_X1 g043(.A(new_n198), .B(new_n226), .C1(new_n202), .C2(new_n203), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n227), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n199), .A2(new_n205), .A3(KEYINPUT91), .A4(KEYINPUT17), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n208), .A2(new_n224), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G113), .B(G122), .ZN(new_n234));
  INV_X1    g048(.A(G104), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT18), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n225), .B1(new_n237), .B2(new_n226), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n204), .A2(KEYINPUT18), .A3(G131), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n211), .A2(new_n213), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n209), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT88), .B1(new_n240), .B2(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(KEYINPUT88), .A3(G146), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n238), .A2(new_n239), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n233), .A2(new_n236), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n236), .B1(new_n233), .B2(new_n246), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n187), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT92), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(KEYINPUT92), .B(new_n187), .C1(new_n247), .C2(new_n248), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(G475), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n233), .A2(new_n236), .A3(new_n246), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n199), .A2(new_n205), .B1(new_n226), .B2(new_n225), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n214), .B1(new_n215), .B2(new_n217), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n241), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n241), .B2(new_n258), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n257), .B1(new_n261), .B2(G146), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n246), .B1(new_n255), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n236), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n254), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G475), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(new_n187), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT20), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT20), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n266), .A2(new_n270), .A3(new_n267), .A4(new_n187), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g086(.A(KEYINPUT9), .B(G234), .Z(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(G217), .A3(new_n188), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n201), .A2(G128), .ZN(new_n276));
  INV_X1    g090(.A(G128), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G143), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(G134), .ZN(new_n280));
  INV_X1    g094(.A(G122), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G116), .ZN(new_n282));
  INV_X1    g096(.A(G116), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n283), .A2(KEYINPUT93), .A3(G122), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT93), .B1(new_n283), .B2(G122), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G107), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT93), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(new_n281), .B2(G116), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n283), .A2(KEYINPUT93), .A3(G122), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G107), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n282), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n280), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n276), .A2(new_n278), .A3(KEYINPUT13), .ZN(new_n295));
  OR3_X1    g109(.A1(new_n277), .A2(KEYINPUT13), .A3(G143), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(G134), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT94), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT94), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n295), .A2(new_n296), .A3(new_n299), .A4(G134), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT95), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n294), .A2(new_n301), .A3(KEYINPUT95), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n279), .B(G134), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT96), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n291), .B2(KEYINPUT14), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT14), .ZN(new_n310));
  AOI211_X1 g124(.A(KEYINPUT96), .B(new_n310), .C1(new_n289), .C2(new_n290), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n289), .A2(new_n310), .A3(new_n290), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n282), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n309), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n307), .B(new_n293), .C1(new_n314), .C2(new_n292), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n275), .B1(new_n306), .B2(new_n315), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n294), .A2(new_n301), .A3(KEYINPUT95), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT95), .B1(new_n294), .B2(new_n301), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n315), .B(new_n275), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n187), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT97), .ZN(new_n322));
  INV_X1    g136(.A(G478), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(KEYINPUT15), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n274), .ZN(new_n326));
  AOI21_X1  g140(.A(G902), .B1(new_n326), .B2(new_n319), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT97), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n322), .A2(new_n324), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n327), .B1(KEYINPUT15), .B2(new_n323), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n188), .A2(G952), .ZN(new_n334));
  INV_X1    g148(.A(G234), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(new_n193), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  AOI211_X1 g151(.A(new_n187), .B(new_n192), .C1(G234), .C2(G237), .ZN(new_n338));
  XOR2_X1   g152(.A(KEYINPUT21), .B(G898), .Z(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n337), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n253), .A2(new_n272), .A3(new_n333), .A4(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(KEYINPUT78), .A2(G104), .ZN(new_n344));
  NOR2_X1   g158(.A1(KEYINPUT78), .A2(G104), .ZN(new_n345));
  OAI21_X1  g159(.A(G107), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n292), .A3(G104), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n344), .A2(new_n345), .A3(G107), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n346), .B(new_n348), .C1(new_n349), .C2(new_n347), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G101), .ZN(new_n351));
  OR2_X1    g165(.A1(KEYINPUT78), .A2(G104), .ZN(new_n352));
  NAND2_X1  g166(.A1(KEYINPUT78), .A2(G104), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n292), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT3), .ZN(new_n355));
  INV_X1    g169(.A(G101), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n355), .A2(new_n356), .A3(new_n346), .A4(new_n348), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n351), .A2(KEYINPUT4), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(KEYINPUT2), .A2(G113), .ZN(new_n359));
  NAND2_X1  g173(.A1(KEYINPUT2), .A2(G113), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT66), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT66), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT2), .A3(G113), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n359), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G116), .B(G119), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n364), .B(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n350), .A2(new_n369), .A3(G101), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n358), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n283), .A2(KEYINPUT5), .A3(G119), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(new_n365), .B2(KEYINPUT5), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G113), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n364), .A2(new_n365), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n292), .A2(G104), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n344), .A2(new_n345), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n377), .B1(new_n378), .B2(new_n292), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT79), .B1(new_n379), .B2(new_n356), .ZN(new_n380));
  INV_X1    g194(.A(new_n377), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n356), .B1(new_n354), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT79), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n376), .A2(new_n380), .A3(new_n357), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n371), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G110), .B(G122), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n371), .A2(new_n385), .A3(new_n387), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(KEYINPUT6), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(KEYINPUT0), .A2(G128), .ZN(new_n392));
  XNOR2_X1  g206(.A(G143), .B(G146), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n392), .B1(new_n393), .B2(KEYINPUT64), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n201), .A2(G146), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n209), .A2(G143), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT0), .B(G128), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT64), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G125), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n277), .A2(new_n209), .A3(G143), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n201), .B(G146), .C1(new_n277), .C2(KEYINPUT1), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n277), .A2(KEYINPUT1), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n403), .B(new_n404), .C1(new_n397), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n212), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT83), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n402), .A2(new_n410), .A3(new_n407), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G224), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(G953), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n409), .A2(G224), .A3(new_n188), .A4(new_n411), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n386), .A2(new_n417), .A3(new_n388), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n391), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT84), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT84), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n391), .A2(new_n416), .A3(new_n421), .A4(new_n418), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n406), .A2(new_n212), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n212), .B1(new_n394), .B2(new_n400), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT85), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT7), .B1(new_n413), .B2(G953), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  OAI22_X1  g242(.A1(new_n424), .A2(new_n425), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(KEYINPUT85), .B2(new_n427), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n408), .A2(new_n426), .A3(new_n428), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n387), .B(KEYINPUT8), .Z(new_n433));
  NAND3_X1  g247(.A1(new_n380), .A2(new_n384), .A3(new_n357), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n374), .A2(new_n375), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n433), .B1(new_n385), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n432), .A2(new_n438), .A3(KEYINPUT86), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT86), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n430), .A2(new_n431), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n440), .B1(new_n441), .B2(new_n437), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n442), .A3(new_n390), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n187), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n423), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G210), .B1(G237), .B2(G902), .ZN(new_n447));
  XOR2_X1   g261(.A(new_n447), .B(KEYINPUT87), .Z(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G214), .B1(G237), .B2(G902), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n423), .A2(new_n448), .A3(new_n445), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n343), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n192), .A2(G210), .A3(new_n193), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(G101), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G134), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT11), .B1(new_n460), .B2(G137), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT11), .ZN(new_n462));
  INV_X1    g276(.A(G137), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n463), .A3(G134), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n463), .A2(G134), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n226), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  AOI211_X1 g282(.A(G131), .B(new_n466), .C1(new_n461), .C2(new_n464), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n401), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT65), .B1(new_n463), .B2(G134), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT65), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n460), .A3(G137), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n463), .A2(G134), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G131), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n465), .A2(new_n226), .A3(new_n467), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n406), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n470), .A2(new_n367), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n367), .B1(new_n470), .B2(new_n478), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT28), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n470), .A2(new_n367), .A3(new_n478), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT28), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT69), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT69), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n462), .B1(G134), .B2(new_n463), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n460), .A2(KEYINPUT11), .A3(G137), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n467), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G131), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n490), .A2(new_n477), .B1(new_n400), .B2(new_n394), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n406), .A2(new_n476), .A3(new_n477), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n368), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n482), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n486), .B1(new_n494), .B2(KEYINPUT28), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n459), .B1(new_n485), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n491), .B2(new_n492), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n470), .A2(KEYINPUT30), .A3(new_n478), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n368), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n482), .A3(new_n458), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT31), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT68), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT31), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n500), .A2(new_n458), .A3(new_n504), .A4(new_n482), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT68), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n501), .A2(new_n506), .A3(KEYINPUT31), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n496), .A2(new_n503), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(G472), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n187), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT70), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT71), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT32), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n458), .B1(new_n485), .B2(new_n495), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n500), .A2(new_n482), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(new_n458), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT29), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n481), .A2(new_n484), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(KEYINPUT29), .A3(new_n458), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n187), .ZN(new_n522));
  OAI21_X1  g336(.A(G472), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT71), .B1(new_n510), .B2(new_n511), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT32), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n510), .B2(KEYINPUT71), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n514), .B(new_n523), .C1(new_n524), .C2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT76), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT23), .B1(new_n277), .B2(G119), .ZN(new_n529));
  INV_X1    g343(.A(G119), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n529), .B(KEYINPUT73), .C1(new_n530), .C2(G128), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT73), .B1(new_n530), .B2(G128), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n532), .B(KEYINPUT23), .C1(G119), .C2(new_n277), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G110), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n530), .A2(KEYINPUT72), .A3(G128), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT72), .B1(new_n530), .B2(G128), .ZN(new_n537));
  OAI22_X1  g351(.A1(new_n536), .A2(new_n537), .B1(new_n530), .B2(G128), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT24), .B(G110), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n535), .B(new_n540), .C1(new_n219), .C2(new_n223), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n538), .A2(new_n539), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n534), .B2(G110), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n257), .A3(new_n242), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT22), .B(G137), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n545), .B(new_n546), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n541), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n547), .B1(new_n541), .B2(new_n544), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n548), .A2(new_n549), .A3(G902), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n528), .B1(new_n550), .B2(KEYINPUT75), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n541), .A2(new_n544), .ZN(new_n552));
  INV_X1    g366(.A(new_n547), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n541), .A2(new_n544), .A3(new_n547), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n187), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT76), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n551), .A2(KEYINPUT25), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G217), .B1(new_n335), .B2(G902), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT75), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT76), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT25), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n548), .A2(new_n549), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n559), .A2(new_n187), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT82), .B(G469), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n406), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n434), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n380), .A2(new_n384), .A3(new_n357), .A4(new_n406), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n469), .A2(new_n468), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT81), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT12), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n578), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n575), .A2(new_n579), .A3(new_n580), .A4(new_n577), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT80), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n574), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT10), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n358), .A2(new_n401), .A3(new_n370), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n574), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n587), .A2(new_n576), .A3(new_n588), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n192), .A2(G227), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT77), .ZN(new_n593));
  XNOR2_X1  g407(.A(G110), .B(G140), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n583), .A2(new_n584), .A3(new_n591), .A4(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n577), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n595), .B1(new_n599), .B2(new_n591), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n187), .B(new_n571), .C1(new_n597), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(G469), .A2(G902), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n583), .A2(new_n584), .A3(new_n591), .ZN(new_n603));
  INV_X1    g417(.A(new_n595), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n599), .A2(new_n591), .A3(new_n595), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(G469), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n601), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n273), .ZN(new_n609));
  OAI21_X1  g423(.A(G221), .B1(new_n609), .B2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n454), .A2(new_n527), .A3(new_n569), .A4(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  NAND2_X1  g428(.A1(new_n508), .A2(new_n187), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(KEYINPUT98), .A2(G472), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n615), .A2(KEYINPUT98), .A3(G472), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n620), .A2(new_n611), .A3(new_n568), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n253), .A2(new_n272), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n322), .A2(new_n323), .A3(new_n329), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(new_n316), .B2(new_n320), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n326), .A2(KEYINPUT33), .A3(new_n319), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n625), .A2(G478), .A3(new_n187), .A4(new_n626), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n453), .A2(new_n341), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n621), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  NAND2_X1  g447(.A1(new_n253), .A2(new_n272), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n333), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n621), .A2(new_n630), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  NOR2_X1   g452(.A1(new_n553), .A2(KEYINPUT36), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n552), .B(new_n639), .Z(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n567), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n558), .B2(new_n563), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n343), .A2(new_n642), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n423), .A2(new_n448), .A3(new_n445), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n448), .B1(new_n423), .B2(new_n445), .ZN(new_n645));
  INV_X1    g459(.A(new_n451), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n620), .A2(new_n611), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n643), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT37), .B(G110), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  INV_X1    g465(.A(new_n642), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n527), .A2(new_n612), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n338), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(G900), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n655), .A2(KEYINPUT99), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(KEYINPUT99), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n336), .A3(new_n657), .ZN(new_n658));
  AND4_X1   g472(.A1(new_n253), .A2(new_n272), .A3(new_n332), .A4(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n647), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n253), .A2(new_n272), .A3(new_n332), .A4(new_n658), .ZN(new_n662));
  OAI21_X1  g476(.A(KEYINPUT100), .B1(new_n662), .B2(new_n453), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n653), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT101), .B(G128), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G30));
  NOR2_X1   g481(.A1(new_n644), .A2(new_n645), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT38), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n646), .B1(new_n253), .B2(new_n272), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n670), .A2(new_n332), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n658), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n612), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT40), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n669), .A2(new_n671), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n459), .A2(new_n494), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(G472), .A3(new_n501), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n509), .A2(new_n187), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n681), .B(KEYINPUT102), .Z(new_n682));
  OAI211_X1 g496(.A(new_n514), .B(new_n682), .C1(new_n524), .C2(new_n526), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n683), .A2(new_n642), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n676), .B(new_n684), .C1(KEYINPUT40), .C2(new_n674), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G143), .ZN(G45));
  INV_X1    g500(.A(new_n628), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n634), .A2(new_n687), .A3(new_n658), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n453), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n527), .A3(new_n612), .A4(new_n652), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  AND4_X1   g505(.A1(new_n647), .A2(new_n634), .A3(new_n342), .A4(new_n687), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n599), .A2(new_n591), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n604), .ZN(new_n694));
  AOI21_X1  g508(.A(G902), .B1(new_n694), .B2(new_n596), .ZN(new_n695));
  INV_X1    g509(.A(G469), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n601), .B(new_n610), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n692), .A2(new_n569), .A3(new_n527), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  NOR4_X1   g515(.A1(new_n453), .A2(new_n634), .A3(new_n333), .A4(new_n341), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n702), .A2(new_n569), .A3(new_n527), .A4(new_n698), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  NOR2_X1   g518(.A1(new_n453), .A2(new_n697), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n643), .A2(new_n705), .A3(new_n527), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G119), .ZN(G21));
  XOR2_X1   g521(.A(KEYINPUT104), .B(G472), .Z(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n508), .B2(new_n187), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n502), .B(new_n505), .C1(new_n520), .C2(new_n458), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n509), .A3(new_n187), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n713), .A2(new_n568), .A3(new_n341), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n671), .A2(new_n668), .A3(new_n698), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  INV_X1    g530(.A(new_n658), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n717), .B(new_n628), .C1(new_n253), .C2(new_n272), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n709), .A2(new_n642), .A3(new_n712), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n705), .A2(new_n718), .A3(KEYINPUT105), .A4(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n634), .A2(new_n719), .A3(new_n687), .A4(new_n658), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n698), .A2(new_n451), .A3(new_n452), .A4(new_n450), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT106), .B(G125), .Z(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G27));
  XNOR2_X1  g541(.A(new_n602), .B(KEYINPUT107), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n601), .A2(new_n607), .A3(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(new_n730), .B(KEYINPUT108), .Z(new_n731));
  INV_X1    g545(.A(new_n610), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n646), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n668), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n527), .A2(new_n569), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n688), .A2(KEYINPUT42), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n510), .A2(new_n525), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n510), .A2(new_n525), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n523), .A3(new_n742), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n743), .A2(new_n569), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n718), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT42), .B1(new_n745), .B2(new_n736), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G131), .ZN(G33));
  NAND3_X1  g562(.A1(new_n737), .A2(new_n738), .A3(new_n659), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  NAND2_X1  g564(.A1(new_n622), .A2(KEYINPUT111), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n634), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n751), .A2(KEYINPUT43), .A3(new_n687), .A4(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n755));
  OAI211_X1 g569(.A(KEYINPUT110), .B(new_n755), .C1(new_n634), .C2(new_n628), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n755), .B1(new_n634), .B2(new_n628), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n754), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n620), .A3(new_n652), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT44), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n668), .A2(new_n646), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n605), .A2(new_n606), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n605), .A2(KEYINPUT45), .A3(new_n606), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(G469), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n769), .A2(new_n729), .B1(new_n770), .B2(KEYINPUT46), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(KEYINPUT46), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n771), .A2(new_n772), .B1(new_n695), .B2(new_n571), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n732), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n775), .A2(new_n673), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n764), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  INV_X1    g592(.A(new_n763), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n779), .A2(new_n527), .A3(new_n688), .A4(new_n569), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT113), .ZN(new_n781));
  XNOR2_X1  g595(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n775), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n775), .A2(new_n782), .ZN(new_n784));
  OR3_X1    g598(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  NOR2_X1   g600(.A1(new_n683), .A2(new_n568), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n601), .B1(new_n695), .B2(new_n696), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(KEYINPUT49), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n751), .A2(new_n687), .A3(new_n753), .ZN(new_n790));
  INV_X1    g604(.A(new_n788), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT49), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n733), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OR4_X1    g607(.A1(new_n669), .A2(new_n789), .A3(new_n790), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n713), .A2(new_n568), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n760), .A2(new_n646), .A3(new_n337), .A4(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n797), .A2(new_n669), .A3(new_n697), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OAI22_X1  g614(.A1(new_n783), .A2(new_n784), .B1(new_n610), .B2(new_n788), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n760), .A2(new_n337), .A3(new_n796), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n763), .A3(new_n802), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n668), .A2(new_n336), .A3(new_n788), .A4(new_n734), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n787), .A2(new_n622), .A3(new_n628), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n760), .A2(new_n719), .A3(new_n804), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n803), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n795), .B1(new_n800), .B2(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n803), .A2(new_n805), .A3(new_n806), .ZN(new_n809));
  INV_X1    g623(.A(new_n669), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n802), .A2(new_n646), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n799), .B1(new_n811), .B2(new_n697), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n798), .A2(KEYINPUT50), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n809), .A2(KEYINPUT51), .A3(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n808), .A2(new_n334), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n760), .A2(new_n744), .A3(new_n804), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT119), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT48), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n802), .A2(new_n705), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n787), .A2(new_n629), .A3(new_n804), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n816), .A2(new_n819), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n653), .A2(new_n689), .B1(new_n720), .B2(new_n724), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n658), .B(KEYINPUT116), .Z(new_n826));
  AND4_X1   g640(.A1(new_n668), .A2(new_n670), .A3(new_n332), .A4(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n684), .A2(new_n610), .A3(new_n731), .A4(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n824), .A2(new_n825), .A3(new_n665), .A4(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n829), .A2(new_n747), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n699), .A2(new_n703), .A3(new_n706), .A4(new_n715), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n828), .A2(new_n665), .A3(new_n690), .A4(new_n725), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n831), .B1(new_n832), .B2(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n653), .A2(new_n763), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n622), .A2(new_n333), .A3(new_n658), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n749), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n613), .A2(new_n649), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(KEYINPUT114), .A3(new_n631), .A4(new_n636), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n613), .A2(new_n631), .A3(new_n636), .A4(new_n649), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n836), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n736), .A2(new_n722), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT115), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n830), .A2(new_n833), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n845), .A2(KEYINPUT53), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(KEYINPUT53), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n833), .A2(KEYINPUT117), .A3(new_n747), .A4(new_n829), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT53), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(new_n845), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n823), .B(new_n848), .C1(new_n851), .C2(KEYINPUT54), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n846), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n830), .A2(new_n833), .A3(new_n844), .A4(new_n842), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n850), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n845), .A2(KEYINPUT53), .A3(new_n849), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT54), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT118), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n822), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(G952), .A2(G953), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n794), .B1(new_n859), .B2(new_n860), .ZN(G75));
  NAND4_X1  g675(.A1(new_n855), .A2(G902), .A3(new_n856), .A4(new_n448), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n391), .A2(new_n418), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(new_n416), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT55), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT56), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n864), .A2(new_n867), .B1(new_n868), .B2(new_n862), .ZN(new_n869));
  AND4_X1   g683(.A1(KEYINPUT120), .A2(new_n862), .A3(new_n868), .A4(new_n867), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n192), .A2(G952), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(G51));
  NAND2_X1  g686(.A1(new_n729), .A2(KEYINPUT57), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n729), .A2(KEYINPUT57), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n855), .A2(KEYINPUT54), .A3(new_n856), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n873), .B(new_n874), .C1(new_n875), .C2(new_n857), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n600), .B2(new_n597), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n851), .A2(G902), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(G469), .A3(new_n767), .A4(new_n768), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n871), .B1(new_n877), .B2(new_n879), .ZN(G54));
  NAND4_X1  g694(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .A4(new_n266), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n851), .A2(KEYINPUT58), .A3(G902), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n254), .B(new_n265), .C1(new_n882), .C2(new_n267), .ZN(new_n883));
  INV_X1    g697(.A(new_n871), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n881), .A2(new_n883), .A3(new_n884), .ZN(G60));
  NAND2_X1  g699(.A1(G478), .A2(G902), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT59), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n875), .B2(new_n857), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n625), .A2(new_n626), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n884), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n858), .A2(new_n852), .A3(new_n887), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n892), .B2(new_n890), .ZN(G63));
  NAND2_X1  g707(.A1(G217), .A2(G902), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT60), .Z(new_n895));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n640), .B2(KEYINPUT122), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n640), .A2(KEYINPUT122), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n851), .A2(new_n895), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n855), .A2(new_n856), .A3(new_n895), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n871), .B1(new_n900), .B2(new_n566), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n901), .B2(new_n896), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT61), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n899), .B(new_n904), .C1(new_n901), .C2(new_n896), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n903), .A2(new_n905), .ZN(G66));
  OAI21_X1  g720(.A(G953), .B1(new_n340), .B2(new_n413), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n838), .A2(new_n841), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n831), .ZN(new_n910));
  INV_X1    g724(.A(new_n192), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n865), .B1(G898), .B2(new_n192), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(G69));
  NAND3_X1  g728(.A1(new_n685), .A2(new_n665), .A3(new_n824), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT62), .Z(new_n916));
  OAI21_X1  g730(.A(new_n738), .B1(new_n629), .B2(new_n635), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n917), .A2(new_n674), .A3(new_n779), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT124), .Z(new_n919));
  NAND4_X1  g733(.A1(new_n916), .A2(new_n777), .A3(new_n785), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n192), .ZN(new_n921));
  NAND2_X1  g735(.A1(G227), .A2(G900), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n911), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n498), .A2(new_n499), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT123), .Z(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(new_n261), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n921), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  XOR2_X1   g741(.A(KEYINPUT125), .B(G900), .Z(new_n928));
  NOR2_X1   g742(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  AND4_X1   g743(.A1(new_n665), .A2(new_n785), .A3(new_n749), .A4(new_n824), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n744), .A2(new_n671), .A3(new_n668), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n776), .B1(new_n764), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n930), .A2(new_n932), .A3(new_n747), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n929), .B1(new_n933), .B2(new_n192), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n927), .B1(new_n934), .B2(new_n926), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT126), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n927), .B(new_n937), .C1(new_n934), .C2(new_n926), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(G72));
  XNOR2_X1  g753(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n680), .B(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n910), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n920), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n459), .B1(new_n482), .B2(new_n500), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n945), .A2(new_n517), .A3(new_n941), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n846), .A2(new_n847), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n884), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n942), .B1(new_n933), .B2(new_n943), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n949), .B1(new_n517), .B2(new_n950), .ZN(G57));
endmodule


