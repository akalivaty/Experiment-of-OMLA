//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214,
    new_n1215;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G137), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT66), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n474), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n473), .B1(G2105), .B2(new_n480), .ZN(G160));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n482), .B1(new_n478), .B2(new_n462), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n461), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n486), .B(new_n488), .C1(new_n489), .C2(new_n463), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND2_X1  g066(.A1(G114), .A2(G2104), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n478), .B2(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n494), .A2(G2105), .B1(G102), .B2(new_n471), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT69), .A2(G138), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n475), .A2(new_n477), .A3(new_n496), .A4(new_n462), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT4), .ZN(new_n499));
  OAI21_X1  g074(.A(G138), .B1(KEYINPUT69), .B2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n461), .A2(new_n462), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n495), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(G543), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n514), .A2(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(G89), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n516), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT71), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n527), .B(new_n523), .C1(new_n516), .C2(new_n524), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n519), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT70), .B(G51), .Z(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n529), .A2(new_n532), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n516), .A2(new_n537), .B1(new_n538), .B2(new_n519), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n511), .A2(G64), .ZN(new_n540));
  INV_X1    g115(.A(G77), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n541), .B2(new_n507), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n539), .B1(G651), .B2(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n513), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n515), .A2(G43), .A3(G543), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n516), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT72), .Z(G188));
  NAND3_X1  g131(.A1(new_n511), .A2(G91), .A3(new_n515), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n515), .A2(G53), .A3(G543), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n508), .A2(new_n510), .A3(G65), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n563), .B1(new_n562), .B2(new_n564), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(KEYINPUT74), .B1(new_n567), .B2(G651), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n562), .A2(new_n564), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT73), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n570), .A2(KEYINPUT74), .A3(G651), .A4(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n557), .B(new_n561), .C1(new_n568), .C2(new_n573), .ZN(G299));
  INV_X1    g149(.A(new_n539), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n542), .A2(G651), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G301));
  INV_X1    g152(.A(G166), .ZN(G303));
  OAI21_X1  g153(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n579));
  INV_X1    g154(.A(G49), .ZN(new_n580));
  INV_X1    g155(.A(G87), .ZN(new_n581));
  OAI221_X1 g156(.A(new_n579), .B1(new_n580), .B2(new_n519), .C1(new_n581), .C2(new_n516), .ZN(G288));
  AOI22_X1  g157(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n513), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  INV_X1    g160(.A(G48), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n516), .A2(new_n585), .B1(new_n586), .B2(new_n519), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n516), .A2(new_n590), .B1(new_n591), .B2(new_n519), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT75), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n513), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n516), .B2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n511), .A2(KEYINPUT10), .A3(G92), .A4(new_n515), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(new_n513), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n530), .A2(G54), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n597), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n597), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(new_n557), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n570), .A2(G651), .A3(new_n571), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT74), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI211_X1 g189(.A(new_n611), .B(new_n560), .C1(new_n614), .C2(new_n572), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n610), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n610), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n607), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n607), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n461), .A2(new_n471), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT13), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2100), .ZN(new_n627));
  INV_X1    g202(.A(G135), .ZN(new_n628));
  NOR2_X1   g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n630));
  OAI22_X1  g205(.A1(new_n463), .A2(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(G123), .B2(new_n485), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n627), .A2(new_n633), .ZN(G156));
  INV_X1    g209(.A(G14), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT15), .B(G2435), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT16), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n642), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n635), .B1(new_n648), .B2(KEYINPUT76), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n645), .A2(new_n647), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n649), .B(new_n650), .C1(KEYINPUT76), .C2(new_n648), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT77), .ZN(G401));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2067), .B(G2678), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT17), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n661), .B(new_n662), .C1(new_n660), .C2(new_n656), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2096), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n669), .A2(KEYINPUT78), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(KEYINPUT78), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT79), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n667), .A2(new_n668), .ZN(new_n679));
  OR3_X1    g254(.A1(new_n673), .A2(new_n669), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n673), .A2(new_n679), .ZN(new_n682));
  NAND4_X1  g257(.A1(new_n678), .A2(new_n680), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1986), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1991), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n685), .B(new_n688), .ZN(G229));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G23), .ZN(new_n691));
  INV_X1    g266(.A(G288), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n690), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT33), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G1976), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n690), .A2(G6), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n588), .B2(new_n690), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT32), .B(G1981), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n690), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n690), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1971), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n697), .B2(new_n698), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n699), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT82), .B(KEYINPUT34), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(G16), .A2(G24), .ZN(new_n712));
  XOR2_X1   g287(.A(G290), .B(KEYINPUT81), .Z(new_n713));
  AOI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(G16), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1986), .ZN(new_n715));
  NOR2_X1   g290(.A1(G25), .A2(G29), .ZN(new_n716));
  INV_X1    g291(.A(G131), .ZN(new_n717));
  NOR2_X1   g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n719));
  OAI22_X1  g294(.A1(new_n463), .A2(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G119), .B2(new_n485), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT80), .Z(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n716), .B1(new_n723), .B2(G29), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  XOR2_X1   g300(.A(new_n724), .B(new_n725), .Z(new_n726));
  NOR2_X1   g301(.A1(new_n715), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n699), .A2(new_n707), .A3(new_n703), .A4(new_n709), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n711), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(KEYINPUT36), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT36), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n711), .A2(new_n727), .A3(new_n731), .A4(new_n728), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(G171), .A2(G16), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G5), .B2(G16), .ZN(new_n735));
  INV_X1    g310(.A(G1961), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n690), .A2(G19), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n549), .B2(new_n690), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n737), .B1(G1341), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n485), .A2(G129), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n464), .A2(G141), .B1(G105), .B2(new_n471), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT26), .Z(new_n744));
  NAND3_X1  g319(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G29), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G29), .B2(G32), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT27), .B(G1996), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n739), .A2(G1341), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n632), .A2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G28), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n753), .B2(KEYINPUT30), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(KEYINPUT30), .B2(new_n753), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n735), .B2(new_n736), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n740), .A2(new_n750), .A3(new_n751), .A4(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G29), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G26), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT85), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT28), .ZN(new_n762));
  INV_X1    g337(.A(G140), .ZN(new_n763));
  NOR2_X1   g338(.A1(G104), .A2(G2105), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n765));
  OAI22_X1  g340(.A1(new_n463), .A2(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G128), .B2(new_n485), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n762), .B1(new_n767), .B2(new_n759), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT86), .B(G2067), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(G16), .A2(G21), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G286), .B2(new_n690), .ZN(new_n772));
  INV_X1    g347(.A(G1966), .ZN(new_n773));
  OR2_X1    g348(.A1(KEYINPUT24), .A2(G34), .ZN(new_n774));
  NAND2_X1  g349(.A1(KEYINPUT24), .A2(G34), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n774), .A2(new_n759), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G160), .B2(new_n759), .ZN(new_n777));
  OAI221_X1 g352(.A(new_n770), .B1(new_n772), .B2(new_n773), .C1(new_n777), .C2(G2084), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n690), .A2(G4), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n607), .B2(new_n690), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1348), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n759), .A2(G27), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G164), .B2(new_n759), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2078), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n758), .A2(new_n778), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n471), .A2(G103), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT25), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n464), .A2(G139), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n787), .B(new_n788), .C1(new_n462), .C2(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G33), .B(new_n790), .S(G29), .Z(new_n791));
  AOI22_X1  g366(.A1(new_n748), .A2(new_n749), .B1(new_n791), .B2(G2072), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n777), .A2(G2084), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n792), .B(new_n793), .C1(G2072), .C2(new_n791), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT87), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(KEYINPUT23), .B1(new_n615), .B2(new_n690), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n690), .A2(G20), .ZN(new_n798));
  MUX2_X1   g373(.A(KEYINPUT23), .B(new_n797), .S(new_n798), .Z(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(G1956), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n759), .A2(G35), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n490), .B2(G29), .ZN(new_n802));
  MUX2_X1   g377(.A(new_n801), .B(new_n802), .S(KEYINPUT89), .Z(new_n803));
  XOR2_X1   g378(.A(KEYINPUT29), .B(G2090), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n772), .A2(new_n773), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT88), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n785), .A2(new_n796), .A3(new_n800), .A4(new_n808), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT31), .B(G11), .Z(new_n810));
  AND2_X1   g385(.A1(new_n799), .A2(G1956), .ZN(new_n811));
  NOR4_X1   g386(.A1(new_n809), .A2(KEYINPUT90), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT90), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n733), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(G311));
  NAND2_X1  g392(.A1(new_n816), .A2(KEYINPUT91), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT91), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n733), .B(new_n819), .C1(new_n812), .C2(new_n815), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(G150));
  AOI22_X1  g396(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n513), .ZN(new_n823));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  INV_X1    g399(.A(G55), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n516), .A2(new_n824), .B1(new_n825), .B2(new_n519), .ZN(new_n826));
  OAI21_X1  g401(.A(G860), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT93), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT92), .B(KEYINPUT37), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n607), .A2(G559), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT38), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n549), .B1(new_n823), .B2(new_n826), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n823), .A2(new_n826), .ZN(new_n834));
  OAI221_X1 g409(.A(new_n546), .B1(new_n516), .B2(new_n547), .C1(new_n544), .C2(new_n513), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT39), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n832), .B(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n830), .B1(new_n839), .B2(G860), .ZN(G145));
  XNOR2_X1  g415(.A(G160), .B(new_n632), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n490), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT95), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(new_n625), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT95), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n842), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n625), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n494), .A2(G2105), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n471), .A2(G102), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n504), .A2(KEYINPUT94), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT94), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n499), .A2(new_n854), .A3(new_n503), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n852), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n767), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n485), .A2(G130), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n464), .A2(G142), .ZN(new_n859));
  NOR2_X1   g434(.A1(G106), .A2(G2105), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n858), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n745), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n857), .B(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n790), .B(new_n721), .Z(new_n865));
  XOR2_X1   g440(.A(new_n864), .B(new_n865), .Z(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n849), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n844), .A2(new_n848), .A3(new_n866), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g447(.A(new_n620), .B(new_n837), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT96), .B1(new_n615), .B2(new_n606), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT96), .ZN(new_n875));
  NAND3_X1  g450(.A1(G299), .A2(new_n875), .A3(new_n607), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(G299), .B2(new_n607), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n611), .B1(new_n614), .B2(new_n572), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n880), .A2(KEYINPUT97), .A3(new_n561), .A4(new_n606), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n873), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT97), .B1(new_n615), .B2(new_n606), .ZN(new_n884));
  INV_X1    g459(.A(new_n881), .ZN(new_n885));
  AOI211_X1 g460(.A(KEYINPUT96), .B(new_n606), .C1(new_n880), .C2(new_n561), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n875), .B1(G299), .B2(new_n607), .ZN(new_n887));
  OAI22_X1  g462(.A1(new_n884), .A2(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n877), .A2(KEYINPUT41), .A3(new_n882), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n883), .B1(new_n892), .B2(new_n873), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n883), .A2(KEYINPUT98), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(G290), .A2(new_n692), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n593), .A2(G288), .A3(new_n595), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(KEYINPUT99), .A3(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(G166), .B(new_n588), .Z(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT99), .B1(new_n899), .B2(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n906));
  INV_X1    g481(.A(new_n900), .ZN(new_n907));
  AOI21_X1  g482(.A(G288), .B1(new_n593), .B2(new_n595), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n901), .A3(new_n902), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n911), .A2(KEYINPUT100), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n898), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n912), .B1(new_n898), .B2(new_n913), .ZN(new_n915));
  OAI21_X1  g490(.A(G868), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(G868), .B2(new_n834), .ZN(G295));
  OAI21_X1  g492(.A(new_n916), .B1(G868), .B2(new_n834), .ZN(G331));
  NAND2_X1  g493(.A1(new_n905), .A2(new_n910), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT102), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n890), .A2(new_n921), .A3(new_n891), .ZN(new_n922));
  NAND2_X1  g497(.A1(G286), .A2(G171), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n529), .A2(G301), .A3(new_n532), .A4(new_n534), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n833), .A2(new_n836), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n926), .B1(new_n833), .B2(new_n836), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n837), .A2(KEYINPUT101), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n931), .A2(new_n923), .A3(new_n927), .A4(new_n924), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT41), .B1(new_n877), .B2(new_n882), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n933), .B1(new_n934), .B2(KEYINPUT103), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n922), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n888), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n936), .B1(new_n922), .B2(new_n935), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n920), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n933), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n877), .A2(KEYINPUT41), .A3(new_n882), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n943), .B2(new_n934), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(new_n911), .A3(new_n938), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n869), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n941), .A2(KEYINPUT43), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n919), .B(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n944), .A2(new_n938), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n949), .B1(new_n953), .B2(new_n946), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n948), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT44), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n943), .A2(new_n934), .A3(KEYINPUT103), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n888), .A2(KEYINPUT103), .A3(new_n889), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n942), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT104), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(new_n938), .A3(new_n937), .ZN(new_n962));
  AOI211_X1 g537(.A(KEYINPUT43), .B(new_n946), .C1(new_n962), .C2(new_n920), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n951), .A2(new_n952), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n949), .B1(new_n964), .B2(new_n947), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n957), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n956), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n957), .B1(new_n948), .B2(new_n954), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n941), .A2(new_n949), .A3(new_n947), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT43), .B1(new_n953), .B2(new_n946), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT44), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT105), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n968), .A2(new_n973), .ZN(G397));
  NAND2_X1  g549(.A1(new_n480), .A2(G2105), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n469), .A2(G40), .A3(new_n975), .A4(new_n472), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n499), .A2(new_n854), .A3(new_n503), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n854), .B1(new_n499), .B2(new_n503), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n495), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n977), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n767), .B(G2067), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n745), .A2(G1996), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n721), .B(new_n725), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(G290), .B(G1986), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n985), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(G303), .A2(G8), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n995), .B(KEYINPUT55), .Z(new_n996));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n856), .B2(G1384), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n980), .A2(KEYINPUT106), .A3(new_n981), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT50), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n505), .A2(new_n981), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR4_X1   g579(.A1(new_n1000), .A2(G2090), .A3(new_n976), .A4(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n980), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1001), .A2(new_n983), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1006), .A2(new_n1007), .A3(new_n977), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(G1971), .ZN(new_n1009));
  OAI211_X1 g584(.A(G8), .B(new_n996), .C1(new_n1005), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n856), .A2(new_n997), .A3(G1384), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT106), .B1(new_n980), .B2(new_n981), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n977), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n584), .ZN(new_n1015));
  INV_X1    g590(.A(new_n587), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT107), .B(G1981), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(G1981), .B1(new_n584), .B2(new_n587), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT49), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT49), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1020), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1014), .A2(new_n1023), .A3(G8), .A4(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G288), .A2(new_n696), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n696), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1014), .A2(G8), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n976), .B1(new_n998), .B2(new_n999), .ZN(new_n1031));
  INV_X1    g606(.A(G8), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1031), .A2(new_n1032), .A3(new_n1027), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1026), .B(new_n1030), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT109), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1014), .A2(G8), .A3(new_n1028), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT52), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT109), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n1026), .A4(new_n1030), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1011), .A2(new_n1036), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1026), .A2(new_n696), .A3(new_n692), .ZN(new_n1042));
  AOI211_X1 g617(.A(new_n1032), .B(new_n1031), .C1(new_n1042), .C2(new_n1018), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n998), .A2(KEYINPUT50), .A3(new_n999), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT110), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n1001), .B2(KEYINPUT50), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n505), .A2(KEYINPUT110), .A3(new_n1003), .A4(new_n981), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1044), .A2(new_n977), .A3(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G2090), .ZN(new_n1050));
  OAI21_X1  g625(.A(G8), .B1(new_n1050), .B2(new_n1009), .ZN(new_n1051));
  INV_X1    g626(.A(new_n996), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1035), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1010), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1002), .A2(KEYINPUT45), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n998), .A2(new_n999), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n977), .B(new_n1057), .C1(new_n1058), .C2(KEYINPUT45), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n773), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1003), .ZN(new_n1061));
  INV_X1    g636(.A(G2084), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1004), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n977), .A4(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1060), .A2(new_n1064), .A3(G168), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1056), .B1(new_n1065), .B2(G8), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(G8), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1000), .A2(new_n976), .A3(new_n1004), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1069), .A2(new_n1062), .B1(new_n1059), .B2(new_n773), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT51), .B1(new_n1070), .B2(G168), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1066), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1055), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OR2_X1    g649(.A1(KEYINPUT121), .A2(KEYINPUT53), .ZN(new_n1075));
  NAND2_X1  g650(.A1(KEYINPUT121), .A2(KEYINPUT53), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1006), .A2(new_n977), .A3(new_n1007), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1075), .B(new_n1076), .C1(new_n1077), .C2(G2078), .ZN(new_n1078));
  INV_X1    g653(.A(G2078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT53), .ZN(new_n1080));
  OAI221_X1 g655(.A(new_n1078), .B1(new_n1059), .B2(new_n1080), .C1(new_n1069), .C2(G1961), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G171), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1067), .A2(KEYINPUT51), .ZN(new_n1083));
  AOI21_X1  g658(.A(G168), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1084));
  OAI211_X1 g659(.A(G8), .B(new_n1065), .C1(new_n1084), .C2(new_n1056), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1082), .B1(new_n1086), .B2(KEYINPUT62), .ZN(new_n1087));
  AOI211_X1 g662(.A(new_n1041), .B(new_n1043), .C1(new_n1074), .C2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G1956), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1049), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT114), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1049), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT56), .B(G2072), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT116), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1006), .A2(new_n977), .A3(new_n1007), .A4(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT117), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(new_n1093), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT119), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n880), .B2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(new_n615), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1091), .A2(new_n1103), .A3(new_n1093), .A4(new_n1097), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1099), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1014), .A2(G2067), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1061), .A2(new_n977), .A3(new_n1063), .ZN(new_n1108));
  INV_X1    g683(.A(G1348), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1106), .B1(new_n1110), .B2(new_n606), .ZN(new_n1111));
  OAI22_X1  g686(.A1(new_n1069), .A2(G1348), .B1(G2067), .B2(new_n1014), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(KEYINPUT118), .A3(new_n607), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1102), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1091), .A2(new_n1114), .A3(new_n1093), .A4(new_n1097), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1105), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1049), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1092), .B1(new_n1049), .B2(new_n1089), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1096), .B(new_n1121), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1118), .B1(new_n1123), .B2(new_n1114), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1115), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n1118), .A3(new_n1114), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n607), .B1(new_n1110), .B2(KEYINPUT60), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT60), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1112), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT120), .B1(new_n1110), .B2(KEYINPUT60), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1128), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT58), .B(G1341), .Z(new_n1134));
  AOI22_X1  g709(.A1(new_n1014), .A2(new_n1134), .B1(new_n1008), .B2(new_n988), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(new_n835), .ZN(new_n1136));
  XOR2_X1   g711(.A(new_n1136), .B(KEYINPUT59), .Z(new_n1137));
  OAI21_X1  g712(.A(new_n1129), .B1(new_n1112), .B2(new_n1130), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n606), .B1(new_n1112), .B2(new_n1130), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1110), .A2(KEYINPUT120), .A3(KEYINPUT60), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1133), .A2(new_n1137), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1117), .B1(new_n1127), .B2(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1053), .A2(new_n1010), .A3(new_n1054), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1086), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1069), .B2(G1961), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1108), .A2(KEYINPUT122), .A3(new_n736), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n982), .A2(new_n983), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n473), .A2(new_n1080), .ZN(new_n1150));
  INV_X1    g725(.A(G40), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n480), .B(KEYINPUT123), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1151), .B1(new_n1152), .B2(G2105), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1149), .A2(new_n1006), .A3(new_n1150), .A4(new_n1153), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1078), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1147), .A2(new_n1148), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT124), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT124), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1147), .A2(new_n1148), .A3(new_n1158), .A4(new_n1155), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1157), .A2(G171), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT54), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n1081), .B2(G301), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1082), .B(new_n1161), .C1(G171), .C2(new_n1156), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1145), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1143), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1088), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT63), .ZN(new_n1168));
  OR3_X1    g743(.A1(new_n1070), .A2(new_n1032), .A3(G286), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1168), .B1(new_n1055), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT111), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g747(.A(KEYINPUT111), .B(new_n1168), .C1(new_n1055), .C2(new_n1169), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(G8), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1052), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1176), .A2(new_n1036), .A3(new_n1040), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(KEYINPUT112), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT112), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1176), .A2(new_n1036), .A3(new_n1179), .A4(new_n1040), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1169), .A2(new_n1168), .A3(new_n1011), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(KEYINPUT113), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT113), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1181), .A2(new_n1185), .A3(new_n1182), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1174), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n994), .B1(new_n1167), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(KEYINPUT46), .B1(new_n985), .B2(new_n988), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n984), .B1(new_n746), .B2(new_n986), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT46), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n984), .A2(new_n1191), .A3(G1996), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n1193), .B(KEYINPUT125), .Z(new_n1194));
  INV_X1    g769(.A(KEYINPUT47), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n984), .A2(G1986), .A3(G290), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT126), .ZN(new_n1198));
  XOR2_X1   g773(.A(new_n1198), .B(KEYINPUT48), .Z(new_n1199));
  NAND2_X1  g774(.A1(new_n992), .A2(new_n985), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1202));
  INV_X1    g777(.A(G2067), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n767), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n723), .A2(new_n725), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1204), .B1(new_n1205), .B2(new_n990), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(new_n985), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n1196), .A2(new_n1201), .A3(new_n1202), .A4(new_n1207), .ZN(new_n1208));
  XOR2_X1   g783(.A(new_n1208), .B(KEYINPUT127), .Z(new_n1209));
  NAND2_X1  g784(.A1(new_n1188), .A2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g785(.A(G227), .ZN(new_n1212));
  NAND3_X1  g786(.A1(new_n871), .A2(new_n651), .A3(new_n1212), .ZN(new_n1213));
  NOR2_X1   g787(.A1(new_n963), .A2(new_n965), .ZN(new_n1214));
  OR2_X1    g788(.A1(G229), .A2(new_n459), .ZN(new_n1215));
  NOR3_X1   g789(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(G308));
  INV_X1    g790(.A(G308), .ZN(G225));
endmodule


