

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XOR2_X1 U321 ( .A(G15GAT), .B(G127GAT), .Z(n442) );
  XNOR2_X1 U322 ( .A(n343), .B(n325), .ZN(n326) );
  XNOR2_X1 U323 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U324 ( .A(n463), .B(n471), .Z(n537) );
  AND2_X1 U325 ( .A1(G231GAT), .A2(G233GAT), .ZN(n289) );
  XOR2_X1 U326 ( .A(KEYINPUT97), .B(n466), .Z(n290) );
  NOR2_X1 U327 ( .A1(n532), .A2(n534), .ZN(n465) );
  INV_X1 U328 ( .A(KEYINPUT95), .ZN(n323) );
  XNOR2_X1 U329 ( .A(n386), .B(n289), .ZN(n387) );
  INV_X1 U330 ( .A(KEYINPUT7), .ZN(n335) );
  XNOR2_X1 U331 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U332 ( .A(n336), .B(n335), .ZN(n338) );
  XNOR2_X1 U333 ( .A(n426), .B(n340), .ZN(n341) );
  XNOR2_X1 U334 ( .A(n338), .B(n337), .ZN(n360) );
  XNOR2_X1 U335 ( .A(n342), .B(n341), .ZN(n345) );
  NOR2_X1 U336 ( .A1(n496), .A2(n581), .ZN(n497) );
  XOR2_X1 U337 ( .A(n400), .B(n399), .Z(n558) );
  XOR2_X1 U338 ( .A(n347), .B(n346), .Z(n479) );
  XOR2_X1 U339 ( .A(n447), .B(n446), .Z(n534) );
  XOR2_X1 U340 ( .A(n378), .B(n331), .Z(n524) );
  XNOR2_X1 U341 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U342 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT93), .B(KEYINPUT4), .Z(n292) );
  XNOR2_X1 U344 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n291) );
  XNOR2_X1 U345 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U346 ( .A(KEYINPUT90), .B(KEYINPUT1), .Z(n294) );
  XNOR2_X1 U347 ( .A(KEYINPUT5), .B(KEYINPUT6), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U349 ( .A(n296), .B(n295), .Z(n306) );
  XOR2_X1 U350 ( .A(KEYINPUT88), .B(G155GAT), .Z(n298) );
  XNOR2_X1 U351 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U353 ( .A(KEYINPUT87), .B(n299), .Z(n431) );
  XOR2_X1 U354 ( .A(G134GAT), .B(KEYINPUT75), .Z(n339) );
  XOR2_X1 U355 ( .A(KEYINPUT0), .B(KEYINPUT83), .Z(n301) );
  XNOR2_X1 U356 ( .A(G113GAT), .B(G120GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n438) );
  XOR2_X1 U358 ( .A(n339), .B(n438), .Z(n303) );
  NAND2_X1 U359 ( .A1(G225GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U361 ( .A(n431), .B(n304), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n314) );
  XOR2_X1 U363 ( .A(G148GAT), .B(G57GAT), .Z(n308) );
  XNOR2_X1 U364 ( .A(G141GAT), .B(G127GAT), .ZN(n307) );
  XNOR2_X1 U365 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U366 ( .A(G162GAT), .B(G85GAT), .Z(n310) );
  XNOR2_X1 U367 ( .A(G29GAT), .B(G1GAT), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U369 ( .A(n312), .B(n311), .Z(n313) );
  XOR2_X1 U370 ( .A(n314), .B(n313), .Z(n476) );
  XOR2_X1 U371 ( .A(G92GAT), .B(G64GAT), .Z(n316) );
  XNOR2_X1 U372 ( .A(G176GAT), .B(G204GAT), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U374 ( .A(KEYINPUT73), .B(n317), .Z(n378) );
  XOR2_X1 U375 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n319) );
  XNOR2_X1 U376 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n439) );
  XOR2_X1 U378 ( .A(KEYINPUT86), .B(KEYINPUT21), .Z(n321) );
  XNOR2_X1 U379 ( .A(G197GAT), .B(G211GAT), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n321), .B(n320), .ZN(n418) );
  XNOR2_X1 U381 ( .A(n439), .B(n418), .ZN(n327) );
  XNOR2_X1 U382 ( .A(G36GAT), .B(G190GAT), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n322), .B(G218GAT), .ZN(n343) );
  NAND2_X1 U384 ( .A1(G226GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U386 ( .A(n328), .B(KEYINPUT94), .Z(n330) );
  XOR2_X1 U387 ( .A(G169GAT), .B(G8GAT), .Z(n355) );
  XNOR2_X1 U388 ( .A(n355), .B(KEYINPUT76), .ZN(n329) );
  XNOR2_X1 U389 ( .A(n330), .B(n329), .ZN(n331) );
  INV_X1 U390 ( .A(n524), .ZN(n412) );
  XOR2_X1 U391 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n333) );
  NAND2_X1 U392 ( .A1(G232GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U394 ( .A(G92GAT), .B(n334), .ZN(n347) );
  XNOR2_X1 U395 ( .A(G43GAT), .B(G29GAT), .ZN(n336) );
  XOR2_X1 U396 ( .A(KEYINPUT69), .B(KEYINPUT8), .Z(n337) );
  XNOR2_X1 U397 ( .A(n360), .B(n339), .ZN(n342) );
  XOR2_X1 U398 ( .A(G50GAT), .B(G162GAT), .Z(n426) );
  XNOR2_X1 U399 ( .A(KEYINPUT11), .B(G106GAT), .ZN(n340) );
  XOR2_X1 U400 ( .A(G99GAT), .B(G85GAT), .Z(n372) );
  XNOR2_X1 U401 ( .A(n372), .B(n343), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n346) );
  INV_X1 U403 ( .A(n479), .ZN(n404) );
  XOR2_X1 U404 ( .A(KEYINPUT65), .B(G197GAT), .Z(n349) );
  XNOR2_X1 U405 ( .A(KEYINPUT67), .B(KEYINPUT66), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n364) );
  XOR2_X1 U407 ( .A(KEYINPUT68), .B(G15GAT), .Z(n351) );
  XNOR2_X1 U408 ( .A(G113GAT), .B(KEYINPUT29), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U410 ( .A(n352), .B(G50GAT), .Z(n354) );
  XOR2_X1 U411 ( .A(G141GAT), .B(G22GAT), .Z(n427) );
  XNOR2_X1 U412 ( .A(n427), .B(G36GAT), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n359) );
  XOR2_X1 U414 ( .A(n355), .B(KEYINPUT30), .Z(n357) );
  NAND2_X1 U415 ( .A1(G229GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U417 ( .A(n359), .B(n358), .Z(n362) );
  XOR2_X1 U418 ( .A(KEYINPUT70), .B(G1GAT), .Z(n381) );
  XNOR2_X1 U419 ( .A(n360), .B(n381), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n551) );
  INV_X1 U422 ( .A(n551), .ZN(n569) );
  XOR2_X1 U423 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n366) );
  XNOR2_X1 U424 ( .A(G71GAT), .B(G57GAT), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n390) );
  XOR2_X1 U426 ( .A(G78GAT), .B(KEYINPUT72), .Z(n368) );
  XNOR2_X1 U427 ( .A(G148GAT), .B(G106GAT), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n419) );
  XNOR2_X1 U429 ( .A(n390), .B(n419), .ZN(n376) );
  XOR2_X1 U430 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n370) );
  XNOR2_X1 U431 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U433 ( .A(n372), .B(n371), .Z(n374) );
  NAND2_X1 U434 ( .A1(G230GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n378), .B(n377), .ZN(n573) );
  XOR2_X1 U438 ( .A(n573), .B(KEYINPUT41), .Z(n554) );
  NOR2_X1 U439 ( .A1(n569), .A2(n554), .ZN(n380) );
  XNOR2_X1 U440 ( .A(KEYINPUT113), .B(KEYINPUT46), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n401) );
  XOR2_X1 U442 ( .A(n442), .B(G22GAT), .Z(n383) );
  XNOR2_X1 U443 ( .A(n381), .B(G8GAT), .ZN(n382) );
  XNOR2_X1 U444 ( .A(n383), .B(n382), .ZN(n388) );
  XOR2_X1 U445 ( .A(KEYINPUT80), .B(KEYINPUT14), .Z(n385) );
  XNOR2_X1 U446 ( .A(G183GAT), .B(KEYINPUT76), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U448 ( .A(n389), .B(KEYINPUT79), .Z(n392) );
  XNOR2_X1 U449 ( .A(n390), .B(KEYINPUT78), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n400) );
  XOR2_X1 U451 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n394) );
  XNOR2_X1 U452 ( .A(G155GAT), .B(G211GAT), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U454 ( .A(KEYINPUT77), .B(KEYINPUT81), .Z(n396) );
  XNOR2_X1 U455 ( .A(G64GAT), .B(G78GAT), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U457 ( .A(n398), .B(n397), .Z(n399) );
  INV_X1 U458 ( .A(n558), .ZN(n576) );
  NAND2_X1 U459 ( .A1(n401), .A2(n576), .ZN(n402) );
  NOR2_X1 U460 ( .A1(n404), .A2(n402), .ZN(n403) );
  XNOR2_X1 U461 ( .A(KEYINPUT47), .B(n403), .ZN(n409) );
  XOR2_X1 U462 ( .A(n404), .B(KEYINPUT36), .Z(n581) );
  NOR2_X1 U463 ( .A1(n581), .A2(n576), .ZN(n405) );
  XOR2_X1 U464 ( .A(KEYINPUT45), .B(n405), .Z(n406) );
  NOR2_X1 U465 ( .A1(n551), .A2(n406), .ZN(n407) );
  NAND2_X1 U466 ( .A1(n407), .A2(n573), .ZN(n408) );
  NAND2_X1 U467 ( .A1(n409), .A2(n408), .ZN(n411) );
  INV_X1 U468 ( .A(KEYINPUT48), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n533) );
  NOR2_X1 U470 ( .A1(n412), .A2(n533), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n413), .B(KEYINPUT54), .ZN(n414) );
  AND2_X1 U472 ( .A1(n476), .A2(n414), .ZN(n568) );
  XOR2_X1 U473 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n416) );
  NAND2_X1 U474 ( .A1(G228GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U476 ( .A(n417), .B(KEYINPUT23), .Z(n421) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U479 ( .A(KEYINPUT89), .B(KEYINPUT85), .Z(n423) );
  XNOR2_X1 U480 ( .A(G204GAT), .B(G218GAT), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U482 ( .A(n425), .B(n424), .Z(n429) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n471) );
  NAND2_X1 U486 ( .A1(n568), .A2(n471), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n432), .B(KEYINPUT55), .ZN(n448) );
  XOR2_X1 U488 ( .A(G71GAT), .B(G134GAT), .Z(n434) );
  XNOR2_X1 U489 ( .A(G169GAT), .B(G99GAT), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n447) );
  XOR2_X1 U491 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n436) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U494 ( .A(n437), .B(G176GAT), .Z(n441) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U497 ( .A(n443), .B(n442), .Z(n445) );
  XNOR2_X1 U498 ( .A(G43GAT), .B(G190GAT), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U500 ( .A1(n448), .A2(n534), .ZN(n449) );
  XNOR2_X1 U501 ( .A(KEYINPUT120), .B(n449), .ZN(n564) );
  NOR2_X1 U502 ( .A1(n564), .A2(n479), .ZN(n453) );
  XNOR2_X1 U503 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n451) );
  INV_X1 U504 ( .A(G190GAT), .ZN(n450) );
  XNOR2_X1 U505 ( .A(KEYINPUT107), .B(n554), .ZN(n540) );
  INV_X1 U506 ( .A(n540), .ZN(n454) );
  NOR2_X1 U507 ( .A1(n564), .A2(n454), .ZN(n458) );
  XNOR2_X1 U508 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n456) );
  XNOR2_X1 U509 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n455) );
  XNOR2_X1 U510 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  NOR2_X1 U512 ( .A1(n569), .A2(n564), .ZN(n460) );
  XNOR2_X1 U513 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n459) );
  XNOR2_X1 U514 ( .A(n460), .B(n459), .ZN(G1348GAT) );
  XOR2_X1 U515 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n485) );
  NAND2_X1 U516 ( .A1(n573), .A2(n551), .ZN(n461) );
  XNOR2_X1 U517 ( .A(n461), .B(KEYINPUT74), .ZN(n498) );
  XOR2_X1 U518 ( .A(KEYINPUT27), .B(KEYINPUT96), .Z(n462) );
  XOR2_X1 U519 ( .A(n524), .B(n462), .Z(n469) );
  INV_X1 U520 ( .A(n476), .ZN(n521) );
  NAND2_X1 U521 ( .A1(n469), .A2(n521), .ZN(n532) );
  XNOR2_X1 U522 ( .A(KEYINPUT64), .B(KEYINPUT28), .ZN(n463) );
  INV_X1 U523 ( .A(n537), .ZN(n464) );
  NAND2_X1 U524 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n534), .A2(n471), .ZN(n468) );
  XNOR2_X1 U526 ( .A(KEYINPUT98), .B(KEYINPUT26), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n468), .B(n467), .ZN(n567) );
  NAND2_X1 U528 ( .A1(n469), .A2(n567), .ZN(n475) );
  AND2_X1 U529 ( .A1(n534), .A2(n524), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n470), .B(KEYINPUT99), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n472), .A2(n471), .ZN(n473) );
  XOR2_X1 U532 ( .A(KEYINPUT25), .B(n473), .Z(n474) );
  NAND2_X1 U533 ( .A1(n475), .A2(n474), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U535 ( .A1(n290), .A2(n478), .ZN(n494) );
  XOR2_X1 U536 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n481) );
  NAND2_X1 U537 ( .A1(n558), .A2(n479), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n481), .B(n480), .ZN(n482) );
  NAND2_X1 U539 ( .A1(n494), .A2(n482), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n483), .B(KEYINPUT100), .ZN(n509) );
  NOR2_X1 U541 ( .A1(n498), .A2(n509), .ZN(n492) );
  NAND2_X1 U542 ( .A1(n492), .A2(n521), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U545 ( .A1(n492), .A2(n524), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n487), .B(KEYINPUT102), .ZN(n488) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(n488), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U549 ( .A1(n492), .A2(n534), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U551 ( .A(G15GAT), .B(n491), .Z(G1326GAT) );
  NAND2_X1 U552 ( .A1(n492), .A2(n537), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT39), .Z(n501) );
  NAND2_X1 U555 ( .A1(n576), .A2(n494), .ZN(n495) );
  XNOR2_X1 U556 ( .A(KEYINPUT104), .B(n495), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(KEYINPUT37), .ZN(n520) );
  NOR2_X1 U558 ( .A1(n498), .A2(n520), .ZN(n499) );
  XNOR2_X1 U559 ( .A(KEYINPUT38), .B(n499), .ZN(n506) );
  NAND2_X1 U560 ( .A1(n506), .A2(n521), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U562 ( .A1(n524), .A2(n506), .ZN(n502) );
  XNOR2_X1 U563 ( .A(G36GAT), .B(n502), .ZN(G1329GAT) );
  NAND2_X1 U564 ( .A1(n506), .A2(n534), .ZN(n504) );
  XOR2_X1 U565 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G43GAT), .B(n505), .ZN(G1330GAT) );
  XNOR2_X1 U568 ( .A(G50GAT), .B(KEYINPUT106), .ZN(n508) );
  NAND2_X1 U569 ( .A1(n537), .A2(n506), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n508), .B(n507), .ZN(G1331GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n511) );
  NAND2_X1 U572 ( .A1(n569), .A2(n540), .ZN(n519) );
  NOR2_X1 U573 ( .A1(n509), .A2(n519), .ZN(n516) );
  NAND2_X1 U574 ( .A1(n516), .A2(n521), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U576 ( .A(G57GAT), .B(n512), .Z(G1332GAT) );
  XOR2_X1 U577 ( .A(G64GAT), .B(KEYINPUT109), .Z(n514) );
  NAND2_X1 U578 ( .A1(n516), .A2(n524), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n516), .A2(n534), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n515), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U583 ( .A1(n516), .A2(n537), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NOR2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n527) );
  NAND2_X1 U586 ( .A1(n521), .A2(n527), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(KEYINPUT110), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U589 ( .A1(n527), .A2(n524), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n527), .A2(n534), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n526), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(KEYINPUT111), .ZN(n531) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n529) );
  NAND2_X1 U595 ( .A1(n527), .A2(n537), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1339GAT) );
  XOR2_X1 U598 ( .A(G113GAT), .B(KEYINPUT115), .Z(n539) );
  NOR2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n549) );
  NAND2_X1 U600 ( .A1(n534), .A2(n549), .ZN(n535) );
  XNOR2_X1 U601 ( .A(KEYINPUT114), .B(n535), .ZN(n536) );
  NOR2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n546), .A2(n551), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n542) );
  NAND2_X1 U606 ( .A1(n546), .A2(n540), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(n543), .ZN(G1341GAT) );
  NAND2_X1 U609 ( .A1(n546), .A2(n558), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n544), .B(KEYINPUT50), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U613 ( .A1(n546), .A2(n404), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n549), .A2(n567), .ZN(n550) );
  XOR2_X1 U616 ( .A(n550), .B(KEYINPUT117), .Z(n553) );
  INV_X1 U617 ( .A(n553), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n561), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n556) );
  XNOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n561), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT118), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(n560), .ZN(G1346GAT) );
  XOR2_X1 U627 ( .A(G162GAT), .B(KEYINPUT119), .Z(n563) );
  NAND2_X1 U628 ( .A1(n561), .A2(n404), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1347GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n576), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n580) );
  NOR2_X1 U634 ( .A1(n569), .A2(n580), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n580), .ZN(n575) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n580), .ZN(n577) );
  XOR2_X1 U642 ( .A(G211GAT), .B(n577), .Z(G1354GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT62), .Z(n579) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n583) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(n583), .B(n582), .Z(G1355GAT) );
endmodule

