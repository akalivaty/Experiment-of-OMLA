//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT3), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G107), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n187), .A2(KEYINPUT3), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n188), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(G107), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT76), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n193), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(G101), .B1(new_n192), .B2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n196), .A2(G104), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(new_n188), .B2(new_n190), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n194), .A2(KEYINPUT76), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n195), .B1(new_n203), .B2(new_n197), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n199), .A2(KEYINPUT4), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G116), .ZN(new_n208));
  INV_X1    g022(.A(G116), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G119), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT2), .ZN(new_n214));
  INV_X1    g028(.A(G113), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT66), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(KEYINPUT2), .B2(G113), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n212), .A2(new_n218), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n211), .A2(KEYINPUT68), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n208), .A2(new_n210), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n216), .A2(new_n217), .B1(new_n219), .B2(new_n221), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n223), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n202), .B1(new_n201), .B2(new_n204), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n206), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n208), .A2(new_n210), .A3(new_n225), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n225), .B1(new_n208), .B2(new_n210), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n208), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n215), .B1(new_n234), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(G101), .B1(new_n190), .B2(new_n200), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n241), .A2(new_n205), .A3(new_n223), .A4(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n233), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(G110), .B(G122), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n233), .A2(new_n243), .A3(new_n245), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(KEYINPUT6), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT6), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n244), .A2(new_n250), .A3(new_n246), .ZN(new_n251));
  INV_X1    g065(.A(G128), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  INV_X1    g068(.A(G146), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G143), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n252), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G125), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n252), .A2(KEYINPUT1), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n253), .A2(G146), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n256), .A2(KEYINPUT1), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n258), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT80), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n261), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n267), .A2(new_n252), .B1(KEYINPUT1), .B2(new_n256), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n268), .A2(KEYINPUT80), .A3(new_n258), .A4(new_n262), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT0), .A4(G128), .ZN(new_n271));
  XNOR2_X1  g085(.A(G143), .B(G146), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT0), .B(G128), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G125), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G224), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(G953), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n276), .B(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n249), .A2(new_n251), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(G210), .B1(G237), .B2(G902), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT82), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT81), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n266), .A2(new_n285), .A3(new_n269), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(new_n266), .B2(new_n269), .ZN(new_n287));
  INV_X1    g101(.A(new_n275), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT7), .B1(new_n277), .B2(G953), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n284), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n270), .A2(KEYINPUT81), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n275), .ZN(new_n294));
  OAI211_X1 g108(.A(KEYINPUT82), .B(new_n290), .C1(new_n294), .C2(new_n286), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT5), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n240), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n223), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(new_n205), .A3(new_n242), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n205), .A2(new_n242), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n241), .A2(new_n300), .A3(new_n223), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n245), .B(KEYINPUT8), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n270), .A2(new_n291), .A3(new_n275), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n248), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n292), .A2(new_n295), .A3(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n282), .A2(KEYINPUT83), .A3(new_n283), .A4(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n280), .A3(new_n281), .ZN(new_n308));
  INV_X1    g122(.A(new_n283), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n306), .A2(new_n280), .A3(new_n281), .A4(new_n283), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT83), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n307), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT9), .B(G234), .ZN(new_n315));
  OAI21_X1  g129(.A(G221), .B1(new_n315), .B2(G902), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT11), .ZN(new_n318));
  INV_X1    g132(.A(G134), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(G137), .ZN(new_n320));
  INV_X1    g134(.A(G137), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT11), .A3(G134), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(G137), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G131), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT64), .ZN(new_n326));
  INV_X1    g140(.A(G131), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n320), .A2(new_n322), .A3(new_n327), .A4(new_n323), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n324), .A2(KEYINPUT64), .A3(G131), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n257), .A2(new_n262), .A3(new_n263), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n205), .A2(new_n332), .A3(new_n242), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT10), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT10), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n205), .A2(new_n332), .A3(new_n335), .A4(new_n242), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n274), .B1(new_n230), .B2(new_n231), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n338), .A2(KEYINPUT77), .A3(new_n206), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT77), .B1(new_n338), .B2(new_n206), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n331), .B(new_n337), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(G110), .B(G140), .ZN(new_n342));
  INV_X1    g156(.A(G953), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n343), .A2(G227), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n342), .B(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n348));
  INV_X1    g162(.A(new_n331), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n333), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n332), .B1(new_n205), .B2(new_n242), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n329), .A2(KEYINPUT78), .A3(new_n330), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT12), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n300), .A2(new_n262), .A3(new_n268), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n333), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT12), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n357), .A2(KEYINPUT78), .A3(new_n358), .A4(new_n349), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n341), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n347), .A2(new_n350), .B1(new_n360), .B2(new_n345), .ZN(new_n361));
  OAI21_X1  g175(.A(G469), .B1(new_n361), .B2(G902), .ZN(new_n362));
  INV_X1    g176(.A(G469), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n346), .B1(new_n350), .B2(new_n341), .ZN(new_n364));
  AND4_X1   g178(.A1(new_n341), .A2(new_n346), .A3(new_n355), .A4(new_n359), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n363), .B(new_n281), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n317), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(G214), .B1(G237), .B2(G902), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n314), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G217), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n315), .A2(new_n370), .A3(G953), .ZN(new_n371));
  XNOR2_X1  g185(.A(G128), .B(G143), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(KEYINPUT89), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(G134), .ZN(new_n374));
  INV_X1    g188(.A(G122), .ZN(new_n375));
  OR3_X1    g189(.A1(new_n375), .A2(KEYINPUT14), .A3(G116), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT91), .B1(new_n209), .B2(G122), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT91), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n378), .B1(new_n379), .B2(new_n376), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT14), .B1(new_n375), .B2(G116), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT90), .ZN(new_n382));
  OAI21_X1  g196(.A(G107), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G116), .B(G122), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n196), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n374), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n372), .A2(KEYINPUT13), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n253), .A2(G128), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n387), .B(G134), .C1(KEYINPUT13), .C2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n384), .B(new_n196), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n389), .B(new_n390), .C1(new_n373), .C2(G134), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n371), .B1(new_n386), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n386), .A2(new_n391), .A3(new_n371), .ZN(new_n394));
  AOI21_X1  g208(.A(G902), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G478), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n395), .B1(KEYINPUT15), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n394), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n281), .B1(new_n398), .B2(new_n392), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT15), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(G478), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G952), .ZN(new_n403));
  AOI211_X1 g217(.A(G953), .B(new_n403), .C1(G234), .C2(G237), .ZN(new_n404));
  AOI211_X1 g218(.A(new_n281), .B(new_n343), .C1(G234), .C2(G237), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT21), .B(G898), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT85), .ZN(new_n410));
  INV_X1    g224(.A(G237), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n343), .A3(G214), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n253), .ZN(new_n413));
  NOR2_X1   g227(.A1(G237), .A2(G953), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(G143), .A3(G214), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n410), .B1(new_n416), .B2(G131), .ZN(new_n417));
  AOI211_X1 g231(.A(KEYINPUT85), .B(new_n327), .C1(new_n413), .C2(new_n415), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT17), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AND4_X1   g233(.A1(G143), .A2(new_n411), .A3(new_n343), .A4(G214), .ZN(new_n420));
  AOI21_X1  g234(.A(G143), .B1(new_n414), .B2(G214), .ZN(new_n421));
  OAI21_X1  g235(.A(G131), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT85), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n416), .A2(new_n410), .A3(G131), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT17), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n413), .A2(new_n327), .A3(new_n415), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n423), .A2(new_n424), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G140), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G125), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n258), .A2(G140), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT16), .ZN(new_n431));
  OR3_X1    g245(.A1(new_n258), .A2(KEYINPUT16), .A3(G140), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n255), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n432), .A3(G146), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n419), .A2(new_n427), .A3(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G113), .B(G122), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(new_n189), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n416), .A2(KEYINPUT18), .A3(G131), .ZN(new_n441));
  XNOR2_X1  g255(.A(G125), .B(G140), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(new_n255), .ZN(new_n443));
  NAND2_X1  g257(.A1(KEYINPUT18), .A2(G131), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n413), .A2(new_n415), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n441), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n438), .A2(new_n440), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n435), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n442), .B(KEYINPUT19), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(new_n255), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n440), .B1(new_n452), .B2(new_n446), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n409), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(G475), .A2(G902), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n446), .ZN(new_n456));
  INV_X1    g270(.A(new_n440), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n438), .A2(new_n440), .A3(new_n446), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT86), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n454), .A2(new_n455), .A3(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT87), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n461), .A2(new_n466), .A3(new_n463), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT20), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n455), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n458), .B2(new_n459), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT88), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n465), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n440), .B1(new_n438), .B2(new_n446), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n447), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n281), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n408), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT28), .ZN(new_n478));
  INV_X1    g292(.A(new_n274), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n329), .A2(new_n479), .A3(new_n330), .ZN(new_n480));
  INV_X1    g294(.A(new_n323), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n319), .A2(G137), .ZN(new_n482));
  OAI21_X1  g296(.A(G131), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n332), .A2(new_n328), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n229), .ZN(new_n486));
  INV_X1    g300(.A(new_n229), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n480), .A3(new_n484), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n478), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n478), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT71), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n488), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n487), .B1(new_n480), .B2(new_n484), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT28), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT71), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n414), .A2(G210), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(KEYINPUT27), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT26), .B(G101), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n499), .B(new_n500), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n501), .A2(KEYINPUT29), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n492), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT72), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n489), .A2(new_n491), .ZN(new_n505));
  XOR2_X1   g319(.A(new_n501), .B(KEYINPUT69), .Z(new_n506));
  AOI21_X1  g320(.A(KEYINPUT29), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n501), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n480), .A2(KEYINPUT30), .A3(new_n484), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n229), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT30), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n485), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT65), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n485), .A2(KEYINPUT65), .A3(new_n511), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n510), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n508), .B1(new_n516), .B2(new_n493), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n507), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT72), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n492), .A2(new_n497), .A3(new_n519), .A4(new_n502), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n504), .A2(new_n518), .A3(new_n281), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G472), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n506), .B1(new_n495), .B2(new_n490), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT65), .B1(new_n485), .B2(new_n511), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n513), .B(KEYINPUT30), .C1(new_n480), .C2(new_n484), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n229), .B(new_n509), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n493), .A2(new_n508), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n527), .A2(KEYINPUT31), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT31), .B1(new_n527), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n524), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(G472), .A2(G902), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(KEYINPUT32), .A3(new_n532), .ZN(new_n533));
  XOR2_X1   g347(.A(KEYINPUT70), .B(KEYINPUT32), .Z(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT31), .ZN(new_n536));
  INV_X1    g350(.A(new_n528), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n536), .B1(new_n516), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n527), .A2(KEYINPUT31), .A3(new_n528), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n523), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n532), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n535), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n522), .A2(new_n533), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n370), .B1(G234), .B2(new_n281), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(G902), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT75), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT22), .B(G137), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n343), .A2(G221), .A3(G234), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n207), .A2(G128), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n252), .A2(G119), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT24), .B(G110), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(G146), .B1(new_n431), .B2(new_n432), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n556), .B1(new_n448), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G110), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT23), .B1(new_n252), .B2(G119), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT74), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n552), .A2(KEYINPUT74), .A3(KEYINPUT23), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n553), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT73), .ZN(new_n565));
  NAND2_X1  g379(.A1(KEYINPUT23), .A2(G119), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n565), .B1(new_n566), .B2(G128), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n252), .A2(KEYINPUT73), .A3(KEYINPUT23), .A4(G119), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n559), .B1(new_n564), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n558), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n442), .A2(new_n255), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n435), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n564), .A2(new_n559), .A3(new_n569), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n554), .A2(new_n555), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n551), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n564), .A2(new_n569), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n436), .B(new_n556), .C1(new_n579), .C2(new_n559), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n574), .A2(new_n575), .ZN(new_n581));
  INV_X1    g395(.A(new_n573), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n583), .A3(new_n550), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n547), .B1(new_n578), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n577), .A2(new_n584), .A3(KEYINPUT75), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n546), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n544), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n577), .A2(new_n584), .A3(new_n281), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT25), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n577), .A2(new_n584), .A3(KEYINPUT25), .A4(new_n281), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n369), .A2(new_n477), .A3(new_n543), .A4(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT92), .B(G101), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G3));
  OAI211_X1 g412(.A(KEYINPUT93), .B(G472), .C1(new_n540), .C2(G902), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n531), .A2(new_n532), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n531), .A2(new_n281), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT93), .B1(new_n602), .B2(G472), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n367), .A2(new_n595), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n407), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n310), .A2(new_n311), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT94), .B1(new_n608), .B2(new_n368), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT94), .ZN(new_n610));
  INV_X1    g424(.A(new_n368), .ZN(new_n611));
  AOI211_X1 g425(.A(new_n610), .B(new_n611), .C1(new_n310), .C2(new_n311), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT95), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n614), .B1(new_n394), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(new_n398), .B2(new_n392), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n393), .B(new_n394), .C1(new_n615), .C2(new_n614), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n618), .A3(G478), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n396), .A2(new_n281), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n395), .B2(new_n396), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n472), .B2(new_n476), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n606), .A2(new_n607), .A3(new_n613), .A4(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT34), .B(G104), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  AND2_X1   g440(.A1(new_n454), .A2(new_n460), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n455), .A3(new_n462), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n465), .A2(new_n628), .A3(new_n467), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n397), .A2(new_n401), .B1(G475), .B2(new_n475), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n608), .A2(new_n368), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n610), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n608), .A2(KEYINPUT94), .A3(new_n368), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n631), .A2(new_n633), .A3(new_n607), .A4(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n635), .A2(KEYINPUT96), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n613), .A2(new_n637), .A3(new_n607), .A4(new_n631), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n606), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT97), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NAND2_X1  g457(.A1(new_n580), .A2(new_n583), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n551), .A2(KEYINPUT36), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n646), .A2(new_n545), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n594), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n604), .A2(new_n369), .A3(new_n477), .A4(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  INV_X1    g466(.A(new_n366), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n360), .A2(new_n345), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n350), .A2(new_n341), .A3(new_n346), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(G469), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(G469), .A2(G902), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n316), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n648), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n543), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT98), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n633), .A2(new_n634), .ZN(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n405), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n404), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n629), .A2(new_n630), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n662), .B1(new_n663), .B2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n668), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n613), .A2(new_n670), .A3(KEYINPUT98), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n661), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n252), .ZN(G30));
  XNOR2_X1  g487(.A(new_n667), .B(KEYINPUT39), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n367), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT99), .B(KEYINPUT40), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n402), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n472), .B2(new_n476), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n679), .A2(new_n368), .A3(new_n648), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n314), .B(KEYINPUT38), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n516), .A2(new_n537), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n506), .B1(new_n488), .B2(new_n486), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n281), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G472), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n542), .A2(new_n533), .A3(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n677), .A2(new_n680), .A3(new_n681), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  INV_X1    g502(.A(new_n667), .ZN(new_n689));
  AOI211_X1 g503(.A(new_n622), .B(new_n689), .C1(new_n472), .C2(new_n476), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n690), .A2(new_n613), .A3(new_n543), .A4(new_n660), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  NOR2_X1   g506(.A1(new_n364), .A2(new_n365), .ZN(new_n693));
  OAI21_X1  g507(.A(G469), .B1(new_n693), .B2(G902), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n694), .A2(new_n316), .A3(new_n366), .A4(new_n595), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n542), .A2(new_n533), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n695), .B1(new_n696), .B2(new_n522), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n697), .A2(new_n607), .A3(new_n613), .A4(new_n623), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT41), .B(G113), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT100), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n698), .B(new_n700), .ZN(G15));
  INV_X1    g515(.A(new_n697), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n635), .A2(KEYINPUT96), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n702), .B1(new_n703), .B2(new_n638), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n209), .ZN(G18));
  AND4_X1   g519(.A1(new_n476), .A2(new_n408), .A3(new_n472), .A4(new_n649), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n694), .A2(new_n366), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n317), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n706), .A2(new_n613), .A3(new_n543), .A4(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT101), .B(G119), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G21));
  XNOR2_X1  g525(.A(new_n595), .B(KEYINPUT104), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n496), .B1(new_n495), .B2(new_n490), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n489), .A2(KEYINPUT71), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n506), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n492), .A2(KEYINPUT102), .A3(new_n497), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n538), .A2(new_n539), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n541), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT103), .B(G472), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n531), .B2(new_n281), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n712), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n707), .A2(new_n407), .A3(new_n317), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(new_n613), .A3(new_n679), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  NOR3_X1   g542(.A1(new_n721), .A2(new_n724), .A3(new_n648), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n690), .A2(new_n613), .A3(new_n708), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n611), .B1(new_n308), .B2(new_n309), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n307), .A2(new_n733), .A3(new_n313), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n659), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n543), .A2(new_n735), .A3(new_n595), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n472), .A2(new_n476), .ZN(new_n737));
  INV_X1    g551(.A(new_n622), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n667), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n732), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT32), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n540), .B2(new_n541), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n742), .A2(new_n533), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n712), .B1(new_n743), .B2(new_n522), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(KEYINPUT42), .A3(new_n690), .A4(new_n735), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n740), .A2(new_n745), .A3(KEYINPUT105), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n327), .ZN(G33));
  AND2_X1   g565(.A1(new_n735), .A2(new_n595), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(KEYINPUT106), .A3(new_n543), .A4(new_n670), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT106), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n736), .B2(new_n668), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n319), .ZN(G36));
  NAND3_X1  g571(.A1(new_n472), .A2(new_n738), .A3(new_n476), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n758), .B(KEYINPUT43), .Z(new_n759));
  NOR2_X1   g573(.A1(new_n604), .A2(new_n648), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n734), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n759), .A2(KEYINPUT44), .A3(new_n760), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n361), .A2(KEYINPUT45), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n361), .A2(KEYINPUT45), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(G469), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(KEYINPUT46), .A3(new_n657), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT107), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n770), .A2(new_n771), .A3(new_n366), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n771), .B1(new_n770), .B2(new_n366), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT46), .B1(new_n769), .B2(new_n657), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n674), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n775), .A2(new_n317), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n766), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n764), .B1(new_n763), .B2(new_n765), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  OR3_X1    g596(.A1(new_n775), .A2(new_n782), .A3(new_n317), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n782), .B1(new_n775), .B2(new_n317), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT109), .ZN(new_n786));
  NOR4_X1   g600(.A1(new_n739), .A2(new_n543), .A3(new_n595), .A4(new_n734), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n786), .B1(new_n785), .B2(new_n787), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  NAND2_X1  g605(.A1(new_n691), .A2(new_n730), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n672), .A2(new_n792), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n679), .A2(new_n633), .A3(new_n634), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n594), .A2(new_n647), .A3(new_n689), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n316), .B(new_n795), .C1(new_n653), .C2(new_n658), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n362), .A2(new_n366), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(KEYINPUT113), .A3(new_n316), .A4(new_n795), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n798), .A2(new_n686), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n794), .A2(new_n801), .A3(KEYINPUT114), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n679), .A2(new_n633), .A3(new_n634), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n798), .A2(new_n686), .A3(new_n800), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(new_n793), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n661), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n668), .A2(new_n609), .A3(new_n612), .A4(new_n662), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT98), .B1(new_n613), .B2(new_n670), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n691), .A2(new_n730), .ZN(new_n813));
  AND4_X1   g627(.A1(KEYINPUT52), .A2(new_n807), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n808), .A2(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n740), .A2(KEYINPUT105), .A3(new_n745), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT105), .B1(new_n740), .B2(new_n745), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n314), .A2(new_n607), .A3(new_n368), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n472), .A2(new_n476), .A3(new_n402), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n604), .A2(new_n819), .A3(new_n605), .A4(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n650), .A2(new_n821), .A3(KEYINPUT110), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT110), .B1(new_n650), .B2(new_n821), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n604), .A2(new_n819), .A3(new_n623), .A4(new_n605), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n596), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n729), .A2(new_n735), .A3(new_n623), .A4(new_n667), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n397), .A2(new_n476), .A3(new_n401), .A4(new_n667), .ZN(new_n828));
  INV_X1    g642(.A(new_n467), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n466), .B1(new_n461), .B2(new_n463), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n828), .B1(new_n831), .B2(new_n628), .ZN(new_n832));
  INV_X1    g646(.A(new_n734), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n543), .A2(new_n832), .A3(new_n660), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n827), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n753), .B2(new_n755), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n698), .A2(new_n709), .A3(new_n727), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n704), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n818), .A2(new_n826), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT53), .B1(new_n815), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n661), .A2(new_n663), .A3(new_n739), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n841), .B(new_n842), .C1(new_n806), .C2(new_n802), .ZN(new_n843));
  INV_X1    g657(.A(new_n730), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n672), .A2(KEYINPUT112), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT112), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n812), .B2(new_n730), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n843), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n807), .A2(new_n813), .A3(new_n812), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n841), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n838), .A2(new_n836), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n650), .A2(new_n821), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT110), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n650), .A2(new_n821), .A3(KEYINPUT110), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n596), .A3(new_n856), .A4(new_n824), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n852), .A2(new_n750), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n851), .B1(new_n858), .B2(KEYINPUT111), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT111), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n860), .B1(new_n839), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n840), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n793), .A2(KEYINPUT52), .A3(new_n807), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n850), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT53), .B1(new_n858), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT112), .B1(new_n672), .B2(new_n844), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n812), .A2(new_n846), .A3(new_n730), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n871), .A2(new_n843), .B1(new_n841), .B2(new_n849), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n860), .B1(new_n740), .B2(new_n745), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n836), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n697), .B1(new_n636), .B2(new_n639), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n698), .A2(new_n709), .A3(new_n727), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT115), .B1(new_n704), .B2(new_n837), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n874), .A2(new_n826), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n868), .A2(new_n881), .A3(KEYINPUT54), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n865), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n759), .A2(new_n404), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n734), .A2(new_n707), .A3(new_n317), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n729), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n686), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n885), .A2(new_n887), .A3(new_n404), .A4(new_n595), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n472), .A2(new_n476), .A3(new_n622), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n884), .A2(new_n725), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n681), .A2(new_n368), .A3(new_n317), .A4(new_n707), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT50), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n891), .A2(KEYINPUT50), .A3(new_n892), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n707), .A2(new_n316), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n833), .B(new_n891), .C1(new_n785), .C2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(KEYINPUT51), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n884), .A2(new_n744), .A3(new_n885), .ZN(new_n901));
  XOR2_X1   g715(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n902));
  OR2_X1    g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  INV_X1    g718(.A(new_n623), .ZN(new_n905));
  OAI211_X1 g719(.A(G952), .B(new_n343), .C1(new_n888), .C2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n613), .A2(new_n708), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n891), .B2(new_n908), .ZN(new_n909));
  AND4_X1   g723(.A1(new_n900), .A2(new_n903), .A3(new_n904), .A4(new_n909), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n899), .A2(KEYINPUT116), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n899), .A2(KEYINPUT116), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n911), .A2(new_n897), .A3(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n883), .B(new_n910), .C1(KEYINPUT51), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n403), .A2(new_n343), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT118), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n681), .A2(new_n758), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n712), .A2(new_n611), .A3(new_n317), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n707), .B(KEYINPUT49), .Z(new_n920));
  NAND4_X1  g734(.A1(new_n918), .A2(new_n887), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n917), .A2(new_n921), .ZN(G75));
  NOR2_X1   g736(.A1(new_n343), .A2(G952), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n877), .B1(new_n875), .B2(new_n876), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n704), .A2(new_n837), .A3(KEYINPUT115), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n836), .A2(new_n873), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n851), .A2(new_n826), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n860), .B1(new_n815), .B2(new_n839), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(G902), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT56), .B1(new_n933), .B2(G210), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n249), .A2(new_n251), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(new_n279), .Z(new_n936));
  XNOR2_X1  g750(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n924), .B1(new_n934), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n934), .B2(new_n939), .ZN(G51));
  OAI21_X1  g755(.A(KEYINPUT54), .B1(new_n868), .B2(new_n881), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n929), .A2(new_n930), .A3(new_n864), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n657), .B(KEYINPUT57), .Z(new_n945));
  AOI21_X1  g759(.A(new_n693), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n932), .A2(new_n769), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n924), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT120), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(KEYINPUT120), .B(new_n924), .C1(new_n946), .C2(new_n947), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(G54));
  NAND3_X1  g766(.A1(new_n933), .A2(KEYINPUT58), .A3(G475), .ZN(new_n953));
  INV_X1    g767(.A(new_n627), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n955), .A2(new_n956), .A3(new_n923), .ZN(G60));
  INV_X1    g771(.A(KEYINPUT123), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT122), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n617), .A2(new_n618), .ZN(new_n960));
  XNOR2_X1  g774(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(new_n620), .Z(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n864), .B1(new_n929), .B2(new_n930), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n959), .B(new_n964), .C1(new_n882), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n924), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n959), .B1(new_n944), .B2(new_n964), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n958), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n964), .B1(new_n882), .B2(new_n965), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT122), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n971), .A2(KEYINPUT123), .A3(new_n924), .A4(new_n966), .ZN(new_n972));
  INV_X1    g786(.A(new_n962), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n618), .B(new_n617), .C1(new_n883), .C2(new_n973), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n969), .A2(new_n972), .A3(new_n974), .ZN(G63));
  XNOR2_X1  g789(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n370), .A2(new_n281), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n931), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(new_n587), .A3(new_n586), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n931), .A2(new_n646), .A3(new_n978), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n980), .A2(new_n924), .A3(new_n981), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n406), .B2(new_n277), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n826), .A2(new_n838), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n984), .B1(new_n986), .B2(G953), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n935), .B1(G898), .B2(new_n343), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G69));
  AOI21_X1  g803(.A(new_n343), .B1(G227), .B2(G900), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n736), .A2(new_n776), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n623), .B2(new_n820), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n780), .B(new_n992), .C1(new_n788), .C2(new_n789), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n842), .B1(new_n869), .B2(new_n870), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n687), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT62), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n343), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n509), .B1(new_n525), .B2(new_n526), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(new_n449), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT127), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n750), .A2(new_n756), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n1002), .A2(KEYINPUT126), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n777), .A2(new_n794), .A3(new_n744), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n994), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1002), .A2(KEYINPUT126), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  OAI22_X1  g821(.A1(new_n788), .A2(new_n789), .B1(new_n779), .B2(new_n778), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n1007), .A2(new_n1008), .A3(G953), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n999), .B1(G900), .B2(G953), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1001), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1000), .A2(new_n1012), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1009), .A2(new_n1001), .A3(new_n1011), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n990), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n990), .B(KEYINPUT125), .Z(new_n1016));
  OAI211_X1 g830(.A(new_n1000), .B(new_n1016), .C1(new_n1009), .C2(new_n1011), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1015), .A2(new_n1017), .ZN(G72));
  NAND2_X1  g832(.A1(G472), .A2(G902), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT63), .Z(new_n1020));
  OR2_X1    g834(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1020), .B1(new_n1021), .B2(new_n985), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n527), .A2(new_n488), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1023), .A2(new_n501), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1023), .A2(new_n501), .ZN(new_n1026));
  OR3_X1    g840(.A1(new_n993), .A2(new_n985), .A3(new_n996), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1026), .B1(new_n1027), .B2(new_n1020), .ZN(new_n1028));
  INV_X1    g842(.A(new_n517), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1020), .B1(new_n1029), .B2(new_n682), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n924), .B1(new_n863), .B2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g845(.A1(new_n1025), .A2(new_n1028), .A3(new_n1031), .ZN(G57));
endmodule


