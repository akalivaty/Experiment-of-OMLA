//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1027, new_n1028,
    new_n1029, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1046, new_n1047, new_n1048, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT13), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT92), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT15), .ZN(new_n205));
  INV_X1    g004(.A(G43gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G50gat), .ZN(new_n207));
  INV_X1    g006(.A(G50gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G43gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n205), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(G43gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n206), .A2(G50gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT15), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT14), .ZN(new_n218));
  INV_X1    g017(.A(G29gat), .ZN(new_n219));
  INV_X1    g018(.A(G36gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT91), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(KEYINPUT91), .A3(new_n220), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n217), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n204), .B1(new_n215), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n225), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT91), .B1(new_n224), .B2(new_n220), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n216), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G43gat), .B(G50gat), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n231), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n230), .A2(KEYINPUT92), .A3(new_n210), .A4(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G8gat), .ZN(new_n235));
  INV_X1    g034(.A(G22gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G15gat), .ZN(new_n237));
  INV_X1    g036(.A(G15gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G22gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT16), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n237), .B(new_n239), .C1(new_n240), .C2(G1gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT93), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n235), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G15gat), .B(G22gat), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n241), .B1(G1gat), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI221_X1 g045(.A(new_n241), .B1(new_n242), .B2(new_n235), .C1(G1gat), .C2(new_n244), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n221), .A2(new_n216), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n214), .B1(new_n249), .B2(new_n211), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n234), .A2(new_n248), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n248), .B1(new_n251), .B2(new_n234), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n203), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G197gat), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT11), .B(G169gat), .Z(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT12), .ZN(new_n259));
  INV_X1    g058(.A(new_n248), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n234), .A2(new_n251), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT17), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n250), .B1(new_n227), .B2(new_n233), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT17), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n260), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(KEYINPUT18), .B(new_n202), .C1(new_n263), .C2(new_n248), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n254), .B(new_n259), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n263), .A2(new_n264), .ZN(new_n269));
  AOI211_X1 g068(.A(KEYINPUT17), .B(new_n250), .C1(new_n227), .C2(new_n233), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n248), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n202), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n253), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT18), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT94), .B1(new_n268), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n273), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT18), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT12), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n258), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n263), .B(new_n248), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n280), .B1(new_n281), .B2(new_n203), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT94), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n271), .A2(KEYINPUT18), .A3(new_n273), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n278), .A2(new_n282), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n278), .A2(new_n284), .A3(new_n254), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n275), .A2(new_n285), .B1(new_n286), .B2(new_n280), .ZN(new_n287));
  XOR2_X1   g086(.A(G211gat), .B(G218gat), .Z(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT75), .B(G197gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G204gat), .ZN(new_n291));
  INV_X1    g090(.A(G204gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT75), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(G197gat), .ZN(new_n294));
  INV_X1    g093(.A(G197gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(KEYINPUT75), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n292), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT22), .ZN(new_n299));
  INV_X1    g098(.A(G211gat), .ZN(new_n300));
  INV_X1    g099(.A(G218gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n289), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n298), .A2(new_n289), .A3(new_n302), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n307));
  INV_X1    g106(.A(G226gat), .ZN(new_n308));
  INV_X1    g107(.A(G233gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT67), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT25), .ZN(new_n312));
  INV_X1    g111(.A(G169gat), .ZN(new_n313));
  INV_X1    g112(.A(G176gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT23), .ZN(new_n319));
  NAND2_X1  g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT65), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n317), .A2(new_n318), .A3(new_n319), .A4(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(G183gat), .B2(G190gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT24), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n325), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n311), .B1(new_n323), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n328), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT24), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(new_n326), .ZN(new_n334));
  NOR2_X1   g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335));
  AND2_X1   g134(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(G190gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n319), .A2(new_n322), .A3(new_n318), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n338), .A2(KEYINPUT67), .A3(new_n339), .A4(new_n317), .ZN(new_n340));
  AND2_X1   g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n341), .B1(new_n315), .B2(new_n316), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n333), .ZN(new_n343));
  OR2_X1    g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n344), .A3(new_n324), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT64), .B(G176gat), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n342), .B(new_n345), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(new_n312), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n331), .A2(new_n340), .A3(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n315), .A2(KEYINPUT26), .ZN(new_n351));
  NOR2_X1   g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT26), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n320), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n327), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT27), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(KEYINPUT68), .A3(G183gat), .ZN(new_n358));
  AND2_X1   g157(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n356), .B(new_n358), .C1(new_n359), .C2(new_n357), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT27), .B(G183gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(KEYINPUT28), .A3(new_n356), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n355), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n310), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n310), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n370), .B1(new_n350), .B2(new_n366), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n307), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n338), .A2(new_n317), .A3(new_n339), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n373), .A2(new_n311), .B1(new_n348), .B2(new_n312), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n365), .B1(new_n374), .B2(new_n340), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n370), .B1(new_n375), .B2(KEYINPUT29), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT76), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n306), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n306), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n369), .A2(new_n379), .A3(new_n371), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT37), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G8gat), .B(G36gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(G64gat), .B(G92gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(KEYINPUT89), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n371), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT76), .B1(new_n376), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n369), .A2(new_n307), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n379), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT37), .ZN(new_n391));
  INV_X1    g190(.A(new_n380), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT89), .B1(new_n381), .B2(new_n385), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT38), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397));
  XOR2_X1   g196(.A(KEYINPUT72), .B(G120gat), .Z(new_n398));
  INV_X1    g197(.A(G113gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT73), .B(G113gat), .ZN(new_n400));
  INV_X1    g199(.A(G120gat), .ZN(new_n401));
  OAI22_X1  g200(.A1(new_n398), .A2(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G127gat), .ZN(new_n403));
  INV_X1    g202(.A(G134gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(G127gat), .A2(G134gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT1), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n402), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n403), .A2(KEYINPUT69), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT69), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(G127gat), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n404), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT70), .B1(new_n414), .B2(new_n407), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT70), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT69), .B(G127gat), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n416), .B(new_n408), .C1(new_n417), .C2(new_n404), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n399), .A2(new_n401), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT1), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n421), .B1(G113gat), .B2(G120gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT71), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT71), .ZN(new_n426));
  AOI211_X1 g225(.A(new_n426), .B(new_n423), .C1(new_n415), .C2(new_n418), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n410), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G155gat), .ZN(new_n429));
  OR2_X1    g228(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT2), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT80), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT78), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n429), .A2(G162gat), .ZN(new_n436));
  INV_X1    g235(.A(G162gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n437), .A2(G155gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n435), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(G155gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n429), .A2(G162gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT78), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(G141gat), .B(G148gat), .Z(new_n444));
  AND2_X1   g243(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n446));
  OAI21_X1  g245(.A(G155gat), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT80), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT2), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n434), .A2(new_n443), .A3(new_n444), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n444), .A2(new_n433), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(new_n436), .B2(new_n438), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n397), .B1(new_n428), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n412), .A2(G127gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n403), .A2(KEYINPUT69), .ZN(new_n456));
  OAI21_X1  g255(.A(G134gat), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n416), .B1(new_n457), .B2(new_n408), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n414), .A2(KEYINPUT70), .A3(new_n407), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n424), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n426), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n419), .A2(KEYINPUT71), .A3(new_n424), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n453), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n463), .A2(KEYINPUT4), .A3(new_n464), .A4(new_n410), .ZN(new_n465));
  NAND2_X1  g264(.A1(G225gat), .A2(G233gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n454), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n469), .A3(new_n452), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n428), .A2(new_n470), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n450), .A2(KEYINPUT81), .A3(new_n452), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT81), .B1(new_n450), .B2(new_n452), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n472), .A2(new_n473), .A3(new_n469), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n468), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT81), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n453), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n450), .A2(KEYINPUT81), .A3(new_n452), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(KEYINPUT3), .A3(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n479), .A2(KEYINPUT82), .A3(new_n470), .A4(new_n428), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n467), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n464), .B(new_n410), .C1(new_n425), .C2(new_n427), .ZN(new_n482));
  INV_X1    g281(.A(new_n428), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n477), .A2(new_n478), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n466), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT5), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT83), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n481), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n480), .ZN(new_n491));
  INV_X1    g290(.A(new_n467), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT5), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n494), .B1(new_n485), .B2(new_n486), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT83), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  OAI22_X1  g295(.A1(new_n490), .A2(new_n496), .B1(KEYINPUT5), .B2(new_n493), .ZN(new_n497));
  XOR2_X1   g296(.A(G1gat), .B(G29gat), .Z(new_n498));
  XNOR2_X1  g297(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G57gat), .B(G85gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n502), .A2(new_n503), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n497), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT88), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n379), .B1(new_n372), .B2(new_n377), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n376), .A2(new_n387), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT37), .B1(new_n510), .B2(new_n306), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n508), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n306), .B1(new_n388), .B2(new_n389), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n369), .A2(new_n371), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n391), .B1(new_n514), .B2(new_n379), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(KEYINPUT88), .A3(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n384), .A2(KEYINPUT38), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n393), .A2(new_n512), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n390), .A2(new_n384), .A3(new_n392), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT77), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n390), .A2(KEYINPUT77), .A3(new_n384), .A4(new_n392), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n518), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n489), .B1(new_n481), .B2(new_n488), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n493), .A2(KEYINPUT83), .A3(new_n495), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(new_n503), .A3(new_n502), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n396), .A2(new_n507), .A3(new_n523), .A4(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT86), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n485), .B2(new_n486), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n472), .A2(new_n473), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n428), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n533), .A2(KEYINPUT86), .A3(new_n466), .A4(new_n482), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(KEYINPUT39), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT87), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n454), .A2(new_n465), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n491), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n486), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT87), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n531), .A2(new_n540), .A3(KEYINPUT39), .A4(new_n534), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n536), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n466), .B1(new_n491), .B2(new_n537), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT39), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n502), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT40), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n497), .A2(new_n502), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT30), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n521), .A2(new_n522), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n384), .B1(new_n390), .B2(new_n392), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n378), .A2(new_n385), .A3(new_n380), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n552), .B1(KEYINPUT30), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n542), .A2(KEYINPUT40), .A3(new_n545), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n548), .A2(new_n549), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n305), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n368), .B1(new_n558), .B2(new_n303), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n464), .B1(new_n559), .B2(new_n469), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n306), .B1(new_n368), .B2(new_n470), .ZN(new_n561));
  INV_X1    g360(.A(G228gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(new_n309), .ZN(new_n563));
  NOR3_X1   g362(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT29), .B1(new_n304), .B2(new_n305), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n477), .B(new_n478), .C1(new_n566), .C2(KEYINPUT3), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n470), .A2(new_n368), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n379), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n565), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(G22gat), .B1(new_n564), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n559), .A2(new_n469), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n453), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(new_n565), .A3(new_n569), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n561), .B1(new_n532), .B2(new_n572), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n574), .B(new_n236), .C1(new_n575), .C2(new_n565), .ZN(new_n576));
  XNOR2_X1  g375(.A(G78gat), .B(G106gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT31), .B(G50gat), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n577), .B(new_n578), .Z(new_n579));
  INV_X1    g378(.A(KEYINPUT85), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n571), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n571), .A2(new_n576), .B1(new_n580), .B2(new_n579), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n529), .A2(new_n557), .A3(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n551), .A2(new_n554), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n506), .B1(new_n497), .B2(new_n505), .ZN(new_n588));
  INV_X1    g387(.A(new_n506), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n527), .A2(new_n504), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n587), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n584), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n463), .A2(new_n367), .A3(new_n410), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n428), .A2(new_n375), .ZN(new_n595));
  NAND2_X1  g394(.A1(G227gat), .A2(G233gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G71gat), .B(G99gat), .Z(new_n599));
  XNOR2_X1  g398(.A(G15gat), .B(G43gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT33), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n598), .A2(KEYINPUT32), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT74), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT74), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n598), .A2(new_n605), .A3(KEYINPUT32), .A4(new_n602), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n597), .B1(new_n594), .B2(new_n595), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT34), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n598), .A2(KEYINPUT32), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n598), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n612), .A3(new_n601), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n607), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n609), .B1(new_n607), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n593), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n607), .A2(new_n613), .ZN(new_n617));
  INV_X1    g416(.A(new_n609), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n607), .A2(new_n609), .A3(new_n613), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(KEYINPUT36), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n586), .A2(new_n592), .A3(new_n622), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n584), .A2(new_n614), .A3(new_n615), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n587), .B(new_n624), .C1(new_n588), .C2(new_n590), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT35), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n555), .B1(new_n507), .B2(new_n528), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT90), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n614), .B2(new_n615), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n619), .A2(KEYINPUT90), .A3(new_n620), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n584), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT35), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n627), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n626), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n287), .B1(new_n623), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n588), .A2(new_n590), .ZN(new_n636));
  OR2_X1    g435(.A1(G99gat), .A2(G106gat), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n638));
  NAND2_X1  g437(.A1(G99gat), .A2(G106gat), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AND3_X1   g439(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(G99gat), .A2(G106gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(G99gat), .A2(G106gat), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT96), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(G85gat), .ZN(new_n647));
  INV_X1    g446(.A(G92gat), .ZN(new_n648));
  AOI22_X1  g447(.A1(KEYINPUT8), .A2(new_n639), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n640), .A2(new_n643), .A3(new_n646), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n639), .A2(KEYINPUT8), .ZN(new_n651));
  NAND2_X1  g450(.A1(G85gat), .A2(G92gat), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT7), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n647), .A2(new_n648), .ZN(new_n655));
  NAND3_X1  g454(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n651), .A2(new_n654), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT96), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n638), .B1(new_n637), .B2(new_n639), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n650), .B(new_n660), .C1(new_n269), .C2(new_n270), .ZN(new_n661));
  AND3_X1   g460(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n650), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(new_n261), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(G190gat), .B(G218gat), .Z(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  XNOR2_X1  g468(.A(G134gat), .B(G162gat), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n670), .B(new_n671), .Z(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n673), .A2(KEYINPUT97), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(KEYINPUT97), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n668), .B(new_n669), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n668), .A2(new_n669), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n676), .B1(new_n677), .B2(new_n675), .ZN(new_n678));
  NAND2_X1  g477(.A1(G71gat), .A2(G78gat), .ZN(new_n679));
  OR2_X1    g478(.A1(G71gat), .A2(G78gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(G57gat), .B(G64gat), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT9), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n679), .B(new_n680), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n679), .ZN(new_n684));
  INV_X1    g483(.A(G57gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G64gat), .ZN(new_n686));
  INV_X1    g485(.A(G64gat), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G57gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n679), .A2(new_n682), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n684), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT21), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(G231gat), .A2(G233gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G127gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n248), .B1(new_n693), .B2(new_n692), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(G183gat), .B(G211gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT95), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(new_n429), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n701), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n699), .B(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n678), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(G120gat), .B(G148gat), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT100), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT101), .ZN(new_n709));
  XNOR2_X1  g508(.A(G176gat), .B(G204gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n683), .A2(new_n691), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n663), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT10), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n692), .A2(new_n650), .A3(new_n660), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT98), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT98), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n714), .A2(new_n719), .A3(new_n715), .A4(new_n716), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT99), .B1(new_n714), .B2(new_n715), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT99), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n663), .A2(new_n713), .A3(new_n722), .A4(KEYINPUT10), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n718), .A2(new_n720), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(G230gat), .A2(G233gat), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n714), .A2(new_n716), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n726), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n712), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n729), .B(new_n711), .C1(new_n724), .C2(new_n726), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n706), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n635), .A2(new_n636), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g537(.A1(new_n735), .A2(new_n587), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT16), .B(G8gat), .Z(new_n740));
  AND3_X1   g539(.A1(new_n635), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n235), .B1(new_n635), .B2(new_n739), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT42), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(KEYINPUT42), .B2(new_n741), .ZN(G1325gat));
  NAND2_X1  g543(.A1(new_n635), .A2(new_n736), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n616), .A2(new_n621), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n616), .B2(new_n621), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G15gat), .B1(new_n745), .B2(new_n749), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n614), .A2(new_n615), .A3(new_n628), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT90), .B1(new_n619), .B2(new_n620), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n635), .A2(new_n238), .A3(new_n754), .A4(new_n736), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n750), .A2(new_n755), .ZN(G1326gat));
  NOR2_X1   g555(.A1(new_n745), .A2(new_n585), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT43), .B(G22gat), .Z(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1327gat));
  NAND2_X1  g558(.A1(new_n678), .A2(KEYINPUT44), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(new_n623), .B2(new_n634), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n287), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n705), .A3(new_n734), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n678), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n586), .A2(new_n749), .A3(new_n592), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(new_n634), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n762), .B(new_n765), .C1(KEYINPUT44), .C2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n636), .ZN(new_n770));
  OAI21_X1  g569(.A(G29gat), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n764), .A2(new_n766), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n623), .B2(new_n634), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(new_n219), .A3(new_n636), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT45), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n771), .A2(new_n776), .ZN(G1328gat));
  NAND3_X1  g576(.A1(new_n774), .A2(new_n220), .A3(new_n555), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT46), .Z(new_n779));
  OAI21_X1  g578(.A(G36gat), .B1(new_n769), .B2(new_n587), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(G1329gat));
  OAI21_X1  g580(.A(G43gat), .B1(new_n769), .B2(new_n749), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n774), .A2(new_n206), .A3(new_n754), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g584(.A(KEYINPUT48), .ZN(new_n786));
  OAI21_X1  g585(.A(G50gat), .B1(new_n769), .B2(new_n585), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n585), .A2(G50gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n774), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n786), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(KEYINPUT103), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT103), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n774), .A2(new_n792), .A3(new_n788), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(new_n786), .A3(new_n793), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n529), .A2(new_n557), .A3(new_n585), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n614), .A2(new_n615), .A3(new_n593), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT36), .B1(new_n619), .B2(new_n620), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT102), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n616), .A2(new_n621), .A3(new_n746), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n798), .B(new_n799), .C1(new_n627), .C2(new_n585), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n632), .B(new_n587), .C1(new_n588), .C2(new_n590), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n585), .B1(new_n751), .B2(new_n752), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n632), .B1(new_n627), .B2(new_n624), .ZN(new_n804));
  OAI22_X1  g603(.A1(new_n795), .A2(new_n800), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT44), .B1(new_n805), .B2(new_n678), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n761), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(new_n584), .A3(new_n765), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n794), .B1(new_n808), .B2(G50gat), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT104), .B1(new_n790), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n793), .A2(new_n786), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n787), .A2(new_n791), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT104), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n808), .A2(G50gat), .B1(new_n774), .B2(new_n788), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n812), .B(new_n813), .C1(new_n814), .C2(new_n786), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n810), .A2(new_n815), .ZN(G1331gat));
  AND2_X1   g615(.A1(new_n767), .A2(new_n634), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n706), .A2(new_n287), .A3(new_n733), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n636), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(G57gat), .ZN(G1332gat));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT105), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n819), .B(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n587), .A2(KEYINPUT106), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n587), .A2(KEYINPUT106), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n827), .B1(new_n828), .B2(new_n687), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT107), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n822), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n817), .A2(new_n818), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n823), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n819), .A2(KEYINPUT105), .ZN(new_n834));
  AND4_X1   g633(.A1(new_n822), .A2(new_n833), .A3(new_n834), .A4(new_n830), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n831), .A2(new_n835), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n824), .A2(new_n822), .A3(new_n830), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n833), .A2(new_n834), .A3(new_n830), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT108), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n837), .A2(new_n839), .A3(new_n828), .A4(new_n687), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n836), .A2(new_n840), .ZN(G1333gat));
  INV_X1    g640(.A(KEYINPUT50), .ZN(new_n842));
  INV_X1    g641(.A(new_n749), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n833), .A2(new_n843), .A3(new_n834), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(G71gat), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n832), .A2(G71gat), .A3(new_n753), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n842), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  AOI211_X1 g647(.A(KEYINPUT50), .B(new_n846), .C1(new_n844), .C2(G71gat), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(G1334gat));
  NAND2_X1  g649(.A1(new_n824), .A2(new_n584), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(G78gat), .ZN(G1335gat));
  INV_X1    g651(.A(new_n705), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(new_n763), .ZN(new_n854));
  AND4_X1   g653(.A1(KEYINPUT51), .A2(new_n805), .A3(new_n678), .A4(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT51), .B1(new_n768), .B2(new_n854), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n857), .A2(new_n647), .A3(new_n636), .A4(new_n733), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n854), .A2(new_n733), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n762), .B(new_n860), .C1(KEYINPUT44), .C2(new_n768), .ZN(new_n861));
  OAI21_X1  g660(.A(G85gat), .B1(new_n861), .B2(new_n770), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n858), .A2(new_n862), .ZN(G1336gat));
  INV_X1    g662(.A(KEYINPUT109), .ZN(new_n864));
  NOR4_X1   g663(.A1(new_n806), .A2(new_n587), .A3(new_n761), .A4(new_n859), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(new_n648), .ZN(new_n866));
  OAI211_X1 g665(.A(KEYINPUT109), .B(G92gat), .C1(new_n861), .C2(new_n587), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n825), .A2(new_n826), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(G92gat), .A3(new_n734), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT110), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n870), .B1(new_n855), .B2(new_n856), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT111), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(KEYINPUT111), .B(new_n870), .C1(new_n855), .C2(new_n856), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n866), .A2(new_n867), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT52), .ZN(new_n876));
  OAI21_X1  g675(.A(G92gat), .B1(new_n861), .B2(new_n868), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n878), .A3(new_n871), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n876), .A2(new_n879), .ZN(G1337gat));
  NOR3_X1   g679(.A1(new_n753), .A2(G99gat), .A3(new_n734), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n857), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G99gat), .B1(new_n861), .B2(new_n749), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1338gat));
  OAI21_X1  g683(.A(G106gat), .B1(new_n861), .B2(new_n585), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT112), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n585), .A2(G106gat), .A3(new_n734), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n890), .B1(new_n855), .B2(new_n856), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n885), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n886), .A2(new_n887), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n892), .B(new_n893), .ZN(G1339gat));
  INV_X1    g693(.A(new_n732), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT55), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n718), .A2(new_n720), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n721), .A2(new_n723), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n725), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n725), .B1(new_n721), .B2(new_n723), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n896), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n711), .B1(new_n727), .B2(new_n901), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n895), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n899), .A2(new_n901), .A3(new_n725), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n897), .A2(new_n902), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n907), .B(new_n712), .C1(new_n909), .C2(new_n727), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n896), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n272), .B1(new_n266), .B2(new_n253), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(new_n281), .B2(new_n203), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n285), .A2(new_n275), .B1(new_n914), .B2(new_n258), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n678), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n912), .A2(new_n763), .B1(new_n733), .B2(new_n915), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(new_n678), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n705), .A2(new_n918), .B1(new_n736), .B2(new_n287), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(new_n802), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n827), .A2(new_n770), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(G113gat), .B1(new_n922), .B2(new_n287), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n918), .A2(new_n705), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n736), .A2(new_n287), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n636), .ZN(new_n927));
  INV_X1    g726(.A(new_n624), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n868), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n287), .A2(new_n400), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(G1340gat));
  OAI21_X1  g731(.A(G120gat), .B1(new_n922), .B2(new_n734), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n734), .A2(new_n398), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT113), .Z(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n930), .B2(new_n935), .ZN(G1341gat));
  NAND3_X1  g735(.A1(new_n929), .A2(new_n853), .A3(new_n868), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT115), .ZN(new_n938));
  AOI211_X1 g737(.A(new_n455), .B(new_n456), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n922), .A2(new_n417), .A3(new_n705), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT114), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  AOI22_X1  g743(.A1(new_n939), .A2(new_n940), .B1(new_n943), .B2(new_n944), .ZN(G1342gat));
  NOR2_X1   g744(.A1(new_n766), .A2(new_n555), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n404), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n922), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n404), .B1(new_n948), .B2(new_n678), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n947), .B1(new_n949), .B2(KEYINPUT56), .ZN(new_n950));
  OR3_X1    g749(.A1(new_n947), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT116), .B1(new_n947), .B2(KEYINPUT56), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT117), .ZN(G1343gat));
  NAND2_X1  g753(.A1(new_n749), .A2(new_n584), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n927), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n287), .A2(G141gat), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n868), .A3(new_n957), .ZN(new_n958));
  XOR2_X1   g757(.A(new_n958), .B(KEYINPUT120), .Z(new_n959));
  INV_X1    g758(.A(G141gat), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n921), .A2(new_n749), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT57), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n962), .B1(new_n919), .B2(new_n585), .ZN(new_n963));
  INV_X1    g762(.A(new_n916), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n285), .A2(new_n275), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n914), .A2(new_n258), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n965), .A2(new_n733), .A3(new_n966), .ZN(new_n967));
  XNOR2_X1  g766(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n910), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n906), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n970), .B2(new_n287), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT119), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n678), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n967), .B(KEYINPUT119), .C1(new_n970), .C2(new_n287), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n964), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n925), .B1(new_n975), .B2(new_n853), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n585), .A2(new_n962), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n961), .B1(new_n963), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n960), .B1(new_n979), .B2(new_n763), .ZN(new_n980));
  OAI21_X1  g779(.A(KEYINPUT58), .B1(new_n959), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n956), .A2(new_n868), .ZN(new_n982));
  INV_X1    g781(.A(new_n957), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(KEYINPUT58), .B1(new_n984), .B2(KEYINPUT121), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n985), .B1(KEYINPUT121), .B2(new_n984), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n981), .B1(new_n980), .B2(new_n986), .ZN(G1344gat));
  INV_X1    g786(.A(G148gat), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n956), .A2(new_n988), .A3(new_n733), .A4(new_n868), .ZN(new_n989));
  XNOR2_X1  g788(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n961), .A2(new_n734), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n705), .B1(new_n975), .B2(KEYINPUT123), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT123), .ZN(new_n993));
  AOI211_X1 g792(.A(new_n993), .B(new_n964), .C1(new_n973), .C2(new_n974), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n925), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g794(.A(KEYINPUT57), .B1(new_n995), .B2(new_n584), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n926), .A2(new_n977), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n991), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n990), .B1(new_n998), .B2(G148gat), .ZN(new_n999));
  AOI211_X1 g798(.A(KEYINPUT59), .B(new_n988), .C1(new_n979), .C2(new_n733), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n989), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT124), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g802(.A(KEYINPUT124), .B(new_n989), .C1(new_n999), .C2(new_n1000), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(G1345gat));
  NAND3_X1  g804(.A1(new_n956), .A2(new_n853), .A3(new_n868), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n705), .A2(new_n429), .ZN(new_n1007));
  XNOR2_X1  g806(.A(new_n1007), .B(KEYINPUT125), .ZN(new_n1008));
  AOI22_X1  g807(.A1(new_n1006), .A2(new_n429), .B1(new_n979), .B2(new_n1008), .ZN(G1346gat));
  NOR2_X1   g808(.A1(new_n445), .A2(new_n446), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n956), .A2(new_n1010), .A3(new_n946), .ZN(new_n1011));
  AND2_X1   g810(.A1(new_n979), .A2(new_n678), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1011), .B1(new_n1012), .B2(new_n1010), .ZN(new_n1013));
  XOR2_X1   g812(.A(new_n1013), .B(KEYINPUT126), .Z(G1347gat));
  NAND2_X1  g813(.A1(new_n770), .A2(new_n555), .ZN(new_n1015));
  XNOR2_X1  g814(.A(new_n1015), .B(KEYINPUT127), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1016), .A2(new_n920), .ZN(new_n1017));
  NOR3_X1   g816(.A1(new_n1017), .A2(new_n313), .A3(new_n287), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n926), .A2(new_n770), .ZN(new_n1019));
  NOR3_X1   g818(.A1(new_n1019), .A2(new_n928), .A3(new_n868), .ZN(new_n1020));
  AOI21_X1  g819(.A(G169gat), .B1(new_n1020), .B2(new_n763), .ZN(new_n1021));
  NOR2_X1   g820(.A1(new_n1018), .A2(new_n1021), .ZN(G1348gat));
  AOI21_X1  g821(.A(G176gat), .B1(new_n1020), .B2(new_n733), .ZN(new_n1023));
  INV_X1    g822(.A(new_n1017), .ZN(new_n1024));
  AND2_X1   g823(.A1(new_n733), .A2(new_n347), .ZN(new_n1025));
  AOI21_X1  g824(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(G1349gat));
  OAI21_X1  g825(.A(G183gat), .B1(new_n1017), .B2(new_n705), .ZN(new_n1027));
  NAND3_X1  g826(.A1(new_n1020), .A2(new_n363), .A3(new_n853), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g828(.A(new_n1029), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g829(.A1(new_n1020), .A2(new_n356), .A3(new_n678), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n1024), .A2(new_n678), .ZN(new_n1032));
  INV_X1    g831(.A(KEYINPUT61), .ZN(new_n1033));
  NAND3_X1  g832(.A1(new_n1032), .A2(new_n1033), .A3(G190gat), .ZN(new_n1034));
  INV_X1    g833(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g834(.A(new_n1033), .B1(new_n1032), .B2(G190gat), .ZN(new_n1036));
  OAI21_X1  g835(.A(new_n1031), .B1(new_n1035), .B2(new_n1036), .ZN(G1351gat));
  NOR3_X1   g836(.A1(new_n1019), .A2(new_n868), .A3(new_n955), .ZN(new_n1038));
  AOI21_X1  g837(.A(G197gat), .B1(new_n1038), .B2(new_n763), .ZN(new_n1039));
  OR2_X1    g838(.A1(new_n996), .A2(new_n997), .ZN(new_n1040));
  AND2_X1   g839(.A1(new_n1016), .A2(new_n749), .ZN(new_n1041));
  NAND2_X1  g840(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g841(.A(new_n1042), .ZN(new_n1043));
  NOR2_X1   g842(.A1(new_n287), .A2(new_n295), .ZN(new_n1044));
  AOI21_X1  g843(.A(new_n1039), .B1(new_n1043), .B2(new_n1044), .ZN(G1352gat));
  OAI21_X1  g844(.A(G204gat), .B1(new_n1042), .B2(new_n734), .ZN(new_n1046));
  NAND3_X1  g845(.A1(new_n1038), .A2(new_n292), .A3(new_n733), .ZN(new_n1047));
  XOR2_X1   g846(.A(new_n1047), .B(KEYINPUT62), .Z(new_n1048));
  NAND2_X1  g847(.A1(new_n1046), .A2(new_n1048), .ZN(G1353gat));
  NAND3_X1  g848(.A1(new_n1038), .A2(new_n300), .A3(new_n853), .ZN(new_n1050));
  NAND3_X1  g849(.A1(new_n1040), .A2(new_n853), .A3(new_n1041), .ZN(new_n1051));
  AND3_X1   g850(.A1(new_n1051), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1052));
  AOI21_X1  g851(.A(KEYINPUT63), .B1(new_n1051), .B2(G211gat), .ZN(new_n1053));
  OAI21_X1  g852(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(G1354gat));
  OAI21_X1  g853(.A(G218gat), .B1(new_n1042), .B2(new_n766), .ZN(new_n1055));
  NAND3_X1  g854(.A1(new_n1038), .A2(new_n301), .A3(new_n678), .ZN(new_n1056));
  NAND2_X1  g855(.A1(new_n1055), .A2(new_n1056), .ZN(G1355gat));
endmodule


