//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT64), .Z(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT65), .B(G244), .Z(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G116), .A2(G270), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n212), .B1(new_n215), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(G13), .ZN(new_n244));
  NOR3_X1   g0044(.A1(new_n244), .A2(new_n207), .A3(G1), .ZN(new_n245));
  INV_X1    g0045(.A(G68), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT69), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT12), .ZN(new_n248));
  OAI211_X1 g0048(.A(new_n245), .B(new_n246), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n248), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n213), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n245), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n206), .A2(G20), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(G68), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n259), .A2(G77), .B1(G20), .B2(new_n246), .ZN(new_n260));
  INV_X1    g0060(.A(G50), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  AND3_X1   g0064(.A1(new_n264), .A2(KEYINPUT11), .A3(new_n253), .ZN(new_n265));
  AOI21_X1  g0065(.A(KEYINPUT11), .B1(new_n264), .B2(new_n253), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n257), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G232), .A3(G1698), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(G226), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G97), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  OAI211_X1 g0080(.A(G1), .B(G13), .C1(new_n258), .C2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n281), .A2(new_n278), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n279), .B1(G238), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT13), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(KEYINPUT68), .ZN(new_n285));
  AND3_X1   g0085(.A1(new_n276), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n285), .B1(new_n276), .B2(new_n283), .ZN(new_n287));
  OAI21_X1  g0087(.A(G179), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G169), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n276), .A2(new_n283), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT13), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n276), .A2(new_n283), .A3(new_n284), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(KEYINPUT70), .A2(KEYINPUT14), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n288), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n292), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n284), .B1(new_n276), .B2(new_n283), .ZN(new_n297));
  OAI211_X1 g0097(.A(G169), .B(new_n294), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n268), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n261), .B1(new_n206), .B2(G20), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n254), .A2(new_n301), .B1(new_n261), .B2(new_n245), .ZN(new_n302));
  NOR2_X1   g0102(.A1(G50), .A2(G58), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n207), .B1(new_n303), .B2(new_n246), .ZN(new_n304));
  INV_X1    g0104(.A(G150), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n263), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G58), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT8), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT8), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G58), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  AOI211_X1 g0111(.A(new_n304), .B(new_n306), .C1(new_n311), .C2(new_n259), .ZN(new_n312));
  INV_X1    g0112(.A(new_n253), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n302), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n269), .A2(G223), .A3(G1698), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n269), .A2(new_n271), .ZN(new_n316));
  INV_X1    g0116(.A(G222), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n315), .B1(new_n218), .B2(new_n269), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n275), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n279), .B1(G226), .B2(new_n282), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n314), .B1(new_n322), .B2(G169), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n321), .A2(G179), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT9), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n314), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(KEYINPUT9), .B(new_n302), .C1(new_n312), .C2(new_n313), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT10), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n321), .A2(G200), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n319), .A2(G190), .A3(new_n320), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n329), .A2(new_n330), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n327), .A2(new_n332), .A3(new_n328), .ZN(new_n334));
  INV_X1    g0134(.A(new_n331), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT10), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n325), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(G190), .B1(new_n286), .B2(new_n287), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n267), .ZN(new_n339));
  OAI21_X1  g0139(.A(G200), .B1(new_n296), .B2(new_n297), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT67), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT67), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n342), .B(G200), .C1(new_n296), .C2(new_n297), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n339), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n269), .A2(G238), .A3(G1698), .ZN(new_n346));
  INV_X1    g0146(.A(G232), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n346), .B1(new_n203), .B2(new_n269), .C1(new_n316), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n275), .ZN(new_n349));
  INV_X1    g0149(.A(new_n217), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n279), .B1(new_n350), .B2(new_n282), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n289), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n311), .A2(new_n262), .ZN(new_n354));
  INV_X1    g0154(.A(new_n259), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT15), .B(G87), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n354), .B1(new_n207), .B2(new_n218), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n253), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n254), .A2(G77), .A3(new_n255), .ZN(new_n359));
  INV_X1    g0159(.A(new_n245), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n358), .B(new_n359), .C1(G77), .C2(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n353), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n352), .ZN(new_n363));
  INV_X1    g0163(.A(G179), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n361), .B1(G200), .B2(new_n352), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(G190), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n362), .A2(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AND4_X1   g0168(.A1(new_n300), .A2(new_n337), .A3(new_n345), .A4(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT72), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n258), .B2(KEYINPUT3), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT3), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n372), .A2(KEYINPUT72), .A3(G33), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(G20), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n376), .B1(new_n375), .B2(new_n378), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n372), .A2(G33), .ZN(new_n382));
  AOI21_X1  g0182(.A(G20), .B1(new_n382), .B2(new_n374), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT71), .B1(new_n383), .B2(KEYINPUT7), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT71), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n385), .B(new_n377), .C1(new_n269), .C2(G20), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(G68), .B1(new_n381), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n307), .A2(new_n246), .ZN(new_n389));
  NOR2_X1   g0189(.A1(G58), .A2(G68), .ZN(new_n390));
  OAI21_X1  g0190(.A(G20), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n262), .A2(G159), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT16), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n383), .A2(KEYINPUT7), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n377), .B1(new_n269), .B2(G20), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n393), .B1(new_n398), .B2(G68), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n313), .B1(new_n399), .B2(KEYINPUT16), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT74), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT74), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n384), .B(new_n386), .C1(new_n379), .C2(new_n380), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n393), .B1(new_n404), .B2(G68), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n403), .B(new_n400), .C1(new_n405), .C2(KEYINPUT16), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n254), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n311), .A2(new_n255), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n408), .A2(new_n409), .B1(new_n360), .B2(new_n311), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G200), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n282), .A2(G232), .ZN(new_n413));
  INV_X1    g0213(.A(new_n279), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n271), .A2(G226), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n269), .B(new_n416), .C1(G223), .C2(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G87), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n281), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n412), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n419), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n279), .B1(G232), .B2(new_n282), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n420), .B1(new_n423), .B2(G190), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT75), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n424), .B(new_n425), .ZN(new_n426));
  AND4_X1   g0226(.A1(KEYINPUT17), .A2(new_n407), .A3(new_n411), .A4(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n410), .B1(new_n402), .B2(new_n406), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT17), .B1(new_n428), .B2(new_n426), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT16), .ZN(new_n431));
  INV_X1    g0231(.A(new_n380), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n387), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n246), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n431), .B1(new_n436), .B2(new_n393), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n403), .B1(new_n437), .B2(new_n400), .ZN(new_n438));
  INV_X1    g0238(.A(new_n406), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n411), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n423), .A2(new_n364), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(G169), .B2(new_n423), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n440), .A2(KEYINPUT18), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT18), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n428), .B2(new_n442), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n369), .A2(new_n430), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT77), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n382), .A2(new_n374), .A3(G244), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT4), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n451), .A2(new_n452), .B1(G33), .B2(G283), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n269), .A2(KEYINPUT4), .A3(G244), .A4(new_n271), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n452), .B1(new_n269), .B2(G250), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(new_n271), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n450), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n382), .A2(new_n374), .ZN(new_n459));
  INV_X1    g0259(.A(G250), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT4), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G1698), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n462), .A2(KEYINPUT77), .A3(new_n454), .A4(new_n453), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n458), .A2(new_n275), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G190), .ZN(new_n465));
  INV_X1    g0265(.A(G45), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G1), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT5), .B(G41), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n275), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G257), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n275), .A2(new_n277), .ZN(new_n471));
  AND2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n464), .A2(new_n465), .A3(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n453), .B(new_n454), .C1(new_n271), .C2(new_n456), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n281), .B1(new_n480), .B2(new_n450), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n477), .B1(new_n481), .B2(new_n463), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n479), .B1(new_n482), .B2(G200), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n360), .A2(G97), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n258), .A2(G1), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n245), .A2(new_n253), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n486), .B2(G97), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT6), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n488), .A2(new_n202), .A3(G107), .ZN(new_n489));
  XNOR2_X1  g0289(.A(G97), .B(G107), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  OAI22_X1  g0291(.A1(new_n491), .A2(new_n207), .B1(new_n218), .B2(new_n263), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n404), .B2(G107), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n487), .B1(new_n493), .B2(new_n313), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT76), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT76), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n496), .B(new_n487), .C1(new_n493), .C2(new_n313), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n483), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n464), .A2(G179), .A3(new_n478), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n482), .B2(new_n289), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n494), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n382), .A2(new_n374), .A3(G238), .A4(new_n271), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G116), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n502), .B(new_n503), .C1(new_n451), .C2(new_n271), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n275), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n467), .A2(new_n277), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n460), .B1(new_n466), .B2(G1), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(new_n281), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(new_n364), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT78), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n505), .A2(new_n508), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n289), .ZN(new_n513));
  INV_X1    g0313(.A(new_n508), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n504), .B2(new_n275), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(KEYINPUT78), .A3(new_n364), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT19), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n355), .B2(new_n202), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n269), .A2(new_n207), .A3(G68), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n207), .B1(new_n273), .B2(new_n517), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(G87), .B2(new_n204), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n253), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n356), .A2(new_n245), .ZN(new_n524));
  INV_X1    g0324(.A(new_n356), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n486), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n511), .A2(new_n513), .A3(new_n516), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n486), .A2(G87), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n523), .A2(new_n529), .A3(new_n524), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n512), .A2(G200), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n515), .A2(G190), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n498), .A2(new_n501), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT79), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT79), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n498), .A2(new_n537), .A3(new_n501), .A4(new_n534), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n474), .A2(G264), .A3(new_n281), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT82), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n474), .A2(KEYINPUT82), .A3(G264), .A4(new_n281), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n382), .A2(new_n374), .A3(G257), .A4(G1698), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n382), .A2(new_n374), .A3(G250), .A4(new_n271), .ZN(new_n546));
  INV_X1    g0346(.A(G294), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n545), .B(new_n546), .C1(new_n258), .C2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n275), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n544), .A2(new_n476), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n412), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT84), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n544), .A2(new_n476), .A3(new_n549), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n465), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT84), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n550), .A2(new_n555), .A3(new_n412), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n245), .A2(KEYINPUT25), .A3(new_n203), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT81), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT25), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n360), .B2(G107), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(KEYINPUT81), .B(new_n560), .C1(new_n360), .C2(G107), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n486), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n203), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n382), .A2(new_n374), .A3(new_n207), .A4(G87), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT22), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT22), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n269), .A2(new_n569), .A3(new_n207), .A4(G87), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n503), .A2(G20), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT23), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n207), .B2(G107), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT24), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT24), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n571), .A2(new_n579), .A3(new_n576), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n566), .B1(new_n581), .B2(new_n253), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n557), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n253), .ZN(new_n584));
  INV_X1    g0384(.A(new_n566), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n550), .A2(G169), .ZN(new_n587));
  OAI22_X1  g0387(.A1(new_n587), .A2(KEYINPUT83), .B1(new_n364), .B2(new_n550), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n542), .A2(new_n543), .B1(new_n548), .B2(new_n275), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n289), .B1(new_n589), .B2(new_n476), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n586), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n583), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n382), .A2(new_n374), .A3(G257), .A4(new_n271), .ZN(new_n595));
  INV_X1    g0395(.A(G303), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(new_n269), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n269), .A2(G264), .A3(G1698), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n275), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n469), .A2(G270), .B1(new_n471), .B2(new_n475), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n486), .A2(G116), .ZN(new_n602));
  INV_X1    g0402(.A(G116), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n206), .A2(new_n603), .A3(G13), .A4(G20), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n604), .B(KEYINPUT80), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(G20), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n253), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(G20), .B1(G33), .B2(G283), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(G33), .B2(new_n202), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT20), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  AND4_X1   g0410(.A1(KEYINPUT20), .A2(new_n609), .A3(new_n253), .A4(new_n606), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n602), .B(new_n605), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n601), .A2(new_n612), .A3(G169), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n599), .A2(new_n600), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n616), .A2(G179), .A3(new_n612), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n601), .A2(new_n612), .A3(KEYINPUT21), .A4(G169), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(G190), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n612), .B1(new_n601), .B2(G200), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n449), .A2(new_n539), .A3(new_n594), .A4(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n619), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n593), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n513), .A2(new_n509), .A3(new_n527), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n533), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n557), .B2(new_n582), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n625), .A2(new_n501), .A3(new_n498), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n495), .A2(new_n497), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  INV_X1    g0431(.A(new_n627), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n630), .A2(new_n631), .A3(new_n500), .A4(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n626), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n534), .A2(new_n494), .A3(new_n500), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n634), .B1(new_n635), .B2(KEYINPUT26), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n629), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n449), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n407), .A2(new_n426), .A3(new_n411), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT17), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n362), .A2(new_n365), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n300), .B1(new_n344), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n428), .A2(KEYINPUT17), .A3(new_n426), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n447), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n333), .A2(new_n336), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n325), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n638), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g0449(.A(new_n649), .B(KEYINPUT85), .Z(G369));
  NAND3_X1  g0450(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G343), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n612), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n622), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT86), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n624), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n659), .B2(new_n660), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT87), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n663), .A2(G330), .ZN(new_n664));
  INV_X1    g0464(.A(new_n656), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n594), .B1(new_n582), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n593), .B2(new_n665), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n619), .A2(new_n665), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n594), .A2(new_n670), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n590), .A2(new_n591), .B1(new_n553), .B2(G179), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n587), .A2(KEYINPUT83), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n582), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n671), .B1(new_n674), .B2(new_n665), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n668), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n210), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n216), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n464), .A2(new_n478), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n601), .A2(new_n364), .A3(new_n512), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(new_n550), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n515), .A2(new_n544), .A3(new_n549), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n599), .A2(new_n600), .A3(G179), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n482), .A2(new_n689), .A3(KEYINPUT30), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT30), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n616), .A2(G179), .A3(new_n515), .A4(new_n589), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n692), .B1(new_n684), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT88), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT30), .B1(new_n482), .B2(new_n689), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT89), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n690), .B(new_n686), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n694), .A2(KEYINPUT89), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n656), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT31), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT88), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n695), .A2(new_n705), .A3(KEYINPUT31), .A4(new_n656), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n697), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n622), .A2(new_n593), .A3(new_n583), .A4(new_n665), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n536), .B2(new_n538), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G330), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n637), .A2(new_n713), .A3(new_n665), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n534), .A2(new_n500), .A3(new_n631), .A4(new_n494), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n626), .B(KEYINPUT90), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n630), .A2(new_n500), .A3(new_n632), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT26), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n498), .A2(new_n501), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT91), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n674), .B2(new_n619), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n593), .A2(new_n624), .A3(KEYINPUT91), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n721), .A2(new_n628), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n656), .B1(new_n720), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n714), .B1(new_n726), .B2(new_n713), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n712), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n683), .B1(new_n728), .B2(G1), .ZN(G364));
  NOR2_X1   g0529(.A1(new_n244), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n206), .B1(new_n730), .B2(G45), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n678), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n664), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(G330), .B2(new_n663), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n677), .A2(new_n459), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G355), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(G116), .B2(new_n210), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n677), .A2(new_n269), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n216), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n740), .B1(new_n466), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n242), .A2(G45), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n738), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n213), .B1(G20), .B2(new_n289), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n733), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n207), .A2(G179), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(new_n465), .A3(new_n412), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G159), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT94), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT32), .Z(new_n757));
  NOR2_X1   g0557(.A1(new_n207), .A2(new_n364), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n465), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT92), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n760), .A2(KEYINPUT92), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n752), .A2(G190), .A3(G200), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT95), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G58), .A2(new_n765), .B1(new_n771), .B2(G87), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n759), .A2(new_n364), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n758), .A2(new_n465), .A3(G200), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n775), .A2(new_n202), .B1(new_n776), .B2(new_n246), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n752), .A2(new_n465), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n203), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n758), .A2(new_n465), .A3(new_n412), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n269), .B1(new_n780), .B2(new_n218), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n777), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n758), .A2(G190), .A3(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(KEYINPUT93), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n783), .A2(KEYINPUT93), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n772), .B(new_n782), .C1(new_n261), .C2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G322), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n764), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n770), .A2(new_n596), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n459), .B1(new_n780), .B2(new_n792), .C1(new_n775), .C2(new_n547), .ZN(new_n793));
  OR3_X1    g0593(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n776), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT33), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(G317), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(G317), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n795), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n778), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n800), .A2(G283), .B1(new_n754), .B2(G329), .ZN(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT96), .B(G326), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n799), .B(new_n801), .C1(new_n787), .C2(new_n802), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n757), .A2(new_n788), .B1(new_n794), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n751), .B1(new_n804), .B2(new_n748), .ZN(new_n805));
  INV_X1    g0605(.A(new_n747), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n663), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n735), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  NOR2_X1   g0609(.A1(new_n748), .A2(new_n745), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT97), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n733), .B1(new_n811), .B2(G77), .ZN(new_n812));
  INV_X1    g0612(.A(new_n780), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G150), .A2(new_n795), .B1(new_n813), .B2(G159), .ZN(new_n814));
  INV_X1    g0614(.A(G143), .ZN(new_n815));
  INV_X1    g0615(.A(G137), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n814), .B1(new_n764), .B2(new_n815), .C1(new_n816), .C2(new_n787), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT34), .Z(new_n818));
  INV_X1    g0618(.A(G132), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n775), .A2(new_n307), .B1(new_n753), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n269), .B1(new_n778), .B2(new_n246), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n261), .B2(new_n770), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n459), .B1(new_n770), .B2(new_n203), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT98), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n775), .A2(new_n202), .B1(new_n780), .B2(new_n603), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n800), .A2(G87), .ZN(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n828), .B2(new_n776), .C1(new_n792), .C2(new_n753), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n826), .B(new_n829), .C1(G294), .C2(new_n765), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n596), .B2(new_n787), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n818), .A2(new_n823), .B1(new_n825), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n812), .B1(new_n832), .B2(new_n748), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n361), .A2(new_n656), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n368), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT99), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT99), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n368), .A2(new_n837), .A3(new_n834), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n836), .B(new_n838), .C1(new_n642), .C2(new_n665), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n833), .B1(new_n839), .B2(new_n746), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(new_n637), .B2(new_n665), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n836), .A2(new_n838), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n637), .A2(new_n842), .A3(new_n665), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n733), .B1(new_n712), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n712), .A2(new_n845), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT100), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n712), .A2(new_n845), .A3(KEYINPUT100), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n840), .B1(new_n849), .B2(new_n850), .ZN(G384));
  INV_X1    g0651(.A(new_n491), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n852), .A2(KEYINPUT35), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(KEYINPUT35), .ZN(new_n854));
  NOR4_X1   g0654(.A1(new_n853), .A2(new_n854), .A3(new_n603), .A4(new_n215), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT36), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n741), .B(G77), .C1(new_n307), .C2(new_n246), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n261), .A2(G68), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n206), .B(G13), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n642), .A2(new_n656), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n843), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n345), .A2(new_n300), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n267), .A2(new_n665), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n295), .A2(new_n299), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n865), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n400), .B1(KEYINPUT16), .B2(new_n399), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n874), .A2(new_n411), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n654), .B(new_n875), .C1(new_n430), .C2(new_n447), .ZN(new_n876));
  INV_X1    g0676(.A(new_n654), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n443), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n878), .A2(new_n875), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n407), .A2(new_n411), .A3(new_n426), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT37), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n440), .B1(new_n443), .B2(new_n877), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT37), .B1(new_n428), .B2(new_n426), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n873), .B1(new_n876), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n875), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n444), .A2(new_n446), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n641), .A2(new_n644), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n877), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n872), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n889), .B2(new_n654), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT39), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n891), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n440), .B(new_n877), .C1(new_n889), .C2(new_n890), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT101), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(new_n880), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n639), .B(KEYINPUT101), .C1(new_n428), .C2(new_n878), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n884), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n895), .B1(new_n896), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n887), .A2(KEYINPUT39), .A3(new_n892), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n300), .A2(new_n656), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n894), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n646), .A2(new_n647), .ZN(new_n910));
  INV_X1    g0710(.A(new_n325), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n727), .B2(new_n449), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n909), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n839), .B1(new_n869), .B2(new_n866), .ZN(new_n915));
  INV_X1    g0715(.A(new_n708), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n539), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n702), .A2(new_n703), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n694), .A2(KEYINPUT89), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n698), .A2(new_n699), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n691), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT31), .B1(new_n921), .B2(new_n656), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n917), .A2(new_n923), .A3(KEYINPUT102), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT102), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n921), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n704), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n925), .B1(new_n709), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n915), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n896), .B2(new_n904), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT40), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT40), .B1(new_n887), .B2(new_n892), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n929), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n448), .B1(new_n924), .B2(new_n928), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n711), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n935), .B2(new_n934), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n914), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n730), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n938), .B1(G1), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT103), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n914), .A2(new_n937), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n940), .B2(new_n941), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n860), .B1(new_n943), .B2(new_n945), .ZN(G367));
  NAND2_X1  g0746(.A1(new_n630), .A2(new_n656), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n721), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n630), .A2(new_n500), .A3(new_n656), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n671), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT42), .Z(new_n952));
  INV_X1    g0752(.A(new_n950), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n501), .B1(new_n953), .B2(new_n593), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n665), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n530), .A2(new_n665), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n626), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n632), .B2(new_n957), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT104), .Z(new_n960));
  INV_X1    g0760(.A(KEYINPUT43), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n956), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT105), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n960), .A2(new_n961), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n956), .A2(new_n965), .A3(new_n962), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n668), .A2(new_n953), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n678), .B(KEYINPUT41), .Z(new_n970));
  NAND2_X1  g0770(.A1(new_n675), .A2(new_n950), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT106), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT45), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT106), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n971), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT45), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n675), .A2(new_n950), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT44), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n974), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n668), .ZN(new_n981));
  INV_X1    g0781(.A(new_n671), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n667), .B2(new_n670), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n664), .B(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n728), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n970), .B1(new_n985), .B2(new_n728), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n969), .B1(new_n986), .B2(new_n732), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n960), .A2(new_n747), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n750), .B1(new_n677), .B2(new_n525), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n739), .A2(new_n234), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n678), .B(new_n732), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n459), .B1(new_n778), .B2(new_n202), .C1(new_n828), .C2(new_n780), .ZN(new_n992));
  XNOR2_X1  g0792(.A(KEYINPUT107), .B(G317), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n754), .A2(new_n993), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n547), .B2(new_n776), .C1(new_n775), .C2(new_n203), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n992), .B(new_n995), .C1(G303), .C2(new_n765), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n771), .A2(G116), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT46), .ZN(new_n998));
  INV_X1    g0798(.A(new_n787), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n997), .A2(new_n998), .B1(new_n999), .B2(G311), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n996), .B(new_n1000), .C1(new_n998), .C2(new_n997), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT108), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n778), .A2(new_n218), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(new_n459), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT109), .Z(new_n1005));
  AOI22_X1  g0805(.A1(G150), .A2(new_n765), .B1(new_n771), .B2(G58), .ZN(new_n1006));
  INV_X1    g0806(.A(G159), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n775), .A2(new_n246), .B1(new_n776), .B2(new_n1007), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n780), .A2(new_n261), .B1(new_n753), .B2(new_n816), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n999), .A2(G143), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1005), .A2(new_n1006), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1002), .A2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT110), .Z(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT47), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n748), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n988), .B(new_n991), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT111), .Z(new_n1018));
  NAND2_X1  g0818(.A1(new_n987), .A2(new_n1018), .ZN(G387));
  AOI21_X1  g0819(.A(new_n679), .B1(new_n984), .B2(new_n728), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n728), .B2(new_n984), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n667), .A2(new_n806), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n311), .A2(new_n261), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT50), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n680), .B(new_n466), .C1(new_n246), .C2(new_n218), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n739), .B1(new_n1024), .B2(new_n1025), .C1(new_n231), .C2(new_n466), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n680), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n736), .A2(new_n1027), .B1(new_n203), .B2(new_n677), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(KEYINPUT112), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n749), .ZN(new_n1030));
  AOI21_X1  g0830(.A(KEYINPUT112), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n733), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n459), .B1(new_n813), .B2(G68), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n202), .B2(new_n778), .C1(new_n770), .C2(new_n218), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n311), .A2(new_n795), .B1(new_n774), .B2(new_n525), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n305), .B2(new_n753), .C1(new_n787), .C2(new_n1007), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1034), .B(new_n1036), .C1(G50), .C2(new_n765), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT113), .Z(new_n1038));
  OAI22_X1  g0838(.A1(new_n770), .A2(new_n547), .B1(new_n828), .B2(new_n775), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT114), .Z(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n765), .A2(new_n993), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G303), .A2(new_n813), .B1(new_n795), .B2(G311), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(new_n787), .C2(new_n789), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1040), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT49), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n459), .B1(new_n753), .B2(new_n802), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G116), .B2(new_n800), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1038), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1032), .B1(new_n1052), .B2(new_n748), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n984), .A2(new_n732), .B1(new_n1022), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1021), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT115), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1021), .A2(KEYINPUT115), .A3(new_n1054), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(G393));
  INV_X1    g0859(.A(new_n668), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n980), .B(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n984), .A2(new_n728), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n985), .A2(new_n678), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n981), .A2(new_n732), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n239), .A2(new_n740), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n749), .B1(new_n202), .B2(new_n210), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n733), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n999), .A2(G317), .B1(new_n765), .B2(G311), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT52), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n269), .B(new_n779), .C1(G294), .C2(new_n813), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n828), .B2(new_n770), .C1(new_n789), .C2(new_n753), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G303), .A2(new_n795), .B1(new_n774), .B2(G116), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT116), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n1070), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n787), .A2(new_n305), .B1(new_n764), .B2(new_n1007), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT51), .Z(new_n1077));
  NAND2_X1  g0877(.A1(new_n774), .A2(G77), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(new_n815), .B2(new_n753), .C1(new_n261), .C2(new_n776), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n459), .B1(new_n813), .B2(new_n311), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n827), .B(new_n1080), .C1(new_n770), .C2(new_n246), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1077), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1075), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1068), .B1(new_n1083), .B2(new_n748), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n950), .B2(new_n806), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1064), .A2(new_n1065), .A3(new_n1085), .ZN(G390));
  AOI21_X1  g0886(.A(new_n907), .B1(new_n863), .B2(new_n871), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(KEYINPUT38), .B1(new_n891), .B2(new_n885), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n896), .A2(new_n1089), .A3(new_n895), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n428), .B(new_n654), .C1(new_n430), .C2(new_n447), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n900), .A2(new_n901), .B1(new_n883), .B2(new_n882), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n873), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT39), .B1(new_n1093), .B2(new_n892), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1088), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(G330), .B(new_n839), .C1(new_n707), .C2(new_n709), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1096), .A2(new_n870), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1093), .A2(new_n892), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n723), .A2(new_n724), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n628), .A2(new_n498), .A3(new_n501), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n719), .B(new_n717), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n665), .A3(new_n842), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n862), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n907), .B1(new_n1103), .B2(new_n871), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1098), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1095), .A2(new_n1097), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n924), .A2(new_n928), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1107), .A2(G330), .A3(new_n839), .A4(new_n871), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1087), .B1(new_n905), .B2(new_n906), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1098), .A2(new_n1104), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1106), .A2(new_n1112), .A3(new_n732), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n745), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n733), .B1(new_n811), .B2(new_n311), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1078), .B1(new_n547), .B2(new_n753), .C1(new_n203), .C2(new_n776), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G283), .B2(new_n999), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n459), .B1(new_n778), .B2(new_n246), .C1(new_n202), .C2(new_n780), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n771), .B2(G87), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1117), .B(new_n1119), .C1(new_n603), .C2(new_n764), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n771), .A2(G150), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1121), .A2(KEYINPUT53), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1121), .A2(KEYINPUT53), .B1(new_n999), .B2(G128), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n765), .A2(G132), .ZN(new_n1124));
  XOR2_X1   g0924(.A(KEYINPUT54), .B(G143), .Z(new_n1125));
  NAND2_X1  g0925(.A1(new_n813), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1007), .B2(new_n775), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(G137), .B2(new_n795), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .A4(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(G125), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n269), .B1(new_n778), .B2(new_n261), .C1(new_n1130), .C2(new_n753), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT118), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1120), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1115), .B1(new_n1133), .B2(new_n748), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1114), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1113), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT119), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT119), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1113), .A2(new_n1138), .A3(new_n1135), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1106), .A2(new_n1112), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1107), .A2(G330), .A3(new_n449), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT117), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n913), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n711), .B(new_n448), .C1(new_n924), .C2(new_n928), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n713), .B1(new_n1101), .B2(new_n665), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n637), .A2(new_n713), .A3(new_n665), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n449), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n648), .ZN(new_n1149));
  OAI21_X1  g0949(.A(KEYINPUT117), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1096), .A2(new_n870), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1108), .A2(new_n1151), .B1(new_n843), .B2(new_n862), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n862), .B(new_n1102), .C1(new_n1096), .C2(new_n870), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1107), .A2(G330), .A3(new_n839), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1153), .B1(new_n1154), .B2(new_n870), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1144), .B(new_n1150), .C1(new_n1152), .C2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n679), .B1(new_n1141), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1156), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(new_n1106), .A3(new_n1112), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1140), .A2(new_n1160), .ZN(G378));
  INV_X1    g0961(.A(KEYINPUT123), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1150), .A2(new_n1162), .A3(new_n1144), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1162), .B1(new_n1150), .B2(new_n1144), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n1141), .B2(new_n1156), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n314), .A2(new_n877), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n337), .B(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(KEYINPUT40), .A2(new_n930), .B1(new_n932), .B2(new_n929), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n1171), .B2(new_n711), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1170), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n934), .A2(G330), .A3(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1172), .A2(new_n1174), .A3(new_n909), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n909), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1166), .B(KEYINPUT57), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n678), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n909), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1172), .A2(new_n1174), .A3(new_n909), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT57), .B1(new_n1183), .B2(new_n1166), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1178), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n732), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n732), .B(new_n678), .C1(new_n261), .C2(new_n810), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n776), .A2(new_n819), .B1(new_n780), .B2(new_n816), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n765), .A2(G128), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n771), .A2(new_n1125), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1188), .B(new_n1189), .C1(KEYINPUT121), .C2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(KEYINPUT121), .B2(new_n1190), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n787), .A2(new_n1130), .B1(new_n305), .B2(new_n775), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT122), .Z(new_n1194));
  NOR2_X1   g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n800), .A2(G159), .ZN(new_n1199));
  AOI211_X1 g0999(.A(G33), .B(G41), .C1(new_n754), .C2(G124), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n269), .A2(G41), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n356), .B2(new_n780), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G68), .B2(new_n774), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n218), .B2(new_n770), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n778), .A2(new_n307), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G97), .B2(new_n795), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n828), .B2(new_n753), .C1(new_n787), .C2(new_n603), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1205), .B(new_n1208), .C1(G107), .C2(new_n765), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT120), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(KEYINPUT58), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1210), .A2(KEYINPUT58), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1202), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1213), .B(new_n261), .C1(G33), .C2(G41), .ZN(new_n1214));
  AND4_X1   g1014(.A1(new_n1201), .A2(new_n1211), .A3(new_n1212), .A4(new_n1214), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1187), .B1(new_n1173), .B2(new_n746), .C1(new_n1016), .C2(new_n1215), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1186), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1185), .A2(new_n1217), .ZN(G375));
  OAI21_X1  g1018(.A(new_n732), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT124), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n870), .A2(new_n745), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n733), .B1(new_n811), .B2(G68), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n269), .B(new_n1003), .C1(G107), .C2(new_n813), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n202), .B2(new_n770), .C1(new_n828), .C2(new_n764), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G116), .A2(new_n795), .B1(new_n774), .B2(new_n525), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n596), .B2(new_n753), .C1(new_n787), .C2(new_n547), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n459), .B(new_n1206), .C1(G150), .C2(new_n813), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1228), .B1(new_n816), .B2(new_n764), .C1(new_n1007), .C2(new_n770), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n754), .A2(G128), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n795), .A2(new_n1125), .B1(new_n774), .B2(G50), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n787), .C2(new_n819), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1225), .A2(new_n1227), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1223), .B1(new_n1233), .B2(new_n748), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1219), .A2(new_n1220), .B1(new_n1222), .B2(new_n1234), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1221), .A2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1150), .A2(new_n1144), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n970), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1240), .A3(new_n1156), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1236), .A2(new_n1241), .ZN(G381));
  INV_X1    g1042(.A(G375), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1137), .A2(new_n1139), .B1(new_n1159), .B2(new_n1157), .ZN(new_n1244));
  INV_X1    g1044(.A(G390), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(new_n987), .A3(new_n1018), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NOR4_X1   g1047(.A1(G393), .A2(G396), .A3(G384), .A4(G381), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1243), .A2(new_n1244), .A3(new_n1247), .A4(new_n1248), .ZN(G407));
  NAND2_X1  g1049(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G407), .B(G213), .C1(G343), .C2(new_n1250), .ZN(G409));
  NAND2_X1  g1051(.A1(G387), .A2(G390), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1246), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(G393), .A2(G396), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n808), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1252), .B(new_n1246), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1166), .B(new_n1240), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n1186), .A3(new_n1216), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1244), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT125), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1217), .B(G378), .C1(new_n1178), .C2(new_n1184), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1261), .A2(KEYINPUT125), .A3(new_n1244), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n655), .A2(G213), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1239), .B(KEYINPUT60), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1269), .A2(new_n678), .A3(new_n1156), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1270), .A2(new_n1236), .A3(G384), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G384), .B1(new_n1270), .B2(new_n1236), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1267), .A2(new_n1268), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT126), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT62), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1267), .A2(new_n1273), .A3(new_n1277), .A4(new_n1268), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1275), .A2(new_n1276), .A3(new_n1278), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n655), .A2(G213), .A3(G2897), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1273), .B(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT127), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1267), .A2(new_n1282), .A3(new_n1268), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1282), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1281), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1279), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1276), .B1(new_n1288), .B2(new_n1273), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1259), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1257), .A2(new_n1286), .A3(new_n1258), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1291), .B1(new_n1292), .B2(new_n1281), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1288), .A2(KEYINPUT63), .A3(new_n1273), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1293), .B(new_n1294), .C1(KEYINPUT63), .C2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1290), .A2(new_n1296), .ZN(G405));
  NAND2_X1  g1097(.A1(G375), .A2(new_n1244), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1259), .A2(new_n1265), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1265), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1257), .A2(new_n1300), .A3(new_n1258), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1273), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1302), .B(new_n1303), .ZN(G402));
endmodule


