//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT2), .B(G113), .Z(new_n188));
  XNOR2_X1  g002(.A(G116), .B(G119), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT70), .ZN(new_n191));
  OR2_X1    g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n191), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(new_n194), .B2(G107), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT79), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G104), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(new_n197), .A3(G104), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(KEYINPUT79), .A3(G107), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n195), .A2(new_n198), .A3(new_n200), .A4(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT4), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G101), .ZN(new_n204));
  OR2_X1    g018(.A1(new_n202), .A2(G101), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(G101), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n192), .A2(new_n193), .A3(new_n204), .A4(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n194), .A3(G107), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n194), .B2(G107), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n209), .B1(new_n194), .B2(G107), .ZN(new_n212));
  OAI21_X1  g026(.A(G101), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n205), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n188), .A2(new_n189), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n189), .A2(KEYINPUT5), .ZN(new_n216));
  INV_X1    g030(.A(G119), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G116), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n216), .B(G113), .C1(KEYINPUT5), .C2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n214), .A2(new_n215), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n208), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g035(.A(G110), .B(G122), .Z(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n222), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n208), .A2(new_n220), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(KEYINPUT6), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n227));
  INV_X1    g041(.A(G143), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(G146), .ZN(new_n229));
  INV_X1    g043(.A(G146), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(KEYINPUT64), .A3(G143), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n229), .A2(new_n231), .B1(new_n228), .B2(G146), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT0), .A3(G128), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n228), .A2(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(G143), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n234), .A2(new_n235), .B1(KEYINPUT0), .B2(G128), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(KEYINPUT0), .B2(G128), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G125), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G128), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n234), .A2(new_n235), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n229), .A2(new_n231), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n245), .A3(G128), .A4(new_n234), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G125), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n239), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G224), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n250), .A2(G224), .A3(new_n252), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT6), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n221), .A2(new_n257), .A3(new_n222), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n226), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G902), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT81), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n214), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n219), .A2(new_n215), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XOR2_X1   g078(.A(new_n222), .B(KEYINPUT8), .Z(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT7), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n253), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n254), .A2(new_n255), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n251), .A2(new_n267), .A3(new_n253), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n266), .A2(new_n269), .A3(new_n225), .A4(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n259), .A2(new_n260), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G210), .B1(G237), .B2(G902), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n272), .A2(KEYINPUT82), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(KEYINPUT82), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n259), .A2(new_n271), .A3(new_n260), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(G214), .B1(G237), .B2(G902), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n187), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n279), .ZN(new_n281));
  AOI211_X1 g095(.A(KEYINPUT83), .B(new_n281), .C1(new_n275), .C2(new_n277), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT86), .ZN(new_n284));
  INV_X1    g098(.A(G237), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(new_n252), .A3(G214), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n228), .ZN(new_n287));
  NOR2_X1   g101(.A1(G237), .A2(G953), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(G143), .A3(G214), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n284), .B1(new_n290), .B2(G131), .ZN(new_n291));
  INV_X1    g105(.A(G131), .ZN(new_n292));
  AOI211_X1 g106(.A(KEYINPUT86), .B(new_n292), .C1(new_n287), .C2(new_n289), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT17), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n248), .A2(KEYINPUT16), .A3(G140), .ZN(new_n295));
  XNOR2_X1  g109(.A(G125), .B(G140), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(KEYINPUT16), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(new_n230), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n286), .A2(new_n228), .ZN(new_n299));
  AOI21_X1  g113(.A(G143), .B1(new_n288), .B2(G214), .ZN(new_n300));
  OAI21_X1  g114(.A(G131), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT86), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n290), .A2(new_n284), .A3(G131), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n287), .A2(new_n292), .A3(new_n289), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT85), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n287), .A2(KEYINPUT85), .A3(new_n292), .A4(new_n289), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n302), .A2(new_n303), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n294), .B(new_n298), .C1(new_n308), .C2(KEYINPUT17), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n296), .A2(new_n230), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT75), .ZN(new_n311));
  OR2_X1    g125(.A1(new_n296), .A2(new_n230), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(KEYINPUT18), .A2(G131), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n290), .B(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(G113), .B(G122), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(new_n194), .ZN(new_n318));
  XOR2_X1   g132(.A(new_n318), .B(KEYINPUT88), .Z(new_n319));
  NAND3_X1  g133(.A1(new_n309), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n309), .A2(new_n316), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n318), .B1(new_n322), .B2(KEYINPUT89), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT89), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n309), .A2(new_n324), .A3(new_n316), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n321), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G475), .B1(new_n326), .B2(G902), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n297), .A2(G146), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n296), .A2(KEYINPUT87), .A3(KEYINPUT19), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT19), .B1(new_n296), .B2(KEYINPUT87), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n230), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n308), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n316), .ZN(new_n334));
  INV_X1    g148(.A(new_n318), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n320), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT20), .ZN(new_n338));
  INV_X1    g152(.A(G475), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n337), .A2(new_n338), .A3(new_n339), .A4(new_n260), .ZN(new_n340));
  AOI211_X1 g154(.A(G475), .B(G902), .C1(new_n336), .C2(new_n320), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n342));
  OAI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n327), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n252), .A2(G952), .ZN(new_n346));
  NAND2_X1  g160(.A1(G234), .A2(G237), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XOR2_X1   g162(.A(KEYINPUT21), .B(G898), .Z(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(G902), .A3(G953), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G116), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G122), .ZN(new_n353));
  INV_X1    g167(.A(G122), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G116), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n355), .A3(new_n197), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n197), .B1(new_n353), .B2(new_n355), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT90), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n353), .A2(new_n355), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G107), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT90), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n356), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n228), .A2(G128), .ZN(new_n364));
  INV_X1    g178(.A(G128), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G143), .ZN(new_n366));
  INV_X1    g180(.A(G134), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n364), .A2(new_n366), .A3(KEYINPUT13), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n369), .B(G134), .C1(KEYINPUT13), .C2(new_n364), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n359), .A2(new_n363), .A3(new_n368), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n364), .A2(new_n366), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G134), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n357), .B1(new_n373), .B2(new_n368), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT14), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n354), .A2(G116), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n375), .A2(new_n376), .B1(new_n355), .B2(KEYINPUT91), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n375), .A2(new_n352), .A3(KEYINPUT91), .A4(G122), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n378), .B1(new_n375), .B2(new_n376), .ZN(new_n379));
  OAI21_X1  g193(.A(G107), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n374), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n371), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT9), .B(G234), .ZN(new_n383));
  INV_X1    g197(.A(G217), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n383), .A2(new_n384), .A3(G953), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT92), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n371), .A2(new_n381), .A3(new_n385), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n382), .A2(KEYINPUT92), .A3(new_n386), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n390), .A2(KEYINPUT93), .A3(new_n260), .A4(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G478), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(KEYINPUT15), .ZN(new_n394));
  XOR2_X1   g208(.A(new_n392), .B(new_n394), .Z(new_n395));
  NAND3_X1  g209(.A1(new_n345), .A2(new_n351), .A3(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n283), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT32), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT31), .ZN(new_n399));
  OAI211_X1 g213(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n367), .C2(G137), .ZN(new_n400));
  NAND2_X1  g214(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n401));
  INV_X1    g215(.A(G137), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(G134), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  OR3_X1    g218(.A1(new_n402), .A2(KEYINPUT66), .A3(G134), .ZN(new_n405));
  NOR2_X1   g219(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n367), .A2(G137), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n406), .B1(new_n407), .B2(KEYINPUT66), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n404), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT67), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT67), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n404), .A2(new_n408), .A3(new_n411), .A4(new_n405), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(G131), .A3(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n404), .A2(new_n408), .A3(new_n292), .A4(new_n405), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n414), .A2(KEYINPUT68), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT68), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n410), .A2(new_n417), .A3(G131), .A4(new_n412), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n238), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n407), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n367), .A2(G137), .ZN(new_n421));
  OAI21_X1  g235(.A(G131), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n247), .A2(new_n414), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT69), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT69), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n247), .A2(new_n425), .A3(new_n414), .A4(new_n422), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n419), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT30), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n192), .A2(new_n193), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n419), .A2(KEYINPUT30), .A3(new_n423), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n419), .A2(new_n431), .A3(new_n423), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(G101), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n288), .A2(G210), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n434), .A2(new_n435), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT71), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT71), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n434), .A2(new_n442), .A3(new_n435), .A4(new_n439), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n399), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n435), .A2(KEYINPUT28), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n435), .A2(KEYINPUT28), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n428), .A2(new_n432), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n439), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n440), .A2(new_n451), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n444), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(G472), .A2(G902), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n398), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n441), .A2(new_n443), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT31), .ZN(new_n458));
  INV_X1    g272(.A(new_n449), .ZN(new_n459));
  INV_X1    g273(.A(new_n452), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(KEYINPUT32), .A3(new_n454), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n434), .A2(new_n435), .ZN(new_n463));
  INV_X1    g277(.A(new_n439), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT73), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n447), .A2(new_n448), .A3(new_n439), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n463), .A2(KEYINPUT73), .A3(new_n464), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT29), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n467), .A2(new_n468), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n431), .B1(new_n419), .B2(new_n423), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(new_n445), .B2(new_n446), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n464), .A2(new_n470), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G472), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n456), .A2(new_n462), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n365), .A2(G119), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT74), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n217), .A2(G128), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g297(.A(KEYINPUT24), .B(G110), .Z(new_n484));
  AND2_X1   g298(.A1(new_n479), .A2(KEYINPUT23), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n479), .A2(KEYINPUT23), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI22_X1  g301(.A1(new_n483), .A2(new_n484), .B1(G110), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n328), .A3(new_n311), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT76), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n298), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n483), .A2(new_n484), .B1(G110), .B2(new_n487), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n489), .A2(new_n490), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n491), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n252), .A2(G221), .A3(G234), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT22), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(new_n402), .ZN(new_n499));
  OR2_X1    g313(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n499), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n500), .A2(new_n260), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n503));
  OR2_X1    g317(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n384), .B1(G234), .B2(new_n260), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n505), .B(new_n506), .C1(new_n503), .C2(new_n502), .ZN(new_n507));
  INV_X1    g321(.A(new_n506), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT78), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n509), .A2(KEYINPUT78), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n507), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(G221), .B1(new_n383), .B2(G902), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G469), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(new_n260), .ZN(new_n516));
  INV_X1    g330(.A(new_n241), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n246), .B1(new_n517), .B2(new_n232), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n214), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n519), .B1(new_n247), .B2(new_n214), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n416), .A2(new_n418), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT12), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT12), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(G110), .B(G140), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n252), .A2(G227), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT10), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n519), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n207), .A2(new_n238), .A3(new_n204), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n214), .A2(KEYINPUT10), .A3(new_n247), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n416), .A2(new_n418), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n530), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n526), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(new_n521), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n534), .A2(new_n533), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n536), .B1(new_n541), .B2(new_n532), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n530), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(G902), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n516), .B1(new_n544), .B2(new_n515), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n539), .A2(new_n521), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n537), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n540), .B1(new_n525), .B2(new_n524), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n547), .B(G469), .C1(new_n548), .C2(new_n529), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n514), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n397), .A2(new_n478), .A3(new_n512), .A4(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(G101), .ZN(G3));
  INV_X1    g366(.A(G472), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n461), .B2(new_n260), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n453), .A2(new_n455), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n512), .A3(new_n550), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT33), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n390), .A2(new_n558), .A3(new_n391), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n387), .A2(KEYINPUT33), .A3(new_n389), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT94), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n561), .A2(new_n562), .A3(G478), .A4(new_n260), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n390), .A2(new_n260), .A3(new_n391), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n393), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n559), .A2(G478), .A3(new_n260), .A4(new_n560), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT94), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n344), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n272), .A2(new_n273), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n259), .A2(new_n271), .A3(new_n260), .A4(new_n274), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n570), .A2(new_n279), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n351), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n557), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT34), .B(G104), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(G6));
  XNOR2_X1  g390(.A(new_n341), .B(new_n342), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n577), .A2(KEYINPUT95), .ZN(new_n578));
  INV_X1    g392(.A(new_n395), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(KEYINPUT95), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n578), .A2(new_n579), .A3(new_n327), .A4(new_n580), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n557), .A2(new_n573), .A3(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G107), .Z(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT96), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n582), .B(new_n584), .ZN(G9));
  NOR2_X1   g399(.A1(new_n499), .A2(KEYINPUT36), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n496), .B(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n506), .A2(G902), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT97), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n587), .A2(KEYINPUT97), .A3(new_n588), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n507), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n397), .A2(new_n556), .A3(new_n550), .A4(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT99), .B(G110), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT98), .B(KEYINPUT37), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G12));
  NAND2_X1  g414(.A1(new_n545), .A2(new_n549), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n513), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n570), .A2(new_n279), .A3(new_n571), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n348), .B1(G900), .B2(new_n350), .ZN(new_n605));
  XOR2_X1   g419(.A(new_n605), .B(KEYINPUT100), .Z(new_n606));
  NOR2_X1   g420(.A1(new_n581), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n478), .A2(new_n595), .A3(new_n604), .A4(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G128), .ZN(G30));
  INV_X1    g423(.A(new_n472), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n439), .B1(new_n610), .B2(new_n435), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n441), .B2(new_n443), .ZN(new_n612));
  OAI21_X1  g426(.A(G472), .B1(new_n612), .B2(G902), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n456), .A2(new_n462), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT101), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n456), .A2(new_n462), .A3(new_n616), .A4(new_n613), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n606), .B(KEYINPUT39), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n602), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT40), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n619), .A2(new_n595), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n344), .A2(new_n579), .ZN(new_n625));
  AOI211_X1 g439(.A(new_n281), .B(new_n625), .C1(new_n621), .C2(new_n622), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n278), .B(KEYINPUT38), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G143), .ZN(G45));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n630));
  INV_X1    g444(.A(new_n606), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n568), .A2(new_n344), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n568), .A2(new_n344), .A3(new_n631), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT102), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n550), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n478), .A2(new_n572), .A3(new_n595), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G146), .ZN(G48));
  NOR2_X1   g451(.A1(new_n573), .A2(new_n569), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n535), .A2(new_n536), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n546), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n640), .A2(new_n530), .B1(new_n526), .B2(new_n537), .ZN(new_n641));
  OAI21_X1  g455(.A(G469), .B1(new_n641), .B2(G902), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n538), .A2(new_n543), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n643), .A2(new_n515), .A3(new_n260), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n642), .A2(new_n513), .A3(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n478), .A2(new_n512), .A3(new_n638), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT41), .B(G113), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G15));
  NOR2_X1   g462(.A1(new_n581), .A2(new_n573), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n478), .A2(new_n512), .A3(new_n649), .A4(new_n645), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G116), .ZN(G18));
  INV_X1    g465(.A(new_n396), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n645), .A2(KEYINPUT103), .A3(new_n572), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n642), .A2(new_n513), .A3(new_n644), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n654), .B1(new_n655), .B2(new_n603), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n478), .A2(new_n652), .A3(new_n595), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G119), .ZN(G21));
  NOR2_X1   g473(.A1(new_n444), .A2(new_n452), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n473), .A2(new_n439), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n455), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n554), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n573), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n625), .A2(KEYINPUT104), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n625), .A2(KEYINPUT104), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n665), .A2(new_n645), .A3(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n663), .A2(new_n512), .A3(new_n664), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G122), .ZN(G24));
  INV_X1    g483(.A(new_n502), .ZN(new_n670));
  INV_X1    g484(.A(new_n503), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n508), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n593), .B1(new_n672), .B2(new_n505), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n554), .A2(new_n673), .A3(new_n662), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n634), .A2(new_n632), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n674), .A2(KEYINPUT105), .A3(new_n675), .A4(new_n657), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n453), .B2(G902), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n458), .A2(new_n460), .A3(new_n661), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n454), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n675), .A2(new_n678), .A3(new_n680), .A4(new_n595), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n653), .A2(new_n656), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G125), .ZN(G27));
  NOR2_X1   g499(.A1(new_n278), .A2(new_n281), .ZN(new_n686));
  AND4_X1   g500(.A1(new_n550), .A2(new_n686), .A3(new_n632), .A4(new_n634), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(KEYINPUT32), .B1(new_n461), .B2(new_n454), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(KEYINPUT107), .B2(new_n462), .ZN(new_n690));
  OAI211_X1 g504(.A(KEYINPUT107), .B(new_n398), .C1(new_n453), .C2(new_n455), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n477), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n512), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g509(.A(KEYINPUT108), .B(new_n512), .C1(new_n690), .C2(new_n692), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n688), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n478), .A2(new_n687), .A3(new_n512), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n698), .A2(KEYINPUT106), .A3(new_n699), .ZN(new_n703));
  AOI22_X1  g517(.A1(new_n697), .A2(KEYINPUT42), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n292), .ZN(G33));
  NAND2_X1  g519(.A1(new_n478), .A2(new_n512), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n602), .ZN(new_n707));
  INV_X1    g521(.A(new_n686), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n708), .A2(new_n581), .A3(new_n606), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G134), .ZN(G36));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n345), .A2(new_n712), .A3(new_n568), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n344), .B(new_n714), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n715), .A2(new_n568), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n713), .B1(new_n716), .B2(new_n712), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n717), .A2(new_n556), .A3(new_n673), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(KEYINPUT44), .ZN(new_n719));
  OR2_X1    g533(.A1(new_n719), .A2(KEYINPUT111), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n708), .B1(new_n718), .B2(KEYINPUT44), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(KEYINPUT111), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n547), .B1(new_n548), .B2(new_n529), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n515), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT109), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n727), .B2(new_n726), .ZN(new_n730));
  INV_X1    g544(.A(new_n516), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n730), .A2(KEYINPUT46), .A3(new_n731), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n644), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n513), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n620), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n720), .A2(KEYINPUT112), .A3(new_n721), .A4(new_n722), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n725), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G137), .ZN(G39));
  INV_X1    g556(.A(KEYINPUT47), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n736), .A2(KEYINPUT47), .A3(new_n513), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n675), .A3(new_n686), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n478), .A2(new_n512), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G140), .ZN(G42));
  NAND2_X1  g565(.A1(new_n695), .A2(new_n696), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n708), .A2(new_n348), .A3(new_n655), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n713), .B(new_n753), .C1(new_n716), .C2(new_n712), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT48), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n619), .A2(new_n512), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n753), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n757), .B(new_n346), .C1(new_n569), .C2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n663), .A2(new_n512), .A3(new_n347), .A4(new_n346), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n717), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n642), .A2(new_n644), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n513), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n686), .B(new_n762), .C1(new_n746), .C2(new_n764), .ZN(new_n765));
  OR3_X1    g579(.A1(new_n759), .A2(new_n344), .A3(new_n568), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n755), .A2(new_n674), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n627), .A2(new_n279), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n655), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n762), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n770), .A2(new_n771), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(new_n775));
  OR3_X1    g589(.A1(new_n768), .A2(KEYINPUT51), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT51), .B1(new_n768), .B2(new_n775), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n760), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n665), .A2(new_n666), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n595), .A2(new_n602), .A3(new_n603), .A4(new_n606), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n618), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n608), .A2(new_n636), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n782), .A3(new_n684), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n781), .A2(new_n782), .A3(new_n684), .A4(KEYINPUT114), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n785), .A2(KEYINPUT52), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT52), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND4_X1   g603(.A1(new_n395), .A2(new_n578), .A3(new_n327), .A4(new_n580), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n478), .A2(new_n595), .A3(new_n631), .A4(new_n790), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n602), .B(new_n708), .C1(new_n791), .C2(new_n681), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n569), .B1(new_n395), .B2(new_n344), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n351), .B(new_n793), .C1(new_n280), .C2(new_n282), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n596), .B(new_n551), .C1(new_n557), .C2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n646), .A2(new_n650), .A3(new_n668), .A4(new_n658), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n792), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  AOI211_X1 g611(.A(new_n699), .B(new_n688), .C1(new_n695), .C2(new_n696), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n702), .A2(new_n703), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n797), .B(new_n710), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT53), .B1(new_n789), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n608), .A2(new_n636), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n683), .B2(new_n676), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n804), .B1(new_n806), .B2(new_n781), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n800), .A2(new_n788), .A3(new_n803), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n802), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(KEYINPUT115), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT114), .B1(new_n806), .B2(new_n781), .ZN(new_n813));
  INV_X1    g627(.A(new_n786), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n804), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n785), .A2(KEYINPUT52), .A3(new_n786), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n801), .A2(KEYINPUT53), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n800), .A2(new_n788), .A3(new_n807), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n817), .B1(new_n818), .B2(KEYINPUT53), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n812), .B1(new_n819), .B2(KEYINPUT54), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n815), .A2(new_n816), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n803), .B1(new_n821), .B2(new_n800), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n788), .A2(new_n807), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n801), .A3(KEYINPUT53), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(KEYINPUT54), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n778), .B(new_n811), .C1(new_n820), .C2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n761), .A2(new_n682), .A3(new_n717), .ZN(new_n828));
  OAI22_X1  g642(.A1(new_n827), .A2(new_n828), .B1(G952), .B2(G953), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n627), .A2(new_n514), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n281), .B1(new_n763), .B2(KEYINPUT49), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n830), .A2(new_n716), .A3(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n758), .B(new_n832), .C1(KEYINPUT49), .C2(new_n763), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n829), .A2(new_n833), .ZN(G75));
  NAND3_X1  g648(.A1(new_n825), .A2(G210), .A3(G902), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n226), .A2(new_n258), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(new_n256), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT55), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n835), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n839), .B1(new_n835), .B2(new_n836), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n252), .A2(G952), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(G51));
  NAND2_X1  g657(.A1(new_n731), .A2(KEYINPUT57), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n825), .A2(KEYINPUT54), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n844), .B1(new_n846), .B2(new_n826), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n731), .A2(KEYINPUT57), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n643), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OR3_X1    g663(.A1(new_n809), .A2(new_n260), .A3(new_n730), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n842), .B1(new_n849), .B2(new_n850), .ZN(G54));
  NAND2_X1  g665(.A1(KEYINPUT58), .A2(G475), .ZN(new_n852));
  AOI211_X1 g666(.A(new_n260), .B(new_n852), .C1(new_n822), .C2(new_n824), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n842), .B1(new_n853), .B2(new_n337), .ZN(new_n854));
  INV_X1    g668(.A(new_n852), .ZN(new_n855));
  OAI211_X1 g669(.A(G902), .B(new_n855), .C1(new_n802), .C2(new_n808), .ZN(new_n856));
  INV_X1    g670(.A(new_n337), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n856), .A2(KEYINPUT117), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT117), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n854), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT118), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n854), .B(new_n862), .C1(new_n858), .C2(new_n859), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n863), .ZN(G60));
  OAI21_X1  g678(.A(new_n811), .B1(new_n820), .B2(new_n826), .ZN(new_n865));
  XNOR2_X1  g679(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n393), .A2(new_n260), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n866), .B(new_n867), .Z(new_n868));
  AOI21_X1  g682(.A(new_n561), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n561), .ZN(new_n870));
  INV_X1    g684(.A(new_n868), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n809), .A2(new_n810), .ZN(new_n872));
  AOI211_X1 g686(.A(new_n870), .B(new_n871), .C1(new_n872), .C2(new_n845), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n869), .A2(new_n842), .A3(new_n873), .ZN(G63));
  XNOR2_X1  g688(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n384), .A2(new_n260), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n875), .B(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n822), .B2(new_n824), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n842), .B1(new_n879), .B2(new_n587), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n500), .A2(new_n501), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT121), .Z(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(new_n809), .B2(new_n878), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n880), .B(new_n883), .C1(new_n884), .C2(KEYINPUT61), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(KEYINPUT61), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT123), .Z(new_n887));
  XNOR2_X1  g701(.A(new_n885), .B(new_n887), .ZN(G66));
  NAND2_X1  g702(.A1(new_n349), .A2(G224), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(G953), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n795), .A2(new_n796), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n890), .B1(new_n891), .B2(G953), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n837), .B1(G898), .B2(new_n252), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n892), .B(new_n893), .ZN(G69));
  OAI21_X1  g708(.A(new_n710), .B1(new_n747), .B2(new_n749), .ZN(new_n895));
  AND4_X1   g709(.A1(new_n572), .A2(new_n738), .A3(new_n779), .A4(new_n752), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n895), .A2(new_n704), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n740), .A2(new_n898), .A3(new_n806), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n740), .B2(new_n806), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n897), .B(new_n252), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n430), .A2(new_n433), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n330), .A2(new_n331), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n902), .B(new_n903), .Z(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(G900), .B2(G953), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n750), .A2(new_n740), .ZN(new_n906));
  INV_X1    g720(.A(new_n706), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n907), .A2(new_n621), .A3(new_n686), .A4(new_n793), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n628), .A2(KEYINPUT62), .A3(new_n806), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT62), .B1(new_n628), .B2(new_n806), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n252), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n901), .A2(new_n905), .B1(new_n912), .B2(new_n904), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n901), .B2(new_n905), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n252), .B1(G227), .B2(G900), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n901), .A2(new_n905), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n912), .A2(new_n904), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n918), .B(new_n919), .C1(KEYINPUT124), .C2(new_n916), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n917), .A2(new_n921), .ZN(G72));
  NOR4_X1   g736(.A1(new_n906), .A2(new_n795), .A3(new_n911), .A4(new_n796), .ZN(new_n923));
  XNOR2_X1  g737(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n553), .A2(new_n260), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n924), .B(new_n925), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n439), .B(new_n463), .C1(new_n923), .C2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n457), .A2(new_n467), .A3(new_n469), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n819), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n928), .B(new_n930), .C1(G952), .C2(new_n252), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n897), .B(new_n891), .C1(new_n899), .C2(new_n900), .ZN(new_n932));
  AOI211_X1 g746(.A(new_n439), .B(new_n463), .C1(new_n932), .C2(new_n926), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n931), .A2(new_n933), .ZN(G57));
endmodule


