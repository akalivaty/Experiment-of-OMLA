//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  AOI21_X1  g005(.A(G128), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT64), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n188), .A2(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n197), .B(new_n198), .C1(new_n199), .C2(G128), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n202), .A2(new_n189), .A3(new_n191), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n195), .A2(new_n200), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G137), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n206), .A2(G137), .ZN(new_n209));
  OAI21_X1  g023(.A(G131), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n206), .B2(G137), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT11), .A3(G134), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n212), .A2(new_n214), .A3(new_n215), .A4(new_n207), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n205), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g032(.A(G116), .B(G119), .Z(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT2), .B(G113), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT65), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g035(.A(KEYINPUT2), .B(G113), .Z(new_n222));
  XNOR2_X1  g036(.A(G116), .B(G119), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n221), .A2(new_n225), .B1(new_n219), .B2(new_n220), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n199), .A2(KEYINPUT0), .A3(G128), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  OR2_X1    g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n190), .A2(G146), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n228), .B(new_n229), .C1(new_n230), .C2(new_n196), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n212), .A2(new_n207), .A3(new_n214), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G131), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n216), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n218), .A2(new_n226), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n226), .B1(new_n218), .B2(new_n236), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT28), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n218), .A2(new_n226), .A3(new_n236), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT28), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n243));
  INV_X1    g057(.A(G210), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n244), .A2(G237), .A3(G953), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n243), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g060(.A(KEYINPUT26), .B(G101), .Z(new_n247));
  AND2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n246), .A2(new_n247), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n239), .A2(KEYINPUT29), .A3(new_n242), .A4(new_n250), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n239), .A2(new_n242), .A3(new_n250), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT29), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n218), .A2(new_n236), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n255), .B1(new_n232), .B2(new_n235), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n226), .B1(new_n218), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n237), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n253), .B1(new_n259), .B2(new_n250), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n187), .B(new_n251), .C1(new_n252), .C2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT68), .A3(G472), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT68), .B1(new_n261), .B2(G472), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n240), .A2(new_n250), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n256), .B2(new_n258), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT31), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n239), .A2(new_n242), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n246), .B(new_n247), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n267), .A2(new_n268), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n205), .A2(new_n217), .B1(new_n232), .B2(new_n235), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n271), .B1(new_n226), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n218), .A2(new_n257), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n219), .A2(new_n220), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n219), .A2(KEYINPUT65), .A3(new_n220), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n224), .B1(new_n222), .B2(new_n223), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n274), .A2(KEYINPUT30), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n275), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT67), .A3(KEYINPUT31), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n269), .A2(new_n272), .A3(new_n273), .A4(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT32), .ZN(new_n286));
  NOR2_X1   g100(.A1(G472), .A2(G902), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n286), .B1(new_n285), .B2(new_n287), .ZN(new_n289));
  OAI22_X1  g103(.A1(new_n263), .A2(new_n264), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT9), .B(G234), .ZN(new_n291));
  OAI21_X1  g105(.A(G221), .B1(new_n291), .B2(G902), .ZN(new_n292));
  XOR2_X1   g106(.A(new_n292), .B(KEYINPUT74), .Z(new_n293));
  INV_X1    g107(.A(G104), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT3), .B1(new_n294), .B2(G107), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n296));
  INV_X1    g110(.A(G107), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(G104), .ZN(new_n298));
  INV_X1    g112(.A(G101), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n294), .A2(G107), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n295), .A2(new_n298), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n294), .A2(G107), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n297), .A2(G104), .ZN(new_n303));
  OAI21_X1  g117(.A(G101), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT10), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n205), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n295), .A2(new_n298), .A3(new_n300), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G101), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(KEYINPUT4), .A3(new_n301), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT4), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT76), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT76), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT4), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n299), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n309), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n311), .A2(new_n232), .A3(new_n317), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n203), .A2(new_n192), .A3(new_n194), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n306), .B1(new_n319), .B2(new_n305), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n308), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n235), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n323));
  INV_X1    g137(.A(new_n235), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n308), .A2(new_n318), .A3(new_n320), .A4(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(G110), .B(G140), .ZN(new_n327));
  INV_X1    g141(.A(G227), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(G953), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n327), .B(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n321), .A2(KEYINPUT78), .A3(new_n235), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n326), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n197), .B1(new_n199), .B2(G128), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n301), .B(new_n304), .C1(new_n333), .C2(new_n203), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n195), .A2(new_n200), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n305), .A2(new_n204), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n235), .ZN(new_n338));
  XOR2_X1   g152(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n330), .ZN(new_n341));
  NOR2_X1   g155(.A1(KEYINPUT77), .A2(KEYINPUT12), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n337), .A2(new_n235), .A3(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n340), .A2(new_n341), .A3(new_n325), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n332), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G469), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n187), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(G902), .B1(new_n332), .B2(new_n344), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(KEYINPUT79), .A3(new_n346), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n325), .A2(new_n323), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n317), .A2(new_n227), .A3(new_n231), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n354), .A2(new_n311), .B1(new_n334), .B2(new_n306), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n324), .B1(new_n355), .B2(new_n308), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n331), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n341), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n340), .A2(new_n325), .A3(new_n343), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n330), .B(KEYINPUT75), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n346), .B1(new_n363), .B2(new_n187), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n293), .B1(new_n352), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G140), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G125), .ZN(new_n368));
  INV_X1    g182(.A(G125), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G140), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT71), .ZN(new_n371));
  OR3_X1    g185(.A1(new_n369), .A2(KEYINPUT71), .A3(G140), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT72), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT16), .ZN(new_n375));
  INV_X1    g189(.A(new_n368), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT16), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n371), .B2(new_n372), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n380), .A2(new_n374), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n188), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(G237), .A2(G953), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(G143), .A3(G214), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(G143), .B1(new_n383), .B2(G214), .ZN(new_n386));
  OAI21_X1  g200(.A(G131), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT17), .ZN(new_n388));
  INV_X1    g202(.A(G237), .ZN(new_n389));
  INV_X1    g203(.A(G953), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(G214), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n190), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n215), .A3(new_n384), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n387), .A2(new_n388), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n384), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(KEYINPUT17), .A3(G131), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n369), .A2(KEYINPUT71), .A3(G140), .ZN(new_n398));
  XNOR2_X1  g212(.A(G125), .B(G140), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(KEYINPUT71), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT72), .B1(new_n400), .B2(new_n377), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n401), .A2(G146), .A3(new_n378), .A4(new_n375), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n382), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G113), .B(G122), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(new_n294), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n399), .A2(new_n188), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n373), .B2(new_n188), .ZN(new_n407));
  NAND2_X1  g221(.A1(KEYINPUT18), .A2(G131), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n392), .A2(new_n384), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n395), .A2(KEYINPUT18), .A3(G131), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n403), .A2(new_n405), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n368), .A2(new_n370), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT19), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n400), .B2(new_n414), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n416), .A2(new_n188), .B1(new_n387), .B2(new_n393), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n402), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n411), .ZN(new_n419));
  INV_X1    g233(.A(new_n405), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n412), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(G475), .A2(G902), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT20), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n422), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  INV_X1    g241(.A(new_n412), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n405), .B1(new_n403), .B2(new_n411), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n187), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n425), .A2(new_n427), .B1(G475), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n190), .A2(G128), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n201), .A2(G143), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n433), .A3(new_n206), .ZN(new_n434));
  XNOR2_X1  g248(.A(G116), .B(G122), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(new_n297), .ZN(new_n436));
  INV_X1    g250(.A(G122), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G116), .ZN(new_n438));
  INV_X1    g252(.A(G116), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G122), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n438), .A2(new_n440), .A3(new_n297), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n434), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n190), .A2(G128), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT13), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(new_n432), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n201), .A2(G143), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT13), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n206), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n435), .A2(new_n297), .ZN(new_n449));
  INV_X1    g263(.A(new_n434), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n206), .B1(new_n432), .B2(new_n433), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT14), .ZN(new_n453));
  OAI21_X1  g267(.A(G107), .B1(new_n440), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(new_n453), .B2(new_n435), .ZN(new_n455));
  OAI22_X1  g269(.A1(new_n442), .A2(new_n448), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G217), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n291), .A2(new_n457), .A3(G953), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n458), .ZN(new_n460));
  OAI221_X1 g274(.A(new_n460), .B1(new_n452), .B2(new_n455), .C1(new_n448), .C2(new_n442), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n461), .A3(new_n187), .ZN(new_n462));
  INV_X1    g276(.A(G478), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(KEYINPUT15), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n464), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n459), .A2(new_n461), .A3(new_n187), .A4(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n431), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G214), .B1(G237), .B2(G902), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT80), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n390), .A2(G952), .ZN(new_n472));
  INV_X1    g286(.A(G234), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n472), .B1(new_n473), .B2(new_n389), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(G902), .B(G953), .C1(new_n473), .C2(new_n389), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(KEYINPUT84), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT21), .B(G898), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n280), .A2(new_n311), .A3(new_n317), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n439), .A2(KEYINPUT5), .A3(G119), .ZN(new_n482));
  INV_X1    g296(.A(G113), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n223), .A2(KEYINPUT5), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n221), .A2(new_n225), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n305), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n481), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G110), .B(G122), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n481), .A2(new_n490), .A3(new_n488), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(KEYINPUT6), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n495), .A3(new_n491), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n232), .A2(new_n369), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n390), .A2(G224), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(KEYINPUT81), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n195), .A2(new_n200), .A3(new_n204), .A4(new_n369), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n497), .B2(new_n500), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n494), .A2(new_n496), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT7), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n506), .B1(new_n497), .B2(new_n500), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n221), .A2(new_n225), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n508), .A2(new_n277), .B1(new_n309), .B2(new_n316), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n509), .A2(new_n311), .B1(new_n487), .B2(new_n486), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n507), .B1(new_n510), .B2(new_n490), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n500), .B(new_n506), .C1(new_n369), .C2(new_n232), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n485), .A2(new_n484), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n508), .A2(new_n305), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n490), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT83), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n485), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n223), .A2(KEYINPUT83), .A3(KEYINPUT5), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n484), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n305), .B1(new_n521), .B2(new_n508), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n512), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(G902), .B1(new_n511), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(G210), .B1(G237), .B2(G902), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n504), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n526), .B1(new_n504), .B2(new_n525), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n471), .B(new_n480), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n468), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT22), .B(G137), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n390), .A2(G221), .A3(G234), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n201), .A2(G119), .ZN(new_n535));
  INV_X1    g349(.A(G119), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G128), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT24), .B(G110), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT70), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT23), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n536), .B2(G128), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n537), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT69), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT69), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n543), .A2(new_n544), .A3(new_n547), .A4(new_n537), .ZN(new_n548));
  AND4_X1   g362(.A1(new_n541), .A2(new_n546), .A3(G110), .A4(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G110), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n550), .B1(new_n545), .B2(KEYINPUT69), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n541), .B1(new_n551), .B2(new_n548), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n540), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n382), .B2(new_n402), .ZN(new_n554));
  OR2_X1    g368(.A1(new_n545), .A2(G110), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n538), .A2(new_n539), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n555), .A2(new_n556), .B1(new_n188), .B2(new_n399), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n402), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n534), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n546), .A2(G110), .A3(new_n548), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT70), .ZN(new_n562));
  INV_X1    g376(.A(new_n402), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n380), .A2(new_n374), .B1(new_n377), .B2(new_n376), .ZN(new_n564));
  AOI21_X1  g378(.A(G146), .B1(new_n564), .B2(new_n401), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n562), .B(new_n540), .C1(new_n563), .C2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(new_n558), .A3(new_n533), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n560), .A2(new_n567), .A3(new_n187), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT73), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT25), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n457), .B1(G234), .B2(new_n187), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n568), .A2(new_n570), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n560), .A2(new_n567), .A3(KEYINPUT25), .A4(new_n187), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(KEYINPUT73), .A3(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n560), .A2(new_n567), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n572), .A2(G902), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n573), .A2(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n290), .A2(new_n366), .A3(new_n530), .A4(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(G101), .ZN(G3));
  NAND2_X1  g395(.A1(new_n285), .A2(new_n287), .ZN(new_n582));
  INV_X1    g396(.A(G472), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n285), .B2(new_n187), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT85), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI211_X1 g400(.A(KEYINPUT85), .B(new_n583), .C1(new_n285), .C2(new_n187), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n579), .A3(new_n366), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n426), .B1(new_n422), .B2(new_n423), .ZN(new_n590));
  INV_X1    g404(.A(new_n423), .ZN(new_n591));
  AOI211_X1 g405(.A(KEYINPUT20), .B(new_n591), .C1(new_n412), .C2(new_n421), .ZN(new_n592));
  INV_X1    g406(.A(G475), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n403), .A2(new_n411), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n420), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n595), .B2(new_n412), .ZN(new_n596));
  OAI22_X1  g410(.A1(new_n590), .A2(new_n592), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT87), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT86), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n456), .A2(new_n599), .A3(new_n460), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT33), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n460), .B1(new_n456), .B2(new_n599), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n456), .A2(new_n599), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n458), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n605), .A2(KEYINPUT87), .A3(KEYINPUT33), .A4(new_n600), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n459), .A2(new_n461), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n463), .A2(G902), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n603), .A2(new_n606), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n462), .A2(new_n463), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n610), .A2(KEYINPUT88), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT88), .B1(new_n610), .B2(new_n611), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n597), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n469), .B(new_n480), .C1(new_n527), .C2(new_n528), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n589), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT34), .B(G104), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  INV_X1    g432(.A(KEYINPUT89), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n425), .A2(new_n619), .A3(new_n427), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n592), .A2(KEYINPUT89), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT90), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n596), .B2(new_n593), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n430), .A2(KEYINPUT90), .A3(G475), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n465), .A2(new_n467), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n615), .A2(new_n622), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n589), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT35), .B(G107), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  AOI21_X1  g446(.A(KEYINPUT67), .B1(new_n283), .B2(KEYINPUT31), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n256), .A2(new_n258), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n265), .B(new_n268), .C1(new_n634), .C2(new_n275), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n270), .A2(new_n271), .B1(new_n267), .B2(new_n268), .ZN(new_n637));
  AOI21_X1  g451(.A(G902), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT85), .B1(new_n638), .B2(new_n583), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n584), .A2(new_n585), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(new_n582), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n566), .A2(new_n558), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n534), .A2(KEYINPUT36), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n642), .B(new_n643), .Z(new_n644));
  INV_X1    g458(.A(new_n578), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n573), .B2(new_n576), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT91), .B1(new_n641), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT91), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n574), .A2(KEYINPUT73), .A3(new_n575), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n571), .A2(new_n572), .ZN(new_n651));
  OAI22_X1  g465(.A1(new_n650), .A2(new_n651), .B1(new_n645), .B2(new_n644), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n588), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n366), .A2(new_n530), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n648), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  AOI21_X1  g471(.A(new_n364), .B1(new_n349), .B2(new_n351), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n504), .A2(new_n525), .ZN(new_n659));
  INV_X1    g473(.A(new_n526), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n504), .A2(new_n525), .A3(new_n526), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n469), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n658), .A2(new_n664), .A3(new_n293), .ZN(new_n665));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n477), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n474), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n622), .A2(new_n627), .A3(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n665), .A2(new_n290), .A3(new_n652), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  INV_X1    g486(.A(new_n293), .ZN(new_n673));
  AND4_X1   g487(.A1(KEYINPUT79), .A2(new_n345), .A3(new_n346), .A4(new_n187), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT79), .B1(new_n350), .B2(new_n346), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n673), .B1(new_n676), .B2(new_n364), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n668), .B(KEYINPUT39), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT38), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n663), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n661), .A2(KEYINPUT38), .A3(new_n662), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n469), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n597), .A2(new_n626), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n237), .A2(new_n238), .A3(new_n250), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n691), .A2(G902), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n259), .A2(new_n271), .ZN(new_n693));
  OAI21_X1  g507(.A(G472), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n694), .B1(new_n288), .B2(new_n289), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n647), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n682), .A2(new_n689), .A3(new_n690), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  INV_X1    g513(.A(new_n664), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n290), .A2(new_n366), .A3(new_n700), .A4(new_n652), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n597), .B(new_n668), .C1(new_n613), .C2(new_n612), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT92), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n613), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n610), .A2(KEYINPUT88), .A3(new_n611), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n707), .A2(KEYINPUT92), .A3(new_n597), .A4(new_n668), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n701), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n188), .ZN(G48));
  OR2_X1    g525(.A1(new_n350), .A2(new_n346), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n673), .B(new_n712), .C1(new_n674), .C2(new_n675), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n614), .A2(new_n615), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n290), .A2(new_n714), .A3(new_n579), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT93), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND4_X1  g533(.A1(new_n290), .A2(new_n628), .A3(new_n714), .A4(new_n579), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NOR2_X1   g535(.A1(new_n713), .A2(new_n664), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n468), .A2(new_n479), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n290), .A3(new_n652), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  NAND2_X1  g539(.A1(new_n577), .A2(new_n578), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n726), .B1(new_n650), .B2(new_n651), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n637), .B1(new_n268), .B2(new_n267), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n287), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n638), .B2(new_n583), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n713), .A2(new_n615), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n688), .A2(KEYINPUT94), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT94), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n597), .A2(new_n734), .A3(new_n626), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n731), .A2(new_n732), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR2_X1   g552(.A1(new_n647), .A2(new_n730), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n739), .A2(new_n722), .A3(new_n704), .A4(new_n708), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT95), .B(G125), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G27));
  INV_X1    g556(.A(KEYINPUT97), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(new_n288), .B2(new_n289), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n582), .A2(KEYINPUT32), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(KEYINPUT97), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n252), .A2(new_n260), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n251), .A2(new_n187), .ZN(new_n749));
  OAI21_X1  g563(.A(G472), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT68), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n262), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n744), .A2(new_n747), .A3(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n754), .A2(new_n579), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n661), .A2(new_n673), .A3(new_n662), .A4(new_n469), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT96), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n326), .A2(new_n331), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n758), .B1(new_n759), .B2(new_n341), .ZN(new_n760));
  AOI211_X1 g574(.A(KEYINPUT96), .B(new_n330), .C1(new_n326), .C2(new_n331), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n362), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n346), .B1(new_n762), .B2(new_n187), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n757), .B1(new_n676), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n709), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n755), .A2(KEYINPUT98), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT98), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n754), .A2(new_n579), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n359), .A2(KEYINPUT96), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n759), .A2(new_n758), .A3(new_n341), .ZN(new_n771));
  AOI22_X1  g585(.A1(new_n770), .A2(new_n771), .B1(new_n360), .B2(new_n361), .ZN(new_n772));
  OAI21_X1  g586(.A(G469), .B1(new_n772), .B2(G902), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n756), .B1(new_n773), .B2(new_n352), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(KEYINPUT42), .A3(new_n704), .A4(new_n708), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n768), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n290), .A3(new_n579), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(new_n709), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n767), .A2(new_n776), .B1(new_n778), .B2(new_n765), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n215), .ZN(G33));
  NAND4_X1  g594(.A1(new_n774), .A2(new_n290), .A3(new_n670), .A4(new_n579), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G134), .ZN(G36));
  NAND3_X1  g596(.A1(new_n641), .A2(KEYINPUT100), .A3(new_n652), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n707), .A2(new_n431), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT43), .B1(new_n431), .B2(KEYINPUT99), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n707), .B(new_n431), .C1(KEYINPUT99), .C2(KEYINPUT43), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT100), .B1(new_n641), .B2(new_n652), .ZN(new_n791));
  OR3_X1    g605(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n346), .A2(new_n187), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n772), .A2(KEYINPUT45), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n346), .B1(new_n363), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n793), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT46), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n352), .B1(new_n797), .B2(KEYINPUT46), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n673), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n661), .A2(new_n662), .A3(new_n469), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n801), .A2(new_n679), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n790), .B1(new_n789), .B2(new_n791), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n792), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n801), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(KEYINPUT47), .B(new_n673), .C1(new_n799), .C2(new_n800), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n709), .A2(new_n290), .A3(new_n579), .A4(new_n802), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  OAI21_X1  g627(.A(new_n765), .B1(new_n777), .B2(new_n709), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT98), .B1(new_n755), .B2(new_n766), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n769), .A2(new_n775), .A3(new_n768), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n648), .A2(new_n653), .A3(new_n654), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT103), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n626), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT103), .B1(new_n465), .B2(new_n467), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n431), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n529), .B1(new_n614), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n588), .A2(new_n579), .A3(new_n366), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n724), .A3(new_n720), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n737), .A2(new_n580), .A3(new_n716), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n818), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n739), .A2(new_n774), .A3(new_n704), .A4(new_n708), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n781), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n745), .A2(new_n746), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n647), .B1(new_n753), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT104), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n820), .A2(new_n821), .A3(new_n669), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n834), .A2(new_n624), .A3(new_n625), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n620), .A2(new_n621), .ZN(new_n836));
  INV_X1    g650(.A(new_n802), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n832), .A2(new_n833), .A3(new_n366), .A4(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n366), .A2(new_n836), .A3(new_n837), .A4(new_n835), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n290), .A2(new_n652), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT104), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n830), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n817), .A2(new_n828), .A3(new_n843), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n290), .A2(new_n366), .A3(new_n700), .A4(new_n652), .ZN(new_n845));
  INV_X1    g659(.A(new_n709), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n669), .A2(KEYINPUT105), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n669), .A2(KEYINPUT105), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n673), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n676), .B2(new_n763), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n696), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n664), .B1(new_n733), .B2(new_n735), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n845), .A2(new_n846), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n671), .A2(new_n740), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n855), .A3(KEYINPUT106), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT106), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n849), .B1(new_n773), .B2(new_n352), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n853), .A2(new_n858), .A3(new_n647), .A4(new_n695), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(new_n701), .B2(new_n709), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n671), .A2(new_n740), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n857), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT52), .B1(new_n856), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n844), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT52), .B1(new_n860), .B2(new_n861), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT53), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n825), .A2(new_n724), .A3(new_n720), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n737), .A2(new_n580), .A3(new_n716), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n868), .A3(new_n655), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n842), .A2(new_n839), .ZN(new_n870));
  INV_X1    g684(.A(new_n830), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n779), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT52), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT106), .B1(new_n854), .B2(new_n855), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n860), .A2(new_n861), .A3(new_n857), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n856), .A2(new_n862), .A3(KEYINPUT52), .ZN(new_n878));
  AND4_X1   g692(.A1(KEYINPUT53), .A2(new_n873), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT54), .B1(new_n866), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n873), .A2(new_n877), .A3(KEYINPUT53), .A4(new_n865), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n873), .A2(new_n877), .A3(new_n878), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(KEYINPUT53), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n727), .A2(new_n474), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n713), .A2(new_n802), .ZN(new_n886));
  INV_X1    g700(.A(new_n695), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n707), .A2(new_n597), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(KEYINPUT109), .A3(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n886), .A2(new_n885), .A3(new_n887), .A4(new_n889), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT109), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n474), .B1(new_n786), .B2(new_n787), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n894), .A2(new_n886), .ZN(new_n895));
  AOI22_X1  g709(.A1(new_n890), .A2(new_n893), .B1(new_n739), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT108), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n686), .A2(new_n687), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n898), .B1(new_n899), .B2(new_n713), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n714), .A2(KEYINPUT108), .A3(new_n686), .A4(new_n687), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n901), .A3(new_n894), .A4(new_n731), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT50), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT110), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT50), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n902), .B(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT110), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n907), .A3(new_n896), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n352), .A2(new_n712), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT101), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n352), .A2(KEYINPUT101), .A3(new_n712), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT107), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT107), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n911), .A2(new_n916), .A3(new_n913), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n915), .A2(new_n293), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n808), .A2(new_n918), .A3(new_n809), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n894), .A2(new_n731), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n920), .A2(new_n837), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n904), .A2(KEYINPUT51), .A3(new_n908), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n920), .A2(new_n722), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n888), .A2(new_n597), .A3(new_n707), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n924), .A2(new_n472), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n895), .A2(new_n755), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n927), .A2(KEYINPUT48), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(KEYINPUT48), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n922), .A2(new_n906), .A3(new_n896), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT51), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n923), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n880), .A2(new_n884), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(G952), .A2(G953), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT111), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n912), .A2(new_n914), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n939), .A2(KEYINPUT49), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(KEYINPUT49), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n686), .A2(new_n673), .A3(new_n471), .ZN(new_n942));
  NOR4_X1   g756(.A1(new_n942), .A2(new_n727), .A3(new_n695), .A4(new_n784), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT102), .Z(new_n945));
  NAND2_X1  g759(.A1(new_n938), .A2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT112), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n938), .A2(KEYINPUT112), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(G75));
  NOR2_X1   g764(.A1(new_n390), .A2(G952), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT115), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n864), .A2(new_n878), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT53), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI211_X1 g769(.A(new_n244), .B(new_n187), .C1(new_n955), .C2(new_n882), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n494), .A2(new_n496), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(new_n503), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT55), .Z(new_n959));
  INV_X1    g773(.A(KEYINPUT114), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT56), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n959), .A2(new_n960), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n952), .B1(new_n956), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT113), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n956), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n955), .A2(new_n882), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n968), .A2(G210), .A3(G902), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(KEYINPUT113), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n967), .A2(new_n970), .A3(new_n962), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n965), .B1(new_n971), .B2(new_n959), .ZN(G51));
  XNOR2_X1  g786(.A(new_n793), .B(KEYINPUT57), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n881), .B1(new_n955), .B2(new_n882), .ZN(new_n974));
  INV_X1    g788(.A(new_n884), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n345), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n968), .A2(G902), .A3(new_n794), .A4(new_n796), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n951), .B1(new_n977), .B2(new_n978), .ZN(G54));
  AND2_X1   g793(.A1(KEYINPUT58), .A2(G475), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n968), .A2(G902), .A3(new_n422), .A4(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT116), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n968), .A2(G902), .A3(new_n980), .ZN(new_n985));
  INV_X1    g799(.A(new_n422), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n951), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n983), .A2(new_n984), .A3(new_n987), .ZN(G60));
  AND3_X1   g802(.A1(new_n603), .A2(new_n606), .A3(new_n608), .ZN(new_n989));
  NAND2_X1  g803(.A1(G478), .A2(G902), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT59), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n989), .B(new_n991), .C1(new_n974), .C2(new_n975), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n952), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n880), .A2(new_n884), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n989), .B1(new_n994), .B2(new_n991), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n993), .A2(new_n995), .ZN(G63));
  INV_X1    g810(.A(KEYINPUT61), .ZN(new_n997));
  NAND2_X1  g811(.A1(G217), .A2(G902), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT60), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(new_n955), .B2(new_n882), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n644), .B(KEYINPUT117), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n577), .B(KEYINPUT118), .Z(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n952), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n997), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1008), .A2(new_n1002), .A3(KEYINPUT61), .A4(new_n952), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(G66));
  NOR2_X1   g824(.A1(new_n828), .A2(G953), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1011), .B(KEYINPUT119), .ZN(new_n1012));
  INV_X1    g826(.A(G224), .ZN(new_n1013));
  OAI21_X1  g827(.A(G953), .B1(new_n478), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n957), .B1(G898), .B2(new_n390), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(G69));
  OR3_X1    g831(.A1(new_n861), .A2(new_n710), .A3(KEYINPUT121), .ZN(new_n1018));
  OAI21_X1  g832(.A(KEYINPUT121), .B1(new_n861), .B2(new_n710), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n805), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT123), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n805), .A2(KEYINPUT123), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OR2_X1    g838(.A1(new_n801), .A2(new_n679), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n755), .A2(new_n853), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n812), .B(new_n781), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1027), .A2(new_n779), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1024), .A2(new_n390), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n256), .A2(new_n276), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1030), .B(new_n416), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1031), .B1(G900), .B2(G953), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1018), .A2(new_n698), .A3(new_n1019), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT62), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n1018), .A2(new_n698), .A3(KEYINPUT62), .A4(new_n1019), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n802), .B1(new_n614), .B2(new_n823), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n680), .A2(new_n290), .A3(new_n579), .A4(new_n1039), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n805), .A2(new_n812), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g855(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(KEYINPUT122), .ZN(new_n1044));
  INV_X1    g858(.A(KEYINPUT122), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1038), .A2(new_n1045), .A3(new_n1042), .ZN(new_n1046));
  AOI21_X1  g860(.A(G953), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g861(.A(new_n1031), .B(KEYINPUT120), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1033), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g863(.A(G953), .B1(new_n328), .B2(new_n666), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n1050), .B1(new_n1048), .B2(KEYINPUT124), .ZN(new_n1051));
  XNOR2_X1  g865(.A(new_n1049), .B(new_n1051), .ZN(G72));
  NAND3_X1  g866(.A1(new_n1024), .A2(new_n828), .A3(new_n1028), .ZN(new_n1053));
  NAND2_X1  g867(.A1(G472), .A2(G902), .ZN(new_n1054));
  XOR2_X1   g868(.A(new_n1054), .B(KEYINPUT63), .Z(new_n1055));
  NAND2_X1  g869(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n634), .A2(new_n240), .ZN(new_n1057));
  NOR2_X1   g871(.A1(new_n1057), .A2(new_n250), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n951), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g873(.A(new_n879), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n864), .A2(new_n865), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1061), .A2(new_n954), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g877(.A(new_n1055), .ZN(new_n1064));
  AOI21_X1  g878(.A(KEYINPUT126), .B1(new_n1057), .B2(new_n271), .ZN(new_n1065));
  NOR2_X1   g879(.A1(new_n1065), .A2(new_n267), .ZN(new_n1066));
  NAND3_X1  g880(.A1(new_n1057), .A2(KEYINPUT126), .A3(new_n271), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n1064), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AND3_X1   g882(.A1(new_n1063), .A2(KEYINPUT127), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g883(.A(KEYINPUT127), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1070));
  OAI21_X1  g884(.A(new_n1059), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g885(.A(new_n693), .ZN(new_n1072));
  AOI211_X1 g886(.A(KEYINPUT122), .B(new_n1041), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1073));
  AOI21_X1  g887(.A(new_n1045), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1074));
  NOR2_X1   g888(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g889(.A(new_n1064), .B1(new_n1075), .B2(new_n828), .ZN(new_n1076));
  AOI21_X1  g890(.A(new_n1072), .B1(new_n1076), .B2(KEYINPUT125), .ZN(new_n1077));
  INV_X1    g891(.A(KEYINPUT125), .ZN(new_n1078));
  NOR3_X1   g892(.A1(new_n1073), .A2(new_n1074), .A3(new_n869), .ZN(new_n1079));
  OAI21_X1  g893(.A(new_n1078), .B1(new_n1079), .B2(new_n1064), .ZN(new_n1080));
  AOI21_X1  g894(.A(new_n1071), .B1(new_n1077), .B2(new_n1080), .ZN(G57));
endmodule


