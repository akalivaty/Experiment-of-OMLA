//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  INV_X1    g001(.A(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT11), .B(G169gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT12), .Z(new_n207));
  INV_X1    g006(.A(G22gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G15gat), .ZN(new_n209));
  INV_X1    g008(.A(G15gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G22gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT87), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G1gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G8gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(new_n212), .A3(G1gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n218), .B1(new_n217), .B2(new_n219), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT84), .ZN(new_n224));
  NAND2_X1  g023(.A1(G43gat), .A2(G50gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(G43gat), .A2(G50gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n224), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G43gat), .ZN(new_n229));
  INV_X1    g028(.A(G50gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(KEYINPUT84), .A3(new_n225), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(new_n232), .A3(KEYINPUT15), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT86), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n231), .A2(new_n225), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(KEYINPUT15), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G29gat), .ZN(new_n238));
  INV_X1    g037(.A(G36gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT14), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT14), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(G29gat), .B2(G36gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT85), .B(G29gat), .Z(new_n244));
  AOI21_X1  g043(.A(new_n243), .B1(G36gat), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n237), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT85), .B(G29gat), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n242), .B(new_n240), .C1(new_n247), .C2(new_n239), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT15), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n231), .A2(KEYINPUT86), .A3(new_n249), .A4(new_n225), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n233), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n223), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n213), .A2(new_n214), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n215), .A2(new_n216), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n219), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G8gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT88), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n258), .A2(new_n259), .A3(new_n220), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n259), .B1(new_n258), .B2(new_n220), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT17), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n249), .B1(new_n235), .B2(new_n224), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n245), .A2(new_n250), .B1(new_n232), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n248), .B1(new_n233), .B2(new_n236), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n246), .A2(KEYINPUT17), .A3(new_n252), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n254), .B1(new_n262), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G229gat), .A2(G233gat), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT18), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n265), .A2(new_n266), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n220), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n271), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT18), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n265), .A2(new_n266), .A3(new_n263), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT17), .B1(new_n246), .B2(new_n252), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT88), .B1(new_n221), .B2(new_n222), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n258), .A2(new_n259), .A3(new_n220), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n275), .B(new_n278), .C1(new_n281), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n223), .A2(new_n253), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n275), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n271), .B(KEYINPUT13), .Z(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n207), .B1(new_n272), .B2(new_n290), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n270), .A2(new_n278), .B1(new_n287), .B2(new_n288), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n275), .B1(new_n281), .B2(new_n284), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n277), .B1(new_n293), .B2(new_n276), .ZN(new_n294));
  INV_X1    g093(.A(new_n207), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n292), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n291), .A2(new_n296), .A3(KEYINPUT89), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT89), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n298), .B(new_n207), .C1(new_n272), .C2(new_n290), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT90), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n297), .A2(KEYINPUT90), .A3(new_n299), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(G1gat), .B(G29gat), .Z(new_n306));
  XNOR2_X1  g105(.A(G57gat), .B(G85gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n308), .B(new_n309), .Z(new_n310));
  INV_X1    g109(.A(KEYINPUT5), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n312));
  INV_X1    g111(.A(G113gat), .ZN(new_n313));
  INV_X1    g112(.A(G120gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316));
  NAND2_X1  g115(.A1(G113gat), .A2(G120gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n315), .A2(new_n317), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT66), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n318), .B(new_n319), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n317), .ZN(new_n323));
  NOR2_X1   g122(.A1(G113gat), .A2(G120gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(G127gat), .A2(G134gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(G127gat), .A2(G134gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n325), .B(new_n316), .C1(new_n328), .C2(KEYINPUT66), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n322), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT71), .B1(G155gat), .B2(G162gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G155gat), .B(G162gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT71), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G141gat), .ZN(new_n336));
  INV_X1    g135(.A(G148gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G141gat), .A2(G148gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT2), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n340), .A2(KEYINPUT72), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(KEYINPUT72), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n338), .B(new_n339), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n335), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n338), .A2(new_n339), .ZN(new_n345));
  INV_X1    g144(.A(G155gat), .ZN(new_n346));
  OR2_X1    g145(.A1(KEYINPUT73), .A2(G162gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(KEYINPUT73), .A2(G162gat), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n333), .B(new_n345), .C1(new_n349), .C2(new_n340), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n312), .B1(new_n330), .B2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(KEYINPUT73), .B(G162gat), .Z(new_n353));
  OAI21_X1  g152(.A(KEYINPUT2), .B1(new_n353), .B2(new_n346), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n333), .A2(new_n338), .A3(new_n339), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n354), .A2(new_n355), .B1(new_n335), .B2(new_n343), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n322), .A2(new_n329), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(KEYINPUT74), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n330), .A2(new_n351), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n352), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n311), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n352), .A2(new_n364), .A3(new_n358), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n357), .B1(new_n351), .B2(KEYINPUT3), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT3), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n356), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n362), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n356), .A2(KEYINPUT4), .A3(new_n357), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n365), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n363), .A2(new_n371), .ZN(new_n372));
  AND4_X1   g171(.A1(KEYINPUT74), .A2(new_n357), .A3(new_n350), .A4(new_n344), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT74), .B1(new_n356), .B2(new_n357), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT4), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n364), .B1(new_n330), .B2(new_n351), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n375), .A2(new_n369), .A3(new_n311), .A4(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n310), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G197gat), .B(G204gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT69), .B(G218gat), .ZN(new_n381));
  INV_X1    g180(.A(G211gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n380), .B1(new_n383), .B2(KEYINPUT22), .ZN(new_n384));
  XNOR2_X1  g183(.A(G211gat), .B(G218gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(KEYINPUT70), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n384), .B(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(G169gat), .A2(G176gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT26), .ZN(new_n390));
  NAND2_X1  g189(.A1(G183gat), .A2(G190gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT26), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(G169gat), .B2(G176gat), .ZN(new_n393));
  AND2_X1   g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n390), .B(new_n391), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT27), .B(G183gat), .ZN(new_n396));
  INV_X1    g195(.A(G190gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT28), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n396), .A2(KEYINPUT28), .A3(new_n397), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n395), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT65), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT24), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(G183gat), .A3(G190gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(G183gat), .B(G190gat), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n403), .B(new_n405), .C1(new_n406), .C2(new_n404), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT25), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n389), .A2(KEYINPUT23), .ZN(new_n410));
  INV_X1    g209(.A(new_n394), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G183gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(G190gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n397), .A2(G183gat), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n404), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n405), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n412), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT64), .B1(new_n389), .B2(KEYINPUT23), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT64), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT23), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n420), .B(new_n421), .C1(G169gat), .C2(G176gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n409), .A2(new_n418), .A3(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n397), .A2(G183gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n413), .A2(G190gat), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT24), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n394), .B1(KEYINPUT23), .B2(new_n389), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n423), .A2(new_n427), .A3(new_n405), .A4(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(new_n408), .A3(new_n407), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n402), .B1(new_n424), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(KEYINPUT29), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  AOI211_X1 g234(.A(new_n433), .B(new_n402), .C1(new_n424), .C2(new_n430), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n388), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n424), .A2(new_n430), .ZN(new_n438));
  INV_X1    g237(.A(new_n402), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n432), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n440), .B(new_n387), .C1(new_n431), .C2(new_n434), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n437), .A2(new_n441), .A3(new_n445), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(KEYINPUT30), .A3(new_n448), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n437), .A2(new_n441), .A3(new_n445), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n445), .B1(new_n437), .B2(new_n441), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT30), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n449), .A2(new_n453), .A3(KEYINPUT78), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT78), .B1(new_n449), .B2(new_n453), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n379), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n366), .A2(new_n368), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n375), .A2(new_n457), .A3(new_n376), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n362), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n459), .B(KEYINPUT39), .C1(new_n362), .C2(new_n360), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT39), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(new_n461), .A3(new_n362), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n462), .A2(KEYINPUT79), .A3(new_n310), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT79), .B1(new_n462), .B2(new_n310), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT40), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(KEYINPUT40), .B(new_n460), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT80), .B1(new_n456), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT78), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n442), .A2(KEYINPUT30), .A3(new_n446), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n449), .A2(new_n453), .A3(KEYINPUT78), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n378), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT80), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n468), .A4(new_n467), .ZN(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n378), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n372), .A2(new_n310), .A3(new_n377), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n479), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n483), .B2(new_n378), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n442), .A2(KEYINPUT37), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n446), .A2(KEYINPUT37), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n486), .B1(new_n451), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n450), .B1(new_n489), .B2(KEYINPUT38), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT38), .B1(new_n447), .B2(new_n487), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT81), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n437), .A2(new_n492), .A3(new_n441), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n493), .B(KEYINPUT37), .C1(new_n492), .C2(new_n441), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n491), .A2(KEYINPUT82), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT82), .B1(new_n491), .B2(new_n494), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n485), .B(new_n490), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n470), .A2(new_n478), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G228gat), .ZN(new_n499));
  INV_X1    g298(.A(G233gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT29), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n368), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n388), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n387), .A2(new_n502), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n356), .B1(new_n506), .B2(new_n367), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n501), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n384), .A2(new_n385), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT29), .B1(new_n384), .B2(new_n385), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT3), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI221_X1 g310(.A(new_n504), .B1(new_n499), .B2(new_n500), .C1(new_n356), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT31), .B(G50gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G78gat), .B(G106gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(G22gat), .ZN(new_n517));
  INV_X1    g316(.A(new_n514), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n508), .A2(new_n512), .A3(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n515), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n517), .B1(new_n515), .B2(new_n519), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT36), .ZN(new_n524));
  NAND2_X1  g323(.A1(G227gat), .A2(G233gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n431), .A2(new_n330), .ZN(new_n526));
  AOI211_X1 g325(.A(new_n357), .B(new_n402), .C1(new_n424), .C2(new_n430), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT34), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n525), .B2(KEYINPUT68), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n528), .B(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G43gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(G71gat), .B(G99gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n526), .A2(new_n527), .A3(new_n525), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT32), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n537), .A2(KEYINPUT33), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT67), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n438), .A2(new_n439), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n357), .ZN(new_n543));
  INV_X1    g342(.A(new_n525), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n431), .A2(new_n330), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n535), .B1(new_n546), .B2(KEYINPUT32), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT67), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT33), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n541), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n536), .A2(KEYINPUT33), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n546), .A2(KEYINPUT32), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n532), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  AOI211_X1 g355(.A(new_n556), .B(new_n531), .C1(new_n541), .C2(new_n551), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n524), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n548), .B1(new_n547), .B2(new_n550), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n554), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n531), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n552), .A2(new_n554), .A3(new_n532), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(KEYINPUT36), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n523), .B1(new_n558), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT35), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n474), .A2(new_n484), .A3(new_n475), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT83), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n555), .A2(new_n557), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n474), .A2(new_n484), .A3(KEYINPUT83), .A4(new_n475), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n569), .A2(new_n570), .A3(new_n522), .A4(new_n571), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n498), .A2(new_n565), .B1(new_n566), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n449), .A2(new_n453), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n484), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n575), .B(KEYINPUT77), .Z(new_n576));
  AOI21_X1  g375(.A(new_n522), .B1(new_n558), .B2(new_n564), .ZN(new_n577));
  AND4_X1   g376(.A1(KEYINPUT35), .A2(new_n522), .A3(new_n562), .A4(new_n563), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n305), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G183gat), .B(G211gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT94), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(new_n346), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n582), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G71gat), .B(G78gat), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT92), .B1(G57gat), .B2(G64gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT9), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(KEYINPUT91), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G57gat), .A2(G64gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n590), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(KEYINPUT91), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n588), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n589), .B1(G57gat), .B2(G64gat), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n587), .A4(new_n593), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT93), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n598), .A2(new_n601), .A3(KEYINPUT93), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n223), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT21), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n611), .B1(new_n602), .B2(new_n609), .ZN(new_n614));
  OR3_X1    g413(.A1(new_n613), .A2(G127gat), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(G127gat), .B1(new_n613), .B2(new_n614), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n608), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n608), .B1(new_n615), .B2(new_n616), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n586), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n615), .A2(new_n616), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(new_n223), .A3(new_n607), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(new_n617), .A3(new_n585), .ZN(new_n623));
  NAND2_X1  g422(.A1(G232gat), .A2(G233gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n624), .B(KEYINPUT95), .Z(new_n625));
  INV_X1    g424(.A(KEYINPUT41), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n631), .A2(G85gat), .A3(G92gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT97), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(G85gat), .ZN(new_n635));
  INV_X1    g434(.A(G92gat), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n633), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .A4(new_n631), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT7), .B1(new_n635), .B2(new_n636), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n634), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(G99gat), .A2(G106gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n645));
  NAND2_X1  g444(.A1(G99gat), .A2(G106gat), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n646), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT98), .B1(new_n648), .B2(new_n643), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AOI22_X1  g450(.A1(KEYINPUT8), .A2(new_n646), .B1(new_n635), .B2(new_n636), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n642), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n642), .B2(new_n652), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n269), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G190gat), .B(G218gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT99), .ZN(new_n659));
  OAI22_X1  g458(.A1(new_n655), .A2(new_n253), .B1(new_n626), .B2(new_n625), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n659), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n625), .A2(new_n626), .ZN(new_n663));
  INV_X1    g462(.A(new_n655), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n663), .B1(new_n664), .B2(new_n273), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n662), .B1(new_n665), .B2(new_n656), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n630), .B1(new_n661), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n659), .B1(new_n657), .B2(new_n660), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n665), .A2(new_n662), .A3(new_n656), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n629), .A3(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n620), .A2(new_n623), .A3(new_n667), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(G230gat), .A2(G233gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT101), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n675));
  OAI21_X1  g474(.A(new_n602), .B1(new_n653), .B2(new_n654), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n642), .A2(new_n652), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n650), .ZN(new_n678));
  INV_X1    g477(.A(new_n602), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n642), .A2(new_n651), .A3(new_n652), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n675), .B1(new_n676), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n605), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n655), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n674), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT102), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n687), .B(new_n674), .C1(new_n682), .C2(new_n684), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n676), .A2(new_n673), .A3(new_n681), .ZN(new_n689));
  XNOR2_X1  g488(.A(G120gat), .B(G148gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT103), .ZN(new_n691));
  XNOR2_X1  g490(.A(G176gat), .B(G204gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n691), .B(new_n692), .Z(new_n693));
  NOR2_X1   g492(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n686), .A2(new_n688), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n685), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n693), .B1(new_n696), .B2(new_n689), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n671), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n580), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n484), .A2(KEYINPUT104), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n484), .A2(KEYINPUT104), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT105), .B(G1gat), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1324gat));
  INV_X1    g506(.A(new_n700), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n474), .A2(new_n475), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT16), .B(G8gat), .Z(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n709), .ZN(new_n712));
  OAI21_X1  g511(.A(G8gat), .B1(new_n700), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  MUX2_X1   g513(.A(new_n711), .B(new_n714), .S(KEYINPUT42), .Z(G1325gat));
  AND2_X1   g514(.A1(new_n558), .A2(new_n564), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G15gat), .B1(new_n700), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n570), .A2(new_n210), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n700), .B2(new_n719), .ZN(G1326gat));
  NOR2_X1   g519(.A1(new_n700), .A2(new_n522), .ZN(new_n721));
  XOR2_X1   g520(.A(KEYINPUT43), .B(G22gat), .Z(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1327gat));
  INV_X1    g522(.A(new_n698), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n620), .A2(new_n623), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n667), .A2(new_n670), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT106), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n580), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n247), .A3(new_n703), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT45), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n498), .A2(new_n565), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n572), .A2(new_n566), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(new_n579), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n727), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT44), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n728), .B1(new_n573), .B2(new_n579), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n300), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n244), .B1(new_n744), .B2(new_n704), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n733), .A2(new_n745), .ZN(G1328gat));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n239), .A3(new_n709), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT46), .Z(new_n748));
  OAI21_X1  g547(.A(G36gat), .B1(new_n744), .B2(new_n712), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1329gat));
  INV_X1    g549(.A(new_n740), .ZN(new_n751));
  AOI211_X1 g550(.A(new_n728), .B(new_n751), .C1(new_n573), .C2(new_n579), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n736), .B2(new_n727), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n716), .B(new_n743), .C1(new_n752), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G43gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n731), .A2(new_n229), .A3(new_n570), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT108), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1330gat));
  OAI21_X1  g559(.A(G50gat), .B1(new_n744), .B2(new_n522), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n731), .A2(new_n230), .A3(new_n523), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT48), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n761), .B2(new_n762), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(G1331gat));
  INV_X1    g565(.A(new_n300), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n767), .A2(new_n671), .A3(new_n724), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n736), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n703), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g570(.A1(new_n769), .A2(new_n709), .ZN(new_n772));
  NOR2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  AND2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n772), .B2(new_n773), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT109), .ZN(G1333gat));
  NAND2_X1  g576(.A1(new_n769), .A2(new_n716), .ZN(new_n778));
  INV_X1    g577(.A(new_n570), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(G71gat), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n778), .A2(G71gat), .B1(new_n769), .B2(new_n780), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1334gat));
  NAND2_X1  g582(.A1(new_n769), .A2(new_n523), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G78gat), .ZN(G1335gat));
  INV_X1    g584(.A(new_n725), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n767), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n724), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n738), .B2(new_n741), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G85gat), .B1(new_n792), .B2(new_n704), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT51), .B1(new_n737), .B2(new_n788), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n739), .A2(new_n795), .A3(new_n787), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n703), .A2(new_n635), .A3(new_n698), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(G1336gat));
  NOR3_X1   g598(.A1(new_n712), .A2(G92gat), .A3(new_n724), .ZN(new_n800));
  OR2_X1    g599(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n739), .B2(new_n787), .ZN(new_n802));
  AND4_X1   g601(.A1(new_n736), .A2(new_n727), .A3(new_n787), .A4(new_n801), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n709), .B(new_n789), .C1(new_n752), .C2(new_n754), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n808), .A3(G92gat), .ZN(new_n809));
  OAI211_X1 g608(.A(KEYINPUT113), .B(new_n800), .C1(new_n802), .C2(new_n803), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n806), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n808), .B1(new_n807), .B2(G92gat), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT52), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n636), .B1(new_n791), .B2(new_n709), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n794), .A2(new_n796), .A3(new_n800), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n814), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n807), .A2(G92gat), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n820), .A2(KEYINPUT114), .A3(new_n817), .A4(new_n816), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n813), .A2(new_n822), .ZN(G1337gat));
  OAI21_X1  g622(.A(G99gat), .B1(new_n792), .B2(new_n717), .ZN(new_n824));
  OR3_X1    g623(.A1(new_n779), .A2(G99gat), .A3(new_n724), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n797), .B2(new_n825), .ZN(G1338gat));
  INV_X1    g625(.A(G106gat), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n791), .B2(new_n523), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n802), .A2(new_n803), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n522), .A2(G106gat), .A3(new_n724), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832));
  INV_X1    g631(.A(new_n830), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n797), .B2(new_n833), .ZN(new_n834));
  OAI22_X1  g633(.A1(new_n831), .A2(new_n832), .B1(new_n834), .B2(new_n828), .ZN(G1339gat));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n699), .A2(new_n836), .A3(new_n300), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n699), .B2(new_n300), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n682), .A2(new_n684), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n673), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n686), .A2(new_n841), .A3(KEYINPUT54), .A4(new_n688), .ZN(new_n842));
  INV_X1    g641(.A(new_n693), .ZN(new_n843));
  XOR2_X1   g642(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n696), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n842), .A2(KEYINPUT55), .A3(new_n845), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n695), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n270), .A2(new_n271), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n287), .A2(new_n288), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n206), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT117), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n855), .B(new_n206), .C1(new_n851), .C2(new_n852), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n727), .A2(new_n854), .A3(new_n296), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n850), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n698), .A2(new_n854), .A3(new_n296), .A4(new_n856), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n850), .B2(new_n300), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n858), .B1(new_n860), .B2(new_n728), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n839), .B1(new_n861), .B2(new_n786), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n779), .A2(new_n523), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n862), .A2(new_n863), .A3(new_n712), .A4(new_n703), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(new_n313), .A3(new_n305), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n862), .A2(new_n703), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n866), .A2(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n712), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n767), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n865), .B1(new_n870), .B2(new_n313), .ZN(G1340gat));
  NOR3_X1   g670(.A1(new_n864), .A2(new_n314), .A3(new_n724), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n698), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n314), .ZN(G1341gat));
  OAI21_X1  g673(.A(G127gat), .B1(new_n864), .B2(new_n725), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n725), .A2(G127gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n868), .B2(new_n876), .ZN(G1342gat));
  INV_X1    g676(.A(G134gat), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n709), .A2(new_n728), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT118), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n867), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n883), .B(new_n884), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n864), .A2(new_n728), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n882), .A2(KEYINPUT56), .B1(G134gat), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(G1343gat));
  AND2_X1   g687(.A1(new_n866), .A2(new_n577), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n712), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n304), .A2(new_n336), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892));
  OAI22_X1  g691(.A1(new_n890), .A2(new_n891), .B1(new_n892), .B2(KEYINPUT58), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n716), .A2(new_n704), .A3(new_n709), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n849), .A2(new_n695), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n302), .A2(new_n303), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT55), .B1(new_n842), .B2(new_n845), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT120), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n859), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n858), .B1(new_n899), .B2(new_n728), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n839), .B1(new_n900), .B2(new_n786), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n522), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(KEYINPUT121), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n862), .A2(new_n523), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n902), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT121), .B1(new_n901), .B2(new_n903), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n767), .B(new_n894), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT58), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n336), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n893), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n894), .B1(new_n907), .B2(new_n908), .ZN(new_n913));
  OAI21_X1  g712(.A(G141gat), .B1(new_n913), .B2(new_n305), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n890), .A2(new_n891), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(new_n892), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n912), .B1(new_n916), .B2(new_n910), .ZN(G1344gat));
  OAI211_X1 g716(.A(new_n698), .B(new_n894), .C1(new_n907), .C2(new_n908), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n337), .A2(KEYINPUT59), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT123), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n305), .A2(new_n699), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n922), .B1(new_n900), .B2(new_n786), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n522), .A2(KEYINPUT57), .ZN(new_n924));
  AOI22_X1  g723(.A1(new_n923), .A2(new_n924), .B1(new_n905), .B2(KEYINPUT57), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n894), .A2(new_n698), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n337), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT59), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT124), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n923), .A2(new_n924), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n905), .A2(KEYINPUT57), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n931), .A2(new_n932), .A3(new_n926), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n930), .B(KEYINPUT59), .C1(new_n933), .C2(new_n337), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n936), .A3(new_n919), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(new_n890), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n337), .A3(new_n698), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1345gat));
  OAI21_X1  g740(.A(G155gat), .B1(new_n913), .B2(new_n725), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n939), .A2(new_n346), .A3(new_n786), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1346gat));
  NAND3_X1  g743(.A1(new_n889), .A2(new_n353), .A3(new_n881), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n913), .A2(new_n728), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n946), .B2(new_n353), .ZN(G1347gat));
  NOR2_X1   g746(.A1(new_n703), .A2(new_n712), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n862), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(new_n863), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n951), .A2(G169gat), .A3(new_n304), .ZN(new_n952));
  AOI21_X1  g751(.A(G169gat), .B1(new_n951), .B2(new_n767), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n952), .A2(new_n953), .ZN(G1348gat));
  NAND2_X1  g753(.A1(new_n951), .A2(new_n698), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(G176gat), .ZN(G1349gat));
  OAI21_X1  g755(.A(new_n413), .B1(new_n950), .B2(new_n725), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n951), .A2(new_n786), .ZN(new_n958));
  OAI221_X1 g757(.A(new_n957), .B1(KEYINPUT125), .B2(KEYINPUT60), .C1(new_n958), .C2(new_n396), .ZN(new_n959));
  NAND2_X1  g758(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n959), .B(new_n960), .ZN(G1350gat));
  OAI22_X1  g760(.A1(new_n950), .A2(new_n728), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n962));
  NAND2_X1  g761(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n962), .B(new_n963), .ZN(G1351gat));
  AND4_X1   g763(.A1(new_n717), .A2(new_n931), .A3(new_n932), .A4(new_n948), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(new_n304), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n203), .B1(new_n966), .B2(KEYINPUT127), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n967), .B1(KEYINPUT127), .B2(new_n966), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n949), .A2(new_n577), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n969), .B(KEYINPUT126), .Z(new_n970));
  NAND3_X1  g769(.A1(new_n970), .A2(new_n203), .A3(new_n767), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n968), .A2(new_n971), .ZN(G1352gat));
  NOR3_X1   g771(.A1(new_n969), .A2(G204gat), .A3(new_n724), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT62), .ZN(new_n974));
  INV_X1    g773(.A(G204gat), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n965), .A2(new_n698), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(G1353gat));
  NAND3_X1  g776(.A1(new_n970), .A2(new_n382), .A3(new_n786), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n965), .A2(new_n786), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n979), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n979), .B2(G211gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(G1354gat));
  AOI21_X1  g781(.A(G218gat), .B1(new_n970), .B2(new_n727), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n728), .A2(new_n381), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n983), .B1(new_n965), .B2(new_n984), .ZN(G1355gat));
endmodule


