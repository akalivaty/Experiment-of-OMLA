//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n580, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT69), .Z(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND3_X1   g041(.A1(KEYINPUT71), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT3), .B1(KEYINPUT71), .B2(G2104), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n474), .A2(new_n476), .A3(G125), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n477), .A2(KEYINPUT70), .B1(G113), .B2(G2104), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n480), .A3(G125), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n472), .B1(new_n482), .B2(G2105), .ZN(G160));
  NAND2_X1  g058(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(new_n475), .ZN(new_n485));
  NAND3_X1  g060(.A1(KEYINPUT71), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(G2105), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n466), .B1(new_n485), .B2(new_n486), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n488), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n466), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n500), .A2(new_n474), .A3(new_n476), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n466), .A2(G138), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(new_n485), .B2(new_n486), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n504), .B2(new_n501), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT72), .B1(new_n508), .B2(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(new_n511), .A3(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(G543), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n513), .A2(new_n514), .A3(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G88), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n524), .A2(new_n508), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n517), .A2(new_n523), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n529), .A2(new_n530), .B1(new_n520), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  INV_X1    g108(.A(G89), .ZN(new_n534));
  OAI221_X1 g109(.A(new_n532), .B1(new_n515), .B2(new_n533), .C1(new_n534), .C2(new_n521), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(G168));
  NAND2_X1  g111(.A1(new_n522), .A2(G90), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n516), .A2(G52), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n508), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  NAND2_X1  g117(.A1(new_n522), .A2(G81), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n516), .A2(G43), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n508), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  AND2_X1   g128(.A1(G53), .A2(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n510), .B1(new_n511), .B2(G651), .ZN(new_n555));
  NOR3_X1   g130(.A1(new_n508), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n514), .B(new_n554), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n509), .A2(new_n512), .B1(KEYINPUT6), .B2(new_n508), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n560), .A2(KEYINPUT73), .A3(new_n554), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(KEYINPUT9), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n557), .A2(new_n558), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n522), .A2(G91), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT75), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G65), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n518), .A2(new_n571), .A3(new_n519), .ZN(new_n572));
  AND2_X1   g147(.A1(KEYINPUT5), .A2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(KEYINPUT5), .A2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT74), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n570), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  AND2_X1   g151(.A1(G78), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n562), .A2(new_n564), .A3(new_n565), .A4(new_n578), .ZN(G299));
  XNOR2_X1  g154(.A(new_n535), .B(KEYINPUT76), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G286));
  OAI21_X1  g156(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n582));
  INV_X1    g157(.A(G49), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  OAI221_X1 g159(.A(new_n582), .B1(new_n515), .B2(new_n583), .C1(new_n584), .C2(new_n521), .ZN(G288));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n521), .B2(new_n587), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n560), .A2(KEYINPUT77), .A3(G86), .A4(new_n520), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n560), .A2(G48), .A3(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n518), .B2(new_n519), .ZN(new_n593));
  AND2_X1   g168(.A1(G73), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n590), .A2(new_n596), .ZN(G305));
  XNOR2_X1  g172(.A(KEYINPUT79), .B(G85), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n522), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  XOR2_X1   g175(.A(KEYINPUT78), .B(G47), .Z(new_n601));
  OAI221_X1 g176(.A(new_n599), .B1(new_n508), .B2(new_n600), .C1(new_n515), .C2(new_n601), .ZN(G290));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NOR2_X1   g178(.A1(G301), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n522), .A2(G92), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n572), .A2(new_n575), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n611), .A2(G651), .B1(G54), .B2(new_n516), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT80), .Z(new_n614));
  AOI21_X1  g189(.A(new_n604), .B1(new_n614), .B2(new_n603), .ZN(G284));
  AOI21_X1  g190(.A(new_n604), .B1(new_n614), .B2(new_n603), .ZN(G321));
  NOR3_X1   g191(.A1(new_n580), .A2(KEYINPUT81), .A3(new_n603), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(G286), .B2(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(G299), .A2(new_n603), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(G297));
  AOI21_X1  g196(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n614), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n614), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n548), .ZN(G323));
  XOR2_X1   g202(.A(KEYINPUT82), .B(KEYINPUT11), .Z(new_n628));
  XNOR2_X1  g203(.A(G323), .B(new_n628), .ZN(G282));
  INV_X1    g204(.A(new_n471), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n479), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT83), .B(G2100), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n632), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n487), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n489), .A2(G123), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n638), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(G2096), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(G2096), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n635), .A2(new_n641), .A3(new_n642), .ZN(G156));
  XOR2_X1   g218(.A(KEYINPUT84), .B(KEYINPUT14), .Z(new_n644));
  XOR2_X1   g219(.A(KEYINPUT15), .B(G2435), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2438), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  AOI21_X1  g222(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n646), .B2(new_n647), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n649), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT85), .ZN(new_n662));
  NOR2_X1   g237(.A1(G2072), .A2(G2078), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n442), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n660), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(KEYINPUT17), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n665), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n660), .B(new_n661), .C1(new_n442), .C2(new_n663), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  NAND3_X1  g244(.A1(new_n666), .A2(new_n662), .A3(new_n660), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n678), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  AOI211_X1 g258(.A(new_n680), .B(new_n683), .C1(new_n675), .C2(new_n679), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G229));
  MUX2_X1   g265(.A(G24), .B(G290), .S(G16), .Z(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(G1986), .Z(new_n692));
  OAI21_X1  g267(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n693));
  INV_X1    g268(.A(G107), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n693), .B1(new_n694), .B2(G2105), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT87), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n487), .A2(G131), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n489), .A2(G119), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  MUX2_X1   g274(.A(G25), .B(new_n699), .S(G29), .Z(new_n700));
  XOR2_X1   g275(.A(KEYINPUT35), .B(G1991), .Z(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT89), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(KEYINPUT36), .ZN(new_n705));
  MUX2_X1   g280(.A(G6), .B(G305), .S(G16), .Z(new_n706));
  XOR2_X1   g281(.A(KEYINPUT32), .B(G1981), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G22), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G166), .B2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(G1971), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n709), .A2(G23), .ZN(new_n714));
  INV_X1    g289(.A(G288), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n709), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT33), .B(G1976), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT88), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n708), .A2(new_n713), .A3(new_n719), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n692), .B(new_n705), .C1(new_n720), .C2(KEYINPUT34), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(KEYINPUT34), .B2(new_n720), .ZN(new_n722));
  OR3_X1    g297(.A1(new_n722), .A2(new_n704), .A3(KEYINPUT36), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n704), .B2(KEYINPUT36), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT91), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT25), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n479), .A2(G127), .ZN(new_n728));
  INV_X1    g303(.A(G115), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n473), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n730), .A2(G2105), .B1(new_n487), .B2(G139), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(KEYINPUT92), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n732), .A2(KEYINPUT92), .ZN(new_n735));
  OAI21_X1  g310(.A(G29), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G33), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(G29), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G2072), .ZN(new_n739));
  INV_X1    g314(.A(G1341), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n548), .A2(new_n709), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n709), .B2(G19), .ZN(new_n742));
  NOR2_X1   g317(.A1(G171), .A2(new_n709), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G5), .B2(new_n709), .ZN(new_n744));
  INV_X1    g319(.A(G1961), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n740), .A2(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G28), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(KEYINPUT30), .ZN(new_n748));
  AOI21_X1  g323(.A(G29), .B1(new_n747), .B2(KEYINPUT30), .ZN(new_n749));
  OR2_X1    g324(.A1(KEYINPUT31), .A2(G11), .ZN(new_n750));
  NAND2_X1  g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n748), .A2(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G29), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n640), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(G26), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT28), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n489), .A2(G128), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT90), .ZN(new_n758));
  OAI21_X1  g333(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n759));
  INV_X1    g334(.A(G116), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(G2105), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n487), .B2(G140), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n756), .B1(new_n763), .B2(G29), .ZN(new_n764));
  INV_X1    g339(.A(G2067), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n754), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n753), .A2(G27), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G164), .B2(new_n753), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G2078), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(KEYINPUT95), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n739), .A2(new_n746), .A3(new_n766), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n753), .A2(G35), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT96), .Z(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n493), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT29), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2090), .ZN(new_n776));
  OAI221_X1 g351(.A(new_n776), .B1(KEYINPUT95), .B2(new_n769), .C1(new_n738), .C2(G2072), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n709), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT23), .ZN(new_n779));
  INV_X1    g354(.A(G299), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(new_n709), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1956), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n771), .A2(new_n777), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n709), .A2(G4), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n614), .B2(new_n709), .ZN(new_n785));
  INV_X1    g360(.A(G1348), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n709), .A2(G21), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G168), .B2(new_n709), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(G1966), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT94), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT24), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n753), .B1(new_n792), .B2(G34), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n792), .B2(G34), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G160), .B2(G29), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(G2084), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT93), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G29), .B2(G32), .ZN(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT26), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n801), .A2(new_n802), .B1(G105), .B2(new_n630), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n487), .A2(G141), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n489), .A2(G129), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G29), .ZN(new_n808));
  MUX2_X1   g383(.A(new_n797), .B(new_n798), .S(new_n808), .Z(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT27), .B(G1996), .ZN(new_n810));
  OAI22_X1  g385(.A1(new_n809), .A2(new_n810), .B1(new_n765), .B2(new_n764), .ZN(new_n811));
  AOI211_X1 g386(.A(new_n796), .B(new_n811), .C1(new_n810), .C2(new_n809), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n795), .A2(G2084), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n740), .A2(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n814));
  AOI211_X1 g389(.A(new_n813), .B(new_n814), .C1(G1966), .C2(new_n789), .ZN(new_n815));
  AND4_X1   g390(.A1(new_n787), .A2(new_n791), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n723), .A2(new_n724), .A3(new_n783), .A4(new_n816), .ZN(G150));
  INV_X1    g392(.A(G150), .ZN(G311));
  NAND2_X1  g393(.A1(new_n522), .A2(G93), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n516), .A2(G55), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n520), .A2(G67), .ZN(new_n821));
  NAND2_X1  g396(.A1(G80), .A2(G543), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G651), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n819), .A2(new_n820), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT97), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT97), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n819), .A2(new_n820), .A3(new_n827), .A4(new_n824), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n548), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n547), .A2(new_n825), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT38), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n614), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n835));
  AOI21_X1  g410(.A(G860), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT98), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n826), .A2(new_n828), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT37), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(G145));
  XNOR2_X1  g417(.A(new_n699), .B(new_n632), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n758), .A2(new_n762), .ZN(new_n845));
  OAI211_X1 g420(.A(KEYINPUT100), .B(new_n502), .C1(new_n504), .C2(new_n501), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n500), .B1(new_n467), .B2(new_n468), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT4), .ZN(new_n849));
  AOI21_X1  g424(.A(KEYINPUT100), .B1(new_n849), .B2(new_n502), .ZN(new_n850));
  OAI211_X1 g425(.A(KEYINPUT101), .B(new_n498), .C1(new_n847), .C2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n505), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n846), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT101), .B1(new_n855), .B2(new_n498), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n845), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n498), .B1(new_n847), .B2(new_n850), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(new_n763), .A3(new_n851), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n857), .A2(new_n807), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n807), .B1(new_n857), .B2(new_n861), .ZN(new_n864));
  OAI21_X1  g439(.A(KEYINPUT102), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n732), .B1(new_n865), .B2(KEYINPUT92), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n487), .A2(G142), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n489), .A2(G130), .ZN(new_n868));
  OR2_X1    g443(.A1(G106), .A2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n869), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n857), .A2(new_n861), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n806), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n862), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n734), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n866), .A2(new_n872), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n732), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n876), .B1(new_n874), .B2(new_n862), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT92), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n878), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n871), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n844), .B1(new_n879), .B2(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(G160), .B(KEYINPUT99), .Z(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n493), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n640), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n872), .B1(new_n866), .B2(new_n878), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n883), .A2(new_n884), .A3(new_n871), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n891), .A3(new_n843), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n886), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n886), .A2(KEYINPUT103), .A3(new_n889), .A4(new_n892), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n889), .B1(new_n886), .B2(new_n892), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(G37), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n897), .A2(KEYINPUT40), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT40), .B1(new_n897), .B2(new_n899), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(G395));
  NAND2_X1  g477(.A1(new_n839), .A2(new_n603), .ZN(new_n903));
  INV_X1    g478(.A(new_n831), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n625), .B(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n613), .A2(G299), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n780), .A2(new_n607), .A3(new_n612), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n906), .A3(new_n908), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n905), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n907), .A2(new_n908), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n914), .A2(new_n915), .B1(new_n905), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n915), .B2(new_n914), .ZN(new_n919));
  XNOR2_X1  g494(.A(G290), .B(G305), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n715), .B(G303), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n920), .B(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n922), .B(KEYINPUT42), .Z(new_n923));
  XNOR2_X1  g498(.A(new_n919), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n903), .B1(new_n924), .B2(new_n603), .ZN(G295));
  OAI21_X1  g500(.A(new_n903), .B1(new_n924), .B2(new_n603), .ZN(G331));
  NOR2_X1   g501(.A1(G286), .A2(G301), .ZN(new_n927));
  NOR2_X1   g502(.A1(G171), .A2(G168), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n831), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(new_n580), .B2(G171), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n904), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n917), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n831), .B(new_n930), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n912), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n922), .ZN(new_n937));
  AOI21_X1  g512(.A(G37), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n910), .A2(new_n939), .A3(new_n911), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n909), .A2(KEYINPUT107), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n934), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n937), .B1(new_n942), .B2(new_n933), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(KEYINPUT108), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n945));
  AOI211_X1 g520(.A(new_n945), .B(new_n937), .C1(new_n942), .C2(new_n933), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n938), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n933), .A2(new_n935), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT105), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n933), .A2(new_n935), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n953), .A3(new_n922), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT43), .B1(new_n954), .B2(new_n938), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT44), .B1(new_n949), .B2(new_n955), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n938), .B(new_n948), .C1(new_n944), .C2(new_n946), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n948), .B1(new_n954), .B2(new_n938), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n957), .B1(new_n958), .B2(KEYINPUT106), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n960));
  AOI211_X1 g535(.A(new_n960), .B(new_n948), .C1(new_n954), .C2(new_n938), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n956), .B1(new_n962), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g538(.A1(G303), .A2(G8), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT55), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n966));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n966), .B1(new_n858), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n848), .A2(KEYINPUT4), .B1(new_n969), .B2(new_n479), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n495), .A2(new_n497), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(G160), .B(G40), .C1(KEYINPUT50), .C2(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n968), .A2(new_n973), .A3(G2090), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n860), .A2(KEYINPUT45), .A3(new_n967), .A4(new_n851), .ZN(new_n975));
  NAND2_X1  g550(.A1(G160), .A2(G40), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n976), .B1(new_n977), .B2(new_n972), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n974), .B1(new_n979), .B2(new_n712), .ZN(new_n980));
  INV_X1    g555(.A(G8), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n965), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT112), .ZN(new_n983));
  INV_X1    g558(.A(G40), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n984), .B(new_n472), .C1(new_n482), .C2(G2105), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(new_n967), .A3(new_n858), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n715), .A2(G1976), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(G8), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT52), .ZN(new_n989));
  AOI21_X1  g564(.A(G1384), .B1(new_n855), .B2(new_n498), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n981), .B1(new_n990), .B2(new_n985), .ZN(new_n991));
  INV_X1    g566(.A(G1976), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT52), .B1(G288), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n987), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1981), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n590), .A2(new_n995), .A3(new_n596), .ZN(new_n996));
  NOR2_X1   g571(.A1(KEYINPUT110), .A2(G86), .ZN(new_n997));
  AND2_X1   g572(.A1(KEYINPUT110), .A2(G86), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n521), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n591), .A2(new_n595), .ZN(new_n1000));
  OAI21_X1  g575(.A(G1981), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n996), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT49), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(KEYINPUT111), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n991), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1003), .B1(new_n1002), .B2(KEYINPUT111), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n989), .B(new_n994), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n979), .A2(new_n712), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n976), .B1(new_n990), .B2(new_n966), .ZN(new_n1009));
  INV_X1    g584(.A(G2090), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1384), .B1(new_n498), .B2(new_n505), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT109), .B1(new_n1011), .B2(new_n966), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n972), .A2(new_n1013), .A3(KEYINPUT50), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(new_n1010), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n981), .B1(new_n1008), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n965), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1007), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1020), .B(new_n965), .C1(new_n980), .C2(new_n981), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n1022));
  INV_X1    g597(.A(G1966), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT45), .B1(new_n858), .B2(new_n967), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1011), .A2(KEYINPUT45), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n985), .A2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1022), .B(new_n1023), .C1(new_n1024), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G2084), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n858), .A2(new_n966), .A3(new_n967), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1015), .A2(new_n1028), .A3(new_n1029), .A4(new_n985), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n985), .B(new_n1025), .C1(new_n990), .C2(KEYINPUT45), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1022), .B1(new_n1032), .B2(new_n1023), .ZN(new_n1033));
  OAI211_X1 g608(.A(G8), .B(new_n580), .C1(new_n1031), .C2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n983), .A2(new_n1019), .A3(new_n1021), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT63), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1008), .A2(new_n1016), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G8), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n965), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n1019), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1019), .A2(new_n1041), .A3(new_n1042), .A4(KEYINPUT114), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1038), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1040), .A2(new_n1007), .A3(new_n965), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n992), .B(new_n715), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n996), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n991), .B2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT56), .B(G2072), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n975), .A2(new_n978), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n1054), .A2(KEYINPUT115), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(KEYINPUT115), .ZN(new_n1056));
  XOR2_X1   g631(.A(new_n1056), .B(KEYINPUT116), .Z(new_n1057));
  AND3_X1   g632(.A1(G299), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1057), .B1(G299), .B2(new_n1055), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1956), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n968), .B2(new_n973), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1053), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1058), .A2(new_n1059), .A3(KEYINPUT117), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n1065));
  NAND2_X1  g640(.A1(G299), .A2(new_n1055), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1057), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(G299), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1065), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1064), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1053), .A2(new_n1062), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n613), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1348), .B1(new_n1009), .B2(new_n1015), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n986), .A2(G2067), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1063), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1053), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT121), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1053), .A2(new_n1060), .A3(new_n1081), .A4(new_n1062), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT61), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NOR4_X1   g661(.A1(new_n1075), .A2(KEYINPUT60), .A3(new_n1076), .A4(new_n613), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1029), .A2(new_n985), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n786), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1076), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(new_n613), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1077), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1087), .B1(new_n1093), .B2(KEYINPUT60), .ZN(new_n1094));
  INV_X1    g669(.A(G1996), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n975), .A2(new_n978), .A3(new_n1095), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT58), .B(G1341), .Z(new_n1097));
  NAND2_X1  g672(.A1(new_n986), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT118), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n986), .A2(new_n1100), .A3(new_n1097), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1096), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n548), .A3(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n986), .A2(new_n1100), .A3(new_n1097), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1100), .B1(new_n986), .B2(new_n1097), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n547), .B1(new_n1107), .B2(new_n1096), .ZN(new_n1108));
  NOR2_X1   g683(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1104), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1086), .A2(new_n1094), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1060), .B1(new_n1053), .B2(new_n1062), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1084), .B1(new_n1063), .B2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(KEYINPUT120), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1078), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n983), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1116));
  OAI21_X1  g691(.A(G8), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1117));
  NOR2_X1   g692(.A1(G168), .A2(new_n981), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT51), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1124));
  OAI22_X1  g699(.A1(new_n1122), .A2(new_n1123), .B1(new_n1124), .B2(new_n1119), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n979), .B2(G2078), .ZN(new_n1127));
  XNOR2_X1  g702(.A(G301), .B(KEYINPUT54), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(new_n745), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n860), .A2(new_n967), .A3(new_n851), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n977), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1126), .A2(G2078), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1132), .A2(new_n985), .A3(new_n975), .A4(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1127), .A2(new_n1130), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1032), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1136), .A2(new_n1133), .B1(new_n1129), .B2(new_n745), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n1127), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1128), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1116), .A2(new_n1125), .A3(new_n1135), .A4(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1047), .B(new_n1051), .C1(new_n1115), .C2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT123), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1078), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1113), .B(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1086), .A2(new_n1094), .A3(new_n1110), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1124), .A2(new_n1119), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1121), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1148), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1139), .A2(new_n1135), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1147), .A2(new_n1116), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(new_n1047), .A4(new_n1051), .ZN(new_n1158));
  AOI21_X1  g733(.A(G301), .B1(new_n1137), .B2(new_n1127), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1116), .B(new_n1159), .C1(new_n1125), .C2(KEYINPUT62), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT124), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1153), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n1116), .A4(new_n1159), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1161), .B(new_n1165), .C1(new_n1162), .C2(new_n1153), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1142), .A2(new_n1158), .A3(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1132), .A2(new_n976), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n763), .B(new_n765), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n806), .B(new_n1095), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n699), .A2(new_n702), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n699), .A2(new_n702), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(G290), .B(G1986), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1168), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1167), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1174), .A2(new_n1168), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1168), .ZN(new_n1179));
  OR3_X1    g754(.A1(new_n1179), .A2(G1986), .A3(G290), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT48), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1178), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1182), .B1(new_n1181), .B2(new_n1180), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1173), .B(KEYINPUT125), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1171), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(G2067), .B2(new_n763), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1183), .B1(new_n1168), .B2(new_n1186), .ZN(new_n1187));
  OR3_X1    g762(.A1(new_n1179), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT46), .B1(new_n1179), .B2(G1996), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1169), .A2(new_n807), .ZN(new_n1190));
  AOI22_X1  g765(.A1(new_n1188), .A2(new_n1189), .B1(new_n1168), .B2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1191), .B(KEYINPUT47), .Z(new_n1192));
  NAND2_X1  g767(.A1(new_n1187), .A2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT126), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1177), .A2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g770(.A1(G227), .A2(new_n464), .ZN(new_n1197));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n1198));
  NOR2_X1   g772(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1200), .A2(new_n658), .ZN(new_n1201));
  NOR3_X1   g775(.A1(G229), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  OAI21_X1  g776(.A(new_n1202), .B1(new_n959), .B2(new_n961), .ZN(new_n1203));
  AOI21_X1  g777(.A(new_n1203), .B1(new_n897), .B2(new_n899), .ZN(G308));
  NAND2_X1  g778(.A1(new_n897), .A2(new_n899), .ZN(new_n1205));
  OAI211_X1 g779(.A(new_n1205), .B(new_n1202), .C1(new_n961), .C2(new_n959), .ZN(G225));
endmodule


