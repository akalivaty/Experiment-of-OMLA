//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n558, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G137), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n463), .A2(new_n470), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT68), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n478), .B1(new_n463), .B2(new_n470), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT69), .Z(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n466), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n483), .A2(new_n485), .B1(new_n464), .B2(G136), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n481), .A2(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G138), .B(new_n470), .C1(new_n461), .C2(new_n462), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(new_n470), .A3(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n490), .B1(new_n463), .B2(new_n492), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n491), .A2(new_n470), .A3(G138), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n471), .A2(new_n494), .A3(KEYINPUT70), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n489), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n500), .B1(new_n476), .B2(G126), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n496), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n497), .B1(new_n496), .B2(new_n501), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT72), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(G543), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(new_n509), .B1(KEYINPUT5), .B2(new_n505), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n505), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(new_n515), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n513), .A2(new_n521), .ZN(G166));
  NAND2_X1  g097(.A1(new_n506), .A2(new_n509), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT73), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n510), .A2(new_n528), .A3(G63), .A4(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n510), .A2(G89), .A3(new_n518), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n534), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n516), .A2(G51), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n530), .A2(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  AOI22_X1  g114(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n512), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n516), .A2(G52), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n519), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(KEYINPUT74), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NOR3_X1   g121(.A1(new_n541), .A2(new_n544), .A3(KEYINPUT74), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  AOI22_X1  g124(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n512), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n516), .A2(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n519), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT75), .ZN(G188));
  AOI22_X1  g136(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n562), .A2(new_n512), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n519), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G91), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n516), .A2(G53), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n564), .A2(new_n566), .A3(new_n568), .ZN(G299));
  INV_X1    g144(.A(G166), .ZN(G303));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT76), .B1(new_n519), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n510), .A2(new_n573), .A3(G87), .A4(new_n518), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n510), .A2(G74), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(G49), .B2(new_n516), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(new_n516), .A2(G48), .ZN(new_n579));
  INV_X1    g154(.A(G86), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n519), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n510), .A2(G61), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n512), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n516), .A2(G47), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n519), .B2(new_n591), .ZN(new_n592));
  OR3_X1    g167(.A1(new_n589), .A2(new_n592), .A3(KEYINPUT77), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT77), .B1(new_n589), .B2(new_n592), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G290));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NOR2_X1   g171(.A1(G301), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n565), .A2(G92), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n525), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n516), .A2(G54), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n597), .B1(new_n596), .B2(new_n607), .ZN(G284));
  AOI21_X1  g183(.A(new_n597), .B1(new_n596), .B2(new_n607), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  AND3_X1   g185(.A1(new_n564), .A2(new_n566), .A3(new_n568), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  XOR2_X1   g187(.A(G280), .B(KEYINPUT78), .Z(G297));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n607), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n471), .A2(new_n467), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n480), .A2(G123), .ZN(new_n624));
  INV_X1    g199(.A(G111), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n625), .A2(KEYINPUT79), .A3(G2105), .ZN(new_n626));
  AOI21_X1  g201(.A(KEYINPUT79), .B1(new_n625), .B2(G2105), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI22_X1  g204(.A1(new_n464), .A2(G135), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n623), .A2(G2100), .B1(new_n631), .B2(G2096), .ZN(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n622), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n632), .B(new_n634), .C1(G2096), .C2(new_n631), .ZN(G156));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(new_n640), .A3(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n645), .A2(new_n648), .ZN(new_n650));
  AND3_X1   g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(G401));
  INV_X1    g226(.A(KEYINPUT18), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n652), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(new_n633), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n655), .B2(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(G2096), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1961), .B(G1966), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT81), .B(KEYINPUT20), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n669), .B(new_n670), .Z(new_n671));
  AND2_X1   g246(.A1(new_n666), .A2(new_n667), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT82), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n665), .A2(new_n672), .A3(new_n668), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT83), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1981), .B(G1986), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  NAND3_X1  g258(.A1(new_n575), .A2(new_n577), .A3(KEYINPUT85), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(KEYINPUT85), .B1(new_n575), .B2(new_n577), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G16), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G16), .B2(G23), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT33), .B(G1976), .Z(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n691), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G22), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G1971), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(G6), .A2(G16), .ZN(new_n699));
  INV_X1    g274(.A(G305), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(G16), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT32), .B(G1981), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n692), .A2(new_n693), .A3(new_n698), .A4(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(KEYINPUT34), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(KEYINPUT34), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n694), .A2(G24), .ZN(new_n707));
  INV_X1    g282(.A(G290), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n694), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(G1986), .Z(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G25), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n480), .A2(G119), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n464), .A2(G131), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n470), .A2(G107), .ZN(new_n715));
  OAI21_X1  g290(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n713), .B(new_n714), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT84), .Z(new_n718));
  OAI21_X1  g293(.A(new_n712), .B1(new_n718), .B2(new_n711), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT35), .B(G1991), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n719), .B(new_n720), .Z(new_n721));
  NAND4_X1  g296(.A1(new_n705), .A2(new_n706), .A3(new_n710), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT36), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n694), .A2(G21), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G168), .B2(new_n694), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT90), .Z(new_n726));
  INV_X1    g301(.A(G1966), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n694), .A2(G5), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G171), .B2(new_n694), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n728), .B(new_n729), .C1(G1961), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n711), .A2(G33), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(new_n470), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT87), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT25), .Z(new_n738));
  AOI211_X1 g313(.A(new_n735), .B(new_n738), .C1(G139), .C2(new_n464), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n733), .B1(new_n739), .B2(new_n711), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(G2072), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(G2072), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT31), .B(G11), .Z(new_n743));
  NOR2_X1   g318(.A1(new_n631), .A2(new_n711), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT30), .B(G28), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n743), .B(new_n744), .C1(new_n711), .C2(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n741), .A2(new_n742), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G1348), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n607), .A2(new_n694), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G4), .B2(new_n694), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n747), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n480), .A2(G129), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n467), .A2(G105), .ZN(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT26), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n753), .B(new_n755), .C1(G141), .C2(new_n464), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  MUX2_X1   g332(.A(G32), .B(new_n757), .S(G29), .Z(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT27), .B(G1996), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G16), .A2(G19), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n555), .B2(G16), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(G1341), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n765), .B2(G34), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G34), .B2(new_n765), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G160), .B2(new_n711), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT89), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n769), .A2(G2084), .B1(G1341), .B2(new_n762), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n751), .A2(new_n760), .A3(new_n763), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n711), .A2(G35), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G162), .B2(new_n711), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT29), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2090), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G1961), .B2(new_n731), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n771), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n769), .A2(G2084), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT91), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n711), .A2(G26), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT28), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n480), .A2(G128), .ZN(new_n782));
  OAI21_X1  g357(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n783));
  INV_X1    g358(.A(G116), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(G2105), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n464), .B2(G140), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G29), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n788), .A2(KEYINPUT86), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(KEYINPUT86), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n781), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G2067), .ZN(new_n792));
  NOR2_X1   g367(.A1(G164), .A2(new_n711), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G27), .B2(new_n711), .ZN(new_n794));
  INV_X1    g369(.A(G2078), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n750), .B2(new_n748), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n694), .A2(G20), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT23), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n611), .B2(new_n694), .ZN(new_n800));
  INV_X1    g375(.A(G1956), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n795), .B2(new_n794), .ZN(new_n803));
  NOR4_X1   g378(.A1(new_n779), .A2(new_n792), .A3(new_n797), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n723), .A2(new_n732), .A3(new_n777), .A4(new_n804), .ZN(G150));
  INV_X1    g380(.A(G150), .ZN(G311));
  NAND2_X1  g381(.A1(new_n607), .A2(G559), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT38), .ZN(new_n808));
  OAI21_X1  g383(.A(KEYINPUT93), .B1(new_n555), .B2(KEYINPUT92), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT92), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT93), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n810), .B(new_n811), .C1(new_n551), .C2(new_n554), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n555), .A2(KEYINPUT92), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(new_n512), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n516), .A2(G55), .ZN(new_n817));
  INV_X1    g392(.A(G93), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n519), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n813), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n809), .A2(new_n820), .A3(new_n814), .A4(new_n812), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n808), .B(new_n824), .Z(new_n825));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n826));
  AOI21_X1  g401(.A(G860), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT94), .Z(new_n829));
  OAI21_X1  g404(.A(G860), .B1(new_n816), .B2(new_n819), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(G145));
  XNOR2_X1  g407(.A(new_n631), .B(G160), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G162), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n757), .B(new_n787), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT95), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n496), .A2(new_n501), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n836), .B1(new_n496), .B2(new_n501), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n835), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n739), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n464), .A2(G142), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(KEYINPUT96), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(KEYINPUT96), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(G118), .B2(new_n470), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n843), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n480), .B2(G130), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(new_n621), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n717), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n842), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n842), .A2(new_n852), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n854), .B1(KEYINPUT97), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n842), .A2(KEYINPUT97), .A3(new_n852), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n834), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n834), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n855), .A2(new_n859), .A3(new_n853), .ZN(new_n860));
  INV_X1    g435(.A(G37), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n858), .A2(KEYINPUT40), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT40), .B1(new_n858), .B2(new_n862), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(G395));
  OAI21_X1  g440(.A(new_n596), .B1(new_n816), .B2(new_n819), .ZN(new_n866));
  XNOR2_X1  g441(.A(G166), .B(KEYINPUT100), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n687), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n687), .A2(new_n867), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n708), .A2(G305), .ZN(new_n871));
  NAND2_X1  g446(.A1(G290), .A2(new_n700), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n870), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n874), .B1(KEYINPUT101), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(KEYINPUT101), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n824), .B(new_n616), .Z(new_n879));
  NAND2_X1  g454(.A1(G299), .A2(KEYINPUT98), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT10), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n598), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n564), .A2(new_n883), .A3(new_n568), .A4(new_n566), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n880), .A2(new_n882), .A3(new_n605), .A4(new_n884), .ZN(new_n885));
  OAI211_X1 g460(.A(KEYINPUT98), .B(G299), .C1(new_n599), .C2(new_n606), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT41), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n879), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n887), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n893), .A2(KEYINPUT99), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n885), .A2(KEYINPUT99), .A3(new_n886), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n892), .B1(new_n879), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n878), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n866), .B1(new_n898), .B2(new_n596), .ZN(G295));
  OAI21_X1  g474(.A(new_n866), .B1(new_n898), .B2(new_n596), .ZN(G331));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n901));
  OAI21_X1  g476(.A(G286), .B1(new_n546), .B2(new_n547), .ZN(new_n902));
  INV_X1    g477(.A(new_n547), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(G168), .A3(new_n545), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n824), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n822), .A2(new_n902), .A3(new_n823), .A4(new_n904), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(KEYINPUT103), .A3(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n907), .A2(KEYINPUT103), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n893), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n889), .A2(new_n890), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n912), .B1(new_n907), .B2(new_n906), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n871), .A2(new_n872), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n870), .B(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n911), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n887), .B1(new_n908), .B2(new_n909), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n874), .B1(new_n918), .B2(new_n913), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n917), .A2(new_n919), .A3(new_n920), .A4(new_n861), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n918), .A2(new_n874), .A3(new_n913), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n891), .A2(new_n908), .A3(new_n909), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n906), .B(new_n907), .C1(new_n894), .C2(new_n895), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n916), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n922), .A2(new_n925), .A3(G37), .ZN(new_n926));
  OAI211_X1 g501(.A(KEYINPUT44), .B(new_n921), .C1(new_n926), .C2(new_n920), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n917), .A2(new_n861), .A3(new_n919), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n932));
  INV_X1    g507(.A(new_n925), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n933), .A2(new_n917), .A3(new_n920), .A4(new_n861), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n930), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n901), .B1(new_n928), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n934), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n929), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(KEYINPUT104), .A3(new_n927), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(G397));
  NOR3_X1   g515(.A1(new_n838), .A2(G1384), .A3(new_n839), .ZN(new_n941));
  XOR2_X1   g516(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n474), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n944), .A2(G40), .A3(new_n468), .A4(new_n465), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n941), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G2067), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n787), .B(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n757), .B(G1996), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT107), .Z(new_n952));
  INV_X1    g527(.A(new_n718), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n953), .A2(new_n720), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(G2067), .B2(new_n787), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n946), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n717), .B(new_n720), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n946), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n952), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT125), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n952), .A2(KEYINPUT125), .A3(new_n959), .ZN(new_n963));
  INV_X1    g538(.A(G1986), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n946), .A2(new_n964), .A3(new_n708), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT48), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n946), .B1(new_n949), .B2(new_n757), .ZN(new_n968));
  INV_X1    g543(.A(G1996), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n946), .A2(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n970), .A2(KEYINPUT46), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(KEYINPUT46), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT124), .B(KEYINPUT47), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n957), .A2(new_n967), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT126), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n957), .A2(new_n967), .A3(KEYINPUT126), .A4(new_n975), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n496), .A2(new_n501), .ZN(new_n981));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(new_n945), .ZN(new_n984));
  XNOR2_X1  g559(.A(KEYINPUT110), .B(G8), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1981), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n582), .A2(new_n586), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n512), .B1(new_n583), .B2(new_n584), .ZN(new_n989));
  OAI21_X1  g564(.A(G1981), .B1(new_n581), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n990), .A3(KEYINPUT111), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT49), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n993));
  NAND3_X1  g568(.A1(G305), .A2(new_n993), .A3(G1981), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n991), .A2(new_n994), .A3(KEYINPUT112), .A4(new_n992), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n992), .B1(new_n991), .B2(new_n994), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n1000), .A2(new_n985), .A3(new_n984), .ZN(new_n1001));
  AOI211_X1 g576(.A(G1976), .B(G288), .C1(new_n999), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n988), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n986), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n981), .A2(KEYINPUT71), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n496), .A2(new_n501), .A3(new_n497), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1384), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(new_n943), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n981), .A2(KEYINPUT95), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1010), .A2(KEYINPUT45), .A3(new_n982), .A4(new_n837), .ZN(new_n1011));
  INV_X1    g586(.A(G40), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n469), .A2(new_n474), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1005), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n982), .B1(new_n502), .B2(new_n503), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n942), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1017), .A2(KEYINPUT108), .A3(new_n1013), .A4(new_n1011), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n697), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1015), .A2(KEYINPUT109), .A3(new_n697), .A4(new_n1018), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1384), .B1(new_n496), .B2(new_n501), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n945), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n1008), .B2(new_n1024), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(G2090), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1021), .A2(new_n1022), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G303), .A2(G8), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT55), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(G8), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n999), .A2(new_n1001), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT85), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G288), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(G1976), .A3(new_n684), .ZN(new_n1036));
  INV_X1    g611(.A(G1976), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(G288), .B2(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1036), .A2(new_n986), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(new_n1036), .B2(new_n986), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1033), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1004), .B1(new_n1032), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n985), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT119), .B1(G286), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n1047), .B(new_n985), .C1(new_n530), .C2(new_n537), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1013), .B1(new_n983), .B2(KEYINPUT50), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(KEYINPUT50), .B2(new_n1016), .ZN(new_n1051));
  INV_X1    g626(.A(G2084), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n982), .B(new_n943), .C1(new_n502), .C2(new_n503), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n945), .B1(new_n983), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1051), .A2(new_n1052), .B1(new_n727), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G8), .ZN(new_n1058));
  OAI211_X1 g633(.A(KEYINPUT51), .B(new_n1049), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1056), .A2(new_n727), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1052), .B(new_n1025), .C1(new_n1008), .C2(new_n1024), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n985), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1049), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1060), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1059), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(new_n1064), .ZN(new_n1069));
  AOI211_X1 g644(.A(KEYINPUT120), .B(new_n1049), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT62), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT53), .B1(new_n1073), .B2(new_n795), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1026), .A2(KEYINPUT116), .ZN(new_n1075));
  INV_X1    g650(.A(G1961), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1077), .B(new_n1025), .C1(new_n1008), .C2(new_n1024), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1053), .A2(new_n1055), .A3(KEYINPUT53), .A4(new_n795), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(G171), .B1(new_n1074), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT120), .B1(new_n1057), .B2(new_n1049), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1068), .A2(new_n1067), .A3(new_n1064), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n1065), .A4(new_n1059), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1072), .A2(new_n1083), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n945), .B1(new_n983), .B2(KEYINPUT50), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1016), .B2(KEYINPUT50), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1091), .A2(G2090), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n985), .B1(new_n1019), .B2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1033), .B(new_n1042), .C1(new_n1093), .C2(new_n1031), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1027), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n1020), .B2(new_n1019), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1058), .B1(new_n1096), .B2(new_n1022), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1094), .B1(new_n1031), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1044), .B1(new_n1089), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1019), .A2(new_n1092), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n1045), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1043), .B1(new_n1101), .B2(new_n1030), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1057), .A2(G286), .A3(new_n985), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1032), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1103), .A2(KEYINPUT63), .A3(new_n1033), .A4(new_n1042), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1030), .A2(KEYINPUT113), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1107), .B1(new_n1097), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1028), .A2(G8), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(KEYINPUT113), .A3(new_n1030), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1106), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1114));
  OAI211_X1 g689(.A(KEYINPUT53), .B(new_n795), .C1(new_n941), .C2(new_n943), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(new_n1014), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1078), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1016), .A2(KEYINPUT50), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1077), .B1(new_n1118), .B2(new_n1025), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1116), .B1(new_n1120), .B2(new_n1076), .ZN(new_n1121));
  AOI21_X1  g696(.A(G2078), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1121), .B(G301), .C1(KEYINPUT53), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1082), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1114), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1121), .B(new_n1127), .C1(KEYINPUT53), .C2(new_n1122), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1116), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n1079), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT122), .B1(new_n1074), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1131), .A3(G171), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1074), .A2(new_n1081), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1133), .B1(new_n1134), .B2(G301), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n611), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1137), .ZN(new_n1140));
  NAND2_X1  g715(.A1(G299), .A2(new_n1140), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1138), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1139), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1091), .A2(new_n801), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT56), .B(G2072), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1017), .A2(new_n1013), .A3(new_n1011), .A4(new_n1146), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1075), .A2(new_n748), .A3(new_n1078), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n984), .A2(new_n947), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT115), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(G299), .B(new_n1137), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1145), .A2(new_n1147), .A3(new_n1154), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1155), .A2(new_n607), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1149), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1153), .A2(KEYINPUT60), .A3(new_n607), .ZN(new_n1158));
  OAI211_X1 g733(.A(KEYINPUT61), .B(new_n1155), .C1(new_n1144), .C2(new_n1148), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n607), .A2(KEYINPUT60), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n607), .A2(KEYINPUT60), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1150), .A2(new_n1152), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1158), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1145), .A2(new_n1147), .A3(new_n1154), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1154), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1017), .A2(new_n969), .A3(new_n1013), .A4(new_n1011), .ZN(new_n1167));
  XOR2_X1   g742(.A(KEYINPUT58), .B(G1341), .Z(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n983), .B2(new_n945), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1170), .A2(new_n555), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1171), .B1(new_n1170), .B2(new_n555), .ZN(new_n1173));
  OAI22_X1  g748(.A1(new_n1166), .A2(KEYINPUT61), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1157), .B1(new_n1163), .B2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1126), .A2(new_n1136), .A3(new_n1098), .A4(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1099), .A2(new_n1113), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n946), .A2(G1986), .A3(G290), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n965), .A2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT106), .Z(new_n1180));
  NOR2_X1   g755(.A1(new_n960), .A2(new_n1180), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1177), .A2(KEYINPUT123), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT123), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n980), .B1(new_n1182), .B2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g759(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1186));
  OR2_X1    g760(.A1(G229), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g761(.A(new_n1187), .B1(new_n858), .B2(new_n862), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n1188), .A2(new_n937), .ZN(G225));
  INV_X1    g763(.A(G225), .ZN(G308));
endmodule


