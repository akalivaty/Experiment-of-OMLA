//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n558, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n634, new_n637, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G236), .A3(G238), .A4(G235), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n453), .A2(G567), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G101), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT68), .A3(G101), .ZN(new_n476));
  OR2_X1    g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n473), .A2(new_n476), .B1(new_n479), .B2(G137), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n468), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n479), .A2(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT70), .Z(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(new_n470), .B2(G112), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT69), .B1(new_n464), .B2(new_n470), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT3), .B(G2104), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n489), .A2(new_n490), .A3(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(G124), .B2(new_n492), .ZN(G162));
  NAND2_X1  g068(.A1(new_n475), .A2(G102), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(new_n474), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n489), .B2(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n494), .B1(new_n497), .B2(new_n470), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n470), .C1(new_n462), .C2(new_n463), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n489), .A2(KEYINPUT4), .A3(G138), .A4(new_n470), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n498), .A2(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  AND2_X1   g086(.A1(G50), .A2(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n510), .A2(G651), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT71), .B1(new_n518), .B2(new_n508), .ZN(new_n519));
  OR2_X1    g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n522), .A2(new_n511), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n513), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n531));
  AND2_X1   g106(.A1(G63), .A2(G651), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n530), .A2(new_n531), .B1(new_n522), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n518), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n511), .A2(KEYINPUT72), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n535), .A2(new_n536), .A3(G543), .ZN(new_n537));
  INV_X1    g112(.A(G51), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  OAI221_X1 g114(.A(new_n533), .B1(new_n537), .B2(new_n538), .C1(new_n525), .C2(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  INV_X1    g116(.A(new_n525), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G90), .ZN(new_n543));
  INV_X1    g118(.A(new_n537), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G52), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n514), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n543), .A2(new_n545), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(new_n542), .A2(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n544), .A2(G43), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n514), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT73), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  AND2_X1   g136(.A1(KEYINPUT74), .A2(G53), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n535), .A2(new_n536), .A3(G543), .A4(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n508), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n525), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G299));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n574));
  AND3_X1   g149(.A1(new_n519), .A2(G88), .A3(new_n524), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n510), .A2(G651), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n511), .A2(new_n512), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n574), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n513), .B(KEYINPUT75), .C1(new_n526), .C2(new_n525), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(G303));
  NAND2_X1  g156(.A1(new_n542), .A2(G87), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n535), .A2(new_n536), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  INV_X1    g160(.A(G49), .ZN(new_n586));
  INV_X1    g161(.A(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n584), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n585), .B1(new_n584), .B2(new_n588), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n582), .B(new_n583), .C1(new_n589), .C2(new_n590), .ZN(G288));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n520), .B2(new_n521), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n593), .B2(new_n594), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT78), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n519), .A2(G86), .A3(new_n524), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n511), .A2(G48), .A3(G543), .ZN(new_n602));
  AND2_X1   g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n604), .B(G651), .C1(new_n596), .C2(new_n598), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n600), .A2(new_n603), .A3(new_n605), .ZN(G305));
  INV_X1    g181(.A(G85), .ZN(new_n607));
  INV_X1    g182(.A(G47), .ZN(new_n608));
  OAI22_X1  g183(.A1(new_n525), .A2(new_n607), .B1(new_n537), .B2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT80), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G72), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G60), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n508), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n514), .B1(new_n614), .B2(KEYINPUT79), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(KEYINPUT79), .B2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n611), .A2(new_n616), .ZN(G290));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NOR2_X1   g193(.A1(G301), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n519), .A2(G92), .A3(new_n524), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT10), .Z(new_n621));
  AOI22_X1  g196(.A1(new_n522), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(new_n514), .ZN(new_n623));
  INV_X1    g198(.A(G54), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n624), .B1(new_n537), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n625), .B2(new_n537), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n621), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT82), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n619), .B1(new_n630), .B2(new_n618), .ZN(G284));
  AOI21_X1  g206(.A(new_n619), .B1(new_n630), .B2(new_n618), .ZN(G321));
  NAND2_X1  g207(.A1(G286), .A2(G868), .ZN(new_n633));
  AOI22_X1  g208(.A1(G299), .A2(new_n618), .B1(KEYINPUT83), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(KEYINPUT83), .B2(new_n633), .ZN(G297));
  OAI21_X1  g210(.A(new_n634), .B1(KEYINPUT83), .B2(new_n633), .ZN(G280));
  INV_X1    g211(.A(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n630), .B1(new_n637), .B2(G860), .ZN(G148));
  NAND2_X1  g213(.A1(new_n554), .A2(new_n618), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n629), .A2(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(new_n618), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g217(.A1(new_n489), .A2(new_n475), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  INV_X1    g220(.A(G2100), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n492), .A2(G123), .ZN(new_n648));
  OAI21_X1  g223(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(KEYINPUT84), .ZN(new_n650));
  INV_X1    g225(.A(G111), .ZN(new_n651));
  AOI22_X1  g226(.A1(new_n649), .A2(KEYINPUT84), .B1(new_n651), .B2(G2105), .ZN(new_n652));
  AOI22_X1  g227(.A1(new_n650), .A2(new_n652), .B1(new_n479), .B2(G135), .ZN(new_n653));
  AND2_X1   g228(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n655), .A2(G2096), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n645), .A2(new_n646), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(G2096), .ZN(new_n658));
  NAND4_X1  g233(.A1(new_n647), .A2(new_n656), .A3(new_n657), .A4(new_n658), .ZN(G156));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT85), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2427), .B(G2438), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2430), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT15), .B(G2435), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(new_n671), .A3(KEYINPUT14), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n666), .A2(new_n673), .ZN(new_n675));
  AND3_X1   g250(.A1(new_n674), .A2(G14), .A3(new_n675), .ZN(G401));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n681));
  AOI21_X1  g256(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n680), .A2(KEYINPUT17), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  MUX2_X1   g260(.A(new_n682), .B(new_n677), .S(new_n685), .Z(new_n686));
  XNOR2_X1  g261(.A(G2096), .B(G2100), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1971), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1961), .B(G1966), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n690), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n690), .A2(new_n693), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT20), .Z(new_n697));
  AOI211_X1 g272(.A(new_n695), .B(new_n697), .C1(new_n690), .C2(new_n694), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  INV_X1    g274(.A(G1981), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n698), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1991), .B(G1996), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT88), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT87), .B(G1986), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(G229));
  INV_X1    g284(.A(KEYINPUT93), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G25), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n492), .A2(G119), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(G95), .A2(G2105), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT90), .ZN(new_n717));
  INV_X1    g292(.A(G107), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n474), .B1(new_n718), .B2(G2105), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n717), .A2(new_n719), .B1(G131), .B2(new_n479), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n712), .B1(new_n721), .B2(new_n711), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G24), .ZN(new_n726));
  INV_X1    g301(.A(G290), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(KEYINPUT91), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(G16), .B1(new_n727), .B2(KEYINPUT91), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n726), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n710), .B(new_n724), .C1(new_n731), .C2(G1986), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G1986), .B2(new_n731), .ZN(new_n733));
  MUX2_X1   g308(.A(G23), .B(G288), .S(G16), .Z(new_n734));
  XOR2_X1   g309(.A(KEYINPUT33), .B(G1976), .Z(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n725), .A2(G22), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G166), .B2(new_n725), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1971), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n725), .A2(G6), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G305), .B2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT32), .B(G1981), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n742), .A2(new_n744), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n734), .A2(new_n735), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n740), .A2(new_n746), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n749), .B2(KEYINPUT34), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n749), .A2(new_n750), .A3(KEYINPUT34), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n733), .B1(KEYINPUT34), .B2(new_n749), .C1(new_n751), .C2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT36), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT31), .B(G11), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT97), .B(G28), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(KEYINPUT30), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(new_n711), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n758), .A2(KEYINPUT30), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n654), .A2(G29), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(KEYINPUT96), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(KEYINPUT96), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n725), .A2(G5), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G171), .B2(new_n725), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n765), .B1(G1961), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n725), .A2(G21), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G168), .B2(new_n725), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT95), .B(G1966), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT98), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n711), .A2(G35), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G162), .B2(new_n711), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT29), .Z(new_n777));
  INV_X1    g352(.A(G2090), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n725), .A2(G20), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT23), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n572), .B2(new_n725), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1956), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n774), .B1(KEYINPUT99), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n711), .A2(G27), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G164), .B2(new_n711), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(G2078), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n711), .A2(G32), .ZN(new_n789));
  NAND3_X1  g364(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT26), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n479), .A2(G141), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n475), .A2(G105), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G129), .B2(new_n492), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n789), .B1(new_n795), .B2(new_n711), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT27), .B(G1996), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n788), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT94), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT25), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n479), .A2(G139), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n489), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n802), .B(new_n803), .C1(new_n470), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(G29), .ZN(new_n806));
  INV_X1    g381(.A(G33), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(G29), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G2072), .ZN(new_n809));
  INV_X1    g384(.A(G2072), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n806), .B(new_n810), .C1(G29), .C2(new_n807), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n711), .B1(KEYINPUT24), .B2(G34), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(KEYINPUT24), .B2(G34), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n481), .B2(G29), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G2084), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n796), .A2(new_n798), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n809), .A2(new_n811), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  AOI211_X1 g392(.A(new_n799), .B(new_n817), .C1(new_n778), .C2(new_n777), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n784), .A2(KEYINPUT99), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n711), .A2(G26), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT28), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n479), .A2(G140), .ZN(new_n822));
  NOR2_X1   g397(.A1(G104), .A2(G2105), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(new_n470), .B2(G116), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G128), .B2(new_n492), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n821), .B1(new_n826), .B2(new_n711), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G2067), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n725), .A2(G19), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n555), .B2(new_n725), .ZN(new_n830));
  OAI22_X1  g405(.A1(G1341), .A2(new_n830), .B1(new_n767), .B2(G1961), .ZN(new_n831));
  AOI211_X1 g406(.A(new_n828), .B(new_n831), .C1(G1341), .C2(new_n830), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n818), .A2(new_n819), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n725), .A2(G4), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n630), .B2(new_n725), .ZN(new_n835));
  INV_X1    g410(.A(G1348), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n785), .A2(new_n833), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n754), .B2(new_n755), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n756), .A2(new_n839), .A3(KEYINPUT100), .ZN(new_n840));
  AOI21_X1  g415(.A(KEYINPUT100), .B1(new_n756), .B2(new_n839), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(G311));
  NAND2_X1  g417(.A1(new_n756), .A2(new_n839), .ZN(G150));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  INV_X1    g419(.A(G67), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n508), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT101), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n514), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n544), .A2(G55), .ZN(new_n850));
  XNOR2_X1  g425(.A(KEYINPUT102), .B(G93), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n849), .B(new_n850), .C1(new_n525), .C2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n555), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT38), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n637), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n857));
  AOI21_X1  g432(.A(G860), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n852), .A2(G860), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT103), .Z(G145));
  INV_X1    g438(.A(KEYINPUT107), .ZN(new_n864));
  INV_X1    g439(.A(G37), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT4), .B1(new_n479), .B2(G138), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n499), .A2(new_n500), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G126), .ZN(new_n870));
  OAI22_X1  g445(.A1(new_n464), .A2(new_n870), .B1(new_n495), .B2(new_n474), .ZN(new_n871));
  AOI22_X1  g446(.A1(new_n871), .A2(G2105), .B1(G102), .B2(new_n475), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT104), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n826), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n795), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(new_n805), .Z(new_n877));
  NAND2_X1  g452(.A1(new_n715), .A2(new_n720), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n644), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n881));
  INV_X1    g456(.A(G118), .ZN(new_n882));
  AOI22_X1  g457(.A1(new_n880), .A2(new_n881), .B1(new_n882), .B2(G2105), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n881), .B2(new_n880), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n479), .A2(G142), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(G130), .B2(new_n492), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n879), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n877), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(G162), .B(G160), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n654), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n877), .A2(new_n888), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n865), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n889), .A2(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n877), .A2(new_n888), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n893), .A2(new_n896), .A3(new_n889), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n864), .B(new_n895), .C1(new_n901), .C2(new_n891), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n891), .B1(new_n899), .B2(new_n900), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT107), .B1(new_n903), .B2(new_n894), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n902), .A2(KEYINPUT40), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT40), .B1(new_n902), .B2(new_n904), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(G395));
  XNOR2_X1  g482(.A(G290), .B(G166), .ZN(new_n908));
  XOR2_X1   g483(.A(G288), .B(G305), .Z(new_n909));
  XOR2_X1   g484(.A(new_n908), .B(new_n909), .Z(new_n910));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n910), .B1(KEYINPUT109), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n852), .B(new_n554), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n640), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n853), .B1(new_n629), .B2(G559), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n918));
  INV_X1    g493(.A(new_n628), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(new_n919), .B2(G299), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n628), .A2(KEYINPUT108), .A3(new_n572), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(G299), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT41), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n923), .A2(KEYINPUT41), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n917), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n911), .A2(KEYINPUT109), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n915), .A2(new_n916), .A3(new_n923), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n928), .B1(new_n926), .B2(new_n929), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n913), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n932), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n934), .A2(new_n930), .A3(new_n912), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(G868), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n852), .A2(new_n618), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n618), .B1(new_n933), .B2(new_n935), .ZN(new_n941));
  INV_X1    g516(.A(new_n939), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT110), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(G295));
  NAND2_X1  g519(.A1(new_n937), .A2(new_n939), .ZN(G331));
  XNOR2_X1  g520(.A(KEYINPUT113), .B(KEYINPUT44), .ZN(new_n946));
  AOI21_X1  g521(.A(G286), .B1(G171), .B2(KEYINPUT112), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n914), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n914), .A2(new_n947), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(G171), .A2(KEYINPUT112), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n951), .B1(new_n948), .B2(new_n949), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n923), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n925), .A2(new_n953), .A3(new_n924), .A4(new_n954), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n910), .ZN(new_n959));
  INV_X1    g534(.A(new_n910), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(new_n956), .A3(new_n957), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n865), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n959), .A2(new_n961), .A3(new_n964), .A4(new_n865), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n946), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n946), .ZN(new_n969));
  AOI211_X1 g544(.A(KEYINPUT111), .B(new_n969), .C1(new_n963), .C2(new_n965), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n968), .A2(new_n970), .ZN(G397));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n874), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n468), .A2(new_n480), .A3(G40), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n973), .B1(new_n498), .B2(new_n503), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n974), .A2(new_n977), .A3(new_n778), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n874), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n975), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(G1971), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(G8), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G8), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n981), .ZN(new_n985));
  INV_X1    g560(.A(G1971), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT104), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT104), .B1(new_n501), .B2(new_n502), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n988), .A2(new_n989), .A3(new_n498), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT50), .B1(new_n990), .B2(G1384), .ZN(new_n991));
  INV_X1    g566(.A(new_n503), .ZN(new_n992));
  AOI21_X1  g567(.A(G1384), .B1(new_n992), .B2(new_n872), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n975), .B1(new_n993), .B2(new_n972), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n994), .A3(new_n778), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n984), .B1(new_n987), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n579), .A2(new_n580), .A3(G8), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT55), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n579), .A2(new_n580), .A3(new_n999), .A4(G8), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  MUX2_X1   g576(.A(new_n983), .B(new_n996), .S(new_n1001), .Z(new_n1002));
  NAND4_X1  g577(.A1(new_n600), .A2(new_n603), .A3(new_n700), .A4(new_n605), .ZN(new_n1003));
  INV_X1    g578(.A(new_n599), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n601), .A2(new_n602), .ZN(new_n1005));
  OAI21_X1  g580(.A(G1981), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT118), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n468), .A2(new_n480), .A3(G40), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n874), .A2(new_n973), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G8), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1010), .A2(KEYINPUT116), .A3(G8), .ZN(new_n1014));
  AOI22_X1  g589(.A1(KEYINPUT49), .A2(new_n1008), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT49), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1007), .A2(KEYINPUT118), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1976), .ZN(new_n1018));
  OR2_X1    g593(.A1(G288), .A2(new_n1018), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1010), .A2(KEYINPUT116), .A3(G8), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT116), .B1(new_n1010), .B2(G8), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1015), .A2(new_n1017), .B1(KEYINPUT52), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT52), .B1(G288), .B2(new_n1018), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1019), .B(new_n1024), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1028), .A2(KEYINPUT117), .A3(new_n1019), .A4(new_n1024), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT45), .B1(new_n874), .B2(new_n973), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1009), .B1(new_n976), .B2(new_n980), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n771), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G2084), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n974), .A2(new_n977), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(G286), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1002), .A2(new_n1023), .A3(new_n1030), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT63), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT119), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(new_n1043), .A3(new_n1040), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1023), .A2(new_n1030), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n983), .A2(new_n1001), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n983), .A2(new_n1001), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(new_n1040), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1045), .A2(new_n1046), .A3(new_n1038), .A4(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1042), .A2(new_n1044), .A3(new_n1049), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1051));
  OR2_X1    g626(.A1(G288), .A2(G1976), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1003), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1045), .A2(new_n1047), .B1(new_n1053), .B2(new_n1028), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G286), .A2(G8), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT123), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1055), .B(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1037), .A2(new_n1058), .A3(new_n1059), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1036), .A2(new_n1057), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n984), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1060), .B(new_n1061), .C1(new_n1065), .C2(new_n1057), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n985), .B2(G2078), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n874), .A2(new_n973), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n980), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1032), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1068), .A2(G2078), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n974), .A2(new_n977), .ZN(new_n1075));
  INV_X1    g650(.A(G1961), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1074), .A2(new_n1077), .A3(KEYINPUT125), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT125), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1069), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(G301), .B(KEYINPUT54), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1076), .B2(new_n1075), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1070), .A2(KEYINPUT114), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1070), .A2(KEYINPUT114), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1084), .A2(new_n1085), .A3(KEYINPUT45), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n979), .A2(new_n1009), .A3(new_n1073), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1083), .B(new_n1069), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1067), .A2(new_n1082), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1002), .A2(new_n1023), .A3(new_n1030), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1010), .ZN(new_n1092));
  INV_X1    g667(.A(G2067), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1075), .A2(new_n836), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(new_n628), .ZN(new_n1095));
  INV_X1    g670(.A(G1956), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n972), .B1(new_n874), .B2(new_n973), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1009), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n979), .A2(new_n981), .A3(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n563), .B(KEYINPUT9), .ZN(new_n1102));
  INV_X1    g677(.A(new_n571), .ZN(new_n1103));
  OR2_X1    g678(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1104));
  NAND2_X1  g679(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(KEYINPUT120), .B(KEYINPUT57), .C1(new_n565), .C2(new_n571), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1099), .A2(new_n1101), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1095), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1106), .ZN(new_n1110));
  AOI21_X1  g685(.A(G1956), .B1(new_n991), .B2(new_n994), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n979), .A2(new_n981), .A3(new_n1100), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(KEYINPUT61), .A3(new_n1108), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT58), .B(G1341), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n985), .A2(G1996), .B1(new_n1092), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n555), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n1117), .B2(new_n555), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1115), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1094), .A2(KEYINPUT60), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1075), .A2(new_n836), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n1124), .A3(KEYINPUT60), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n919), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1094), .A2(KEYINPUT60), .A3(new_n628), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1122), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1121), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1113), .A2(new_n1108), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT121), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n1133));
  AOI211_X1 g708(.A(new_n1133), .B(KEYINPUT61), .C1(new_n1113), .C2(new_n1108), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1114), .B1(new_n1129), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1091), .B1(new_n1136), .B2(KEYINPUT122), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1114), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT61), .B1(new_n1113), .B2(new_n1108), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT121), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1117), .A2(new_n555), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT59), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1117), .A2(new_n1118), .A3(new_n555), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n628), .B1(new_n1094), .B2(KEYINPUT60), .ZN(new_n1145));
  AND4_X1   g720(.A1(KEYINPUT60), .A2(new_n1123), .A3(new_n1124), .A4(new_n628), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1115), .B(new_n1144), .C1(new_n1147), .C2(new_n1122), .ZN(new_n1148));
  OAI211_X1 g723(.A(KEYINPUT122), .B(new_n1138), .C1(new_n1140), .C2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1050), .B(new_n1054), .C1(new_n1137), .C2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1138), .B1(new_n1140), .B2(new_n1148), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1156), .A2(new_n1149), .A3(new_n1091), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1157), .A2(KEYINPUT126), .A3(new_n1050), .A4(new_n1054), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1067), .A2(KEYINPUT62), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT127), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1090), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1067), .A2(KEYINPUT62), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1080), .A2(G171), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1153), .A2(new_n1158), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1086), .A2(new_n1009), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT115), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n721), .A2(new_n723), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n721), .A2(new_n723), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n826), .B(G2067), .ZN(new_n1172));
  INV_X1    g747(.A(G1996), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1172), .B1(new_n1173), .B2(new_n795), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1167), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1166), .A2(G1996), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n795), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1171), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1166), .ZN(new_n1179));
  XNOR2_X1  g754(.A(G290), .B(G1986), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1165), .A2(new_n1181), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1166), .A2(G1986), .A3(G290), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT48), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1178), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1176), .B(KEYINPUT46), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1172), .A2(new_n795), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1186), .B1(new_n1167), .B2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1188), .B(KEYINPUT47), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n826), .A2(new_n1093), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1190), .B1(new_n1191), .B2(new_n1169), .ZN(new_n1192));
  AOI211_X1 g767(.A(new_n1185), .B(new_n1189), .C1(new_n1167), .C2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1182), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g769(.A1(G401), .A2(G227), .A3(new_n460), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n707), .A2(new_n708), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n1197), .B1(new_n902), .B2(new_n904), .ZN(new_n1198));
  AND2_X1   g772(.A1(new_n1198), .A2(new_n966), .ZN(G308));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n966), .ZN(G225));
endmodule


