//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G101), .ZN(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT65), .B1(new_n195), .B2(G143), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G146), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n195), .A2(KEYINPUT64), .A3(G143), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT64), .B1(new_n195), .B2(G143), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n196), .B(new_n199), .C1(new_n200), .C2(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G143), .B(G146), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n202), .A2(new_n205), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G137), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G134), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT11), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n211), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT66), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n209), .A2(G137), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n208), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n217), .A2(KEYINPUT66), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n210), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n213), .B1(new_n215), .B2(new_n218), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n224), .A2(new_n225), .A3(G131), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n207), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n216), .A2(new_n221), .A3(new_n208), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n208), .B1(new_n213), .B2(new_n210), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n195), .A2(G143), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(KEYINPUT1), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n196), .A2(new_n199), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n195), .A2(KEYINPUT64), .A3(G143), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n233), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT1), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n198), .A2(G146), .ZN(new_n241));
  AND4_X1   g055(.A1(new_n240), .A2(new_n232), .A3(new_n241), .A4(G128), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n228), .B(new_n230), .C1(new_n239), .C2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G116), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT68), .B1(new_n244), .B2(G119), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n246));
  INV_X1    g060(.A(G119), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(G116), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(G119), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n245), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G113), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT2), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT2), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G113), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(new_n254), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n257), .A2(new_n245), .A3(new_n249), .A4(new_n248), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n227), .A2(new_n243), .A3(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(KEYINPUT28), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT67), .B1(new_n226), .B2(new_n229), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n228), .A2(new_n264), .A3(new_n230), .ZN(new_n265));
  INV_X1    g079(.A(new_n233), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n202), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n232), .A2(new_n241), .A3(new_n240), .A4(G128), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n263), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n227), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n259), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n194), .B1(new_n262), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n194), .A2(KEYINPUT70), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(new_n227), .B2(new_n243), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n242), .B1(new_n202), .B2(new_n266), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n213), .A2(new_n215), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT66), .B(KEYINPUT11), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n279), .B(new_n210), .C1(new_n280), .C2(new_n213), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n230), .B1(new_n281), .B2(G131), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n278), .B1(new_n282), .B2(KEYINPUT67), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(G131), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n228), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n283), .A2(new_n265), .B1(new_n285), .B2(new_n207), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n277), .B1(new_n286), .B2(new_n276), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n261), .B(new_n275), .C1(new_n287), .C2(new_n260), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT31), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n261), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n270), .A2(new_n276), .A3(new_n227), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n227), .A2(new_n243), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT30), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n291), .B1(new_n295), .B2(new_n259), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(KEYINPUT31), .A3(new_n275), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n273), .B1(new_n290), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(G472), .A2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n187), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT71), .ZN(new_n302));
  INV_X1    g116(.A(new_n273), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT31), .B1(new_n296), .B2(new_n275), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n260), .B1(new_n292), .B2(new_n294), .ZN(new_n305));
  NOR4_X1   g119(.A1(new_n305), .A2(new_n289), .A3(new_n291), .A4(new_n274), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n303), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT32), .A3(new_n299), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n194), .A2(KEYINPUT29), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT28), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n261), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n261), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n293), .A2(new_n259), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n227), .A2(new_n243), .A3(KEYINPUT73), .A4(new_n260), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  AOI211_X1 g132(.A(new_n310), .B(new_n313), .C1(new_n318), .C2(KEYINPUT28), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n309), .B1(new_n319), .B2(G902), .ZN(new_n320));
  INV_X1    g134(.A(G902), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(KEYINPUT28), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n312), .ZN(new_n323));
  OAI211_X1 g137(.A(KEYINPUT74), .B(new_n321), .C1(new_n323), .C2(new_n310), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n291), .A2(KEYINPUT28), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n325), .A2(new_n272), .A3(new_n194), .A4(new_n312), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n262), .A2(KEYINPUT72), .A3(new_n194), .A4(new_n272), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n193), .B1(new_n305), .B2(new_n291), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n328), .A2(new_n329), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n320), .A2(new_n324), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G472), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT71), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n335), .B(new_n187), .C1(new_n298), .C2(new_n300), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n302), .A2(new_n308), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(G475), .A2(G902), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G113), .B(G122), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(G104), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT95), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G237), .ZN(new_n344));
  INV_X1    g158(.A(G953), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(G214), .ZN(new_n346));
  NOR2_X1   g160(.A1(KEYINPUT94), .A2(G143), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n189), .B(G214), .C1(KEYINPUT94), .C2(G143), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(KEYINPUT18), .A3(G131), .ZN(new_n351));
  XNOR2_X1  g165(.A(G125), .B(G140), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(new_n195), .ZN(new_n353));
  NAND2_X1  g167(.A1(KEYINPUT18), .A2(G131), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n348), .A2(new_n349), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n208), .B1(new_n348), .B2(new_n349), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT96), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT17), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n358), .B1(new_n357), .B2(KEYINPUT17), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n350), .A2(G131), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT17), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n348), .A2(new_n349), .A3(new_n208), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G140), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G125), .ZN(new_n367));
  INV_X1    g181(.A(G125), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G140), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT16), .ZN(new_n370));
  OR3_X1    g184(.A1(new_n368), .A2(KEYINPUT16), .A3(G140), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(G146), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(G146), .B1(new_n370), .B2(new_n371), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n365), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n343), .B(new_n356), .C1(new_n361), .C2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT19), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n352), .B(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n372), .B1(new_n379), .B2(G146), .ZN(new_n380));
  INV_X1    g194(.A(new_n364), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(new_n357), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n356), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n341), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n339), .B1(new_n377), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT97), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT20), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n386), .B1(new_n385), .B2(new_n387), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n385), .A2(new_n387), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT9), .B(G234), .ZN(new_n392));
  INV_X1    g206(.A(G217), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n392), .A2(new_n393), .A3(G953), .ZN(new_n394));
  INV_X1    g208(.A(G122), .ZN(new_n395));
  OR3_X1    g209(.A1(new_n395), .A2(KEYINPUT14), .A3(G116), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n244), .A2(G122), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT14), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n395), .A2(G116), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n396), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G107), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n198), .A2(G128), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n231), .A2(G143), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G134), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n403), .A3(new_n209), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G107), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n399), .A2(new_n397), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n401), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT13), .B1(new_n198), .B2(G128), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n402), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT98), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT98), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n415), .A3(new_n402), .ZN(new_n416));
  INV_X1    g230(.A(new_n402), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT13), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G134), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n399), .A2(new_n397), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G107), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n409), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n423), .A2(new_n406), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n411), .B1(new_n425), .B2(KEYINPUT99), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT99), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n420), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n394), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n413), .A2(KEYINPUT98), .B1(KEYINPUT13), .B2(new_n417), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n209), .B1(new_n430), .B2(new_n416), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n423), .A2(new_n406), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT99), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n433), .A2(new_n428), .A3(new_n410), .A4(new_n394), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n321), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G478), .ZN(new_n437));
  NOR2_X1   g251(.A1(KEYINPUT100), .A2(KEYINPUT15), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(KEYINPUT100), .A2(KEYINPUT15), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n394), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n433), .A2(new_n410), .ZN(new_n444));
  INV_X1    g258(.A(new_n428), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(G902), .B1(new_n446), .B2(new_n434), .ZN(new_n447));
  INV_X1    g261(.A(new_n441), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(G234), .A2(G237), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(G952), .A3(new_n345), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n450), .A2(G902), .A3(G953), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(G898), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(new_n455), .B(KEYINPUT101), .Z(new_n456));
  NAND3_X1  g270(.A1(new_n442), .A2(new_n449), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n356), .B1(new_n361), .B2(new_n376), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n341), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n377), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n321), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G475), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n391), .A2(new_n457), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G214), .B1(G237), .B2(G902), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n466));
  INV_X1    g280(.A(G104), .ZN(new_n467));
  OAI21_X1  g281(.A(KEYINPUT3), .B1(new_n467), .B2(G107), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n408), .A3(G104), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(G107), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G101), .ZN(new_n473));
  INV_X1    g287(.A(G101), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n468), .A2(new_n470), .A3(new_n474), .A4(new_n471), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(KEYINPUT4), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT4), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n472), .A2(new_n477), .A3(G101), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n259), .A3(new_n478), .ZN(new_n479));
  OR2_X1    g293(.A1(KEYINPUT87), .A2(KEYINPUT5), .ZN(new_n480));
  NAND2_X1  g294(.A1(KEYINPUT87), .A2(KEYINPUT5), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n480), .A2(G116), .A3(new_n247), .A4(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n480), .A2(new_n481), .ZN(new_n483));
  OAI211_X1 g297(.A(G113), .B(new_n482), .C1(new_n250), .C2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(G104), .B(G107), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT82), .B1(new_n485), .B2(new_n474), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n408), .A2(G104), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n471), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT82), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n489), .A3(G101), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n484), .A2(new_n491), .A3(new_n258), .A4(new_n475), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n479), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(G110), .B(G122), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n466), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n479), .A2(new_n492), .A3(new_n494), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT89), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n479), .A2(new_n492), .A3(KEYINPUT89), .A4(new_n494), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n493), .A2(KEYINPUT88), .A3(new_n495), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT90), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n498), .A2(new_n503), .A3(KEYINPUT90), .A4(new_n504), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n493), .A2(new_n466), .A3(new_n495), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n269), .A2(new_n368), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n207), .A2(G125), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n345), .A2(G224), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n512), .B(new_n514), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n507), .A2(new_n508), .A3(new_n509), .A4(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT91), .B(KEYINPUT8), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n494), .B(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n486), .A2(new_n490), .B1(new_n519), .B2(new_n474), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n258), .B2(new_n484), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n521), .B(KEYINPUT92), .Z(new_n522));
  INV_X1    g336(.A(KEYINPUT5), .ZN(new_n523));
  OAI211_X1 g337(.A(G113), .B(new_n482), .C1(new_n250), .C2(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n520), .A2(new_n258), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n518), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT93), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n512), .A2(new_n527), .A3(KEYINPUT7), .A4(new_n513), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n510), .B(new_n511), .C1(new_n527), .C2(new_n514), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT7), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n529), .B1(new_n530), .B2(new_n514), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n528), .A2(new_n531), .B1(new_n501), .B2(new_n502), .ZN(new_n532));
  AOI21_X1  g346(.A(G902), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(G210), .B1(G237), .B2(G902), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n516), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n516), .B2(new_n533), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n464), .B(new_n465), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n375), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n231), .A2(G119), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n247), .A2(G128), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT24), .B(G110), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT23), .B1(new_n231), .B2(G119), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n231), .A2(G119), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n231), .A2(KEYINPUT23), .A3(G119), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n544), .B1(new_n549), .B2(G110), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n539), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G110), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n547), .A2(KEYINPUT75), .A3(new_n552), .A4(new_n548), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n542), .A2(new_n543), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT23), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n247), .B2(G128), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n556), .A2(new_n548), .A3(new_n552), .A4(new_n541), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT75), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n553), .A2(new_n554), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT76), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n557), .A2(new_n558), .B1(new_n542), .B2(new_n543), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(KEYINPUT76), .A3(new_n553), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n352), .A2(new_n195), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n372), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT77), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT77), .ZN(new_n570));
  AOI211_X1 g384(.A(new_n570), .B(new_n567), .C1(new_n562), .C2(new_n564), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n551), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT22), .B(G137), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n345), .A2(G221), .A3(G234), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n573), .B(new_n574), .Z(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT78), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n393), .B1(G234), .B2(new_n321), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(G902), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT79), .ZN(new_n581));
  INV_X1    g395(.A(new_n575), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n551), .B(new_n582), .C1(new_n569), .C2(new_n571), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n578), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n551), .ZN(new_n586));
  INV_X1    g400(.A(new_n564), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT76), .B1(new_n563), .B2(new_n553), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n568), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n570), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n565), .A2(KEYINPUT77), .A3(new_n568), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n586), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n583), .B(new_n321), .C1(new_n592), .C2(new_n576), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT25), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n578), .A2(KEYINPUT25), .A3(new_n321), .A4(new_n583), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n585), .B1(new_n597), .B2(new_n579), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT85), .ZN(new_n599));
  XNOR2_X1  g413(.A(G110), .B(G140), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n345), .A2(G227), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n600), .B(new_n601), .Z(new_n602));
  XOR2_X1   g416(.A(new_n602), .B(KEYINPUT81), .Z(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n268), .B1(new_n233), .B2(new_n206), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n485), .A2(KEYINPUT82), .A3(new_n474), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n489), .B1(new_n488), .B2(G101), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n605), .B(new_n475), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n269), .B2(new_n520), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT12), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT84), .B1(new_n284), .B2(new_n228), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n610), .B1(new_n609), .B2(new_n611), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n269), .A2(new_n520), .A3(KEYINPUT10), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n608), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n222), .A2(new_n226), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n207), .A2(new_n476), .A3(new_n478), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n615), .A2(new_n617), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n604), .B1(new_n614), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n602), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n615), .A2(new_n617), .A3(new_n619), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n622), .B1(new_n285), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n599), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n609), .A2(new_n611), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT12), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n620), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n620), .A2(new_n602), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n623), .A2(new_n285), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n629), .A2(new_n603), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT85), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n625), .A2(new_n633), .A3(G469), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n622), .A2(KEYINPUT86), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT86), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n620), .A2(new_n636), .A3(new_n602), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n614), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n631), .A2(new_n620), .ZN(new_n639));
  INV_X1    g453(.A(new_n602), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(G469), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n643), .A3(new_n321), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n321), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n634), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(G221), .B1(new_n392), .B2(G902), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT80), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n337), .A2(new_n538), .A3(new_n598), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT102), .B(G101), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G3));
  OAI21_X1  g469(.A(G472), .B1(new_n298), .B2(G902), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n307), .A2(new_n299), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n597), .A2(new_n579), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n584), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n658), .A2(new_n651), .A3(new_n660), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n465), .B(new_n456), .C1(new_n535), .C2(new_n536), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n437), .A2(new_n321), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n447), .B2(new_n437), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n426), .A2(new_n428), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT33), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n446), .A2(new_n434), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n665), .B1(new_n671), .B2(G478), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n389), .A2(new_n390), .ZN(new_n673));
  INV_X1    g487(.A(new_n388), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n462), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n662), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n661), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT34), .B(G104), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G6));
  XNOR2_X1  g495(.A(new_n385), .B(new_n387), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n682), .A2(new_n462), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n448), .B1(new_n670), .B2(new_n321), .ZN(new_n684));
  AOI211_X1 g498(.A(G902), .B(new_n441), .C1(new_n446), .C2(new_n434), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n662), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n661), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT104), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT35), .B(G107), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G9));
  OR2_X1    g507(.A1(new_n577), .A2(KEYINPUT36), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n592), .B(new_n694), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n695), .A2(new_n581), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n579), .B2(new_n597), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n651), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n658), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n538), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT37), .B(G110), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G12));
  OAI21_X1  g516(.A(new_n465), .B1(new_n535), .B2(new_n536), .ZN(new_n703));
  INV_X1    g517(.A(G900), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n452), .B1(new_n453), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n683), .A2(new_n687), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(KEYINPUT105), .B1(new_n703), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n516), .A2(new_n533), .ZN(new_n709));
  INV_X1    g523(.A(new_n534), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n516), .A2(new_n533), .A3(new_n534), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n707), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n713), .A2(new_n714), .A3(new_n715), .A4(new_n465), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n708), .A2(new_n716), .A3(new_n337), .A4(new_n698), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G128), .ZN(G30));
  XOR2_X1   g532(.A(new_n705), .B(KEYINPUT39), .Z(new_n719));
  NAND2_X1  g533(.A1(new_n652), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n720), .B(KEYINPUT40), .Z(new_n721));
  AOI21_X1  g535(.A(new_n686), .B1(new_n675), .B2(new_n462), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n697), .A2(new_n465), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT107), .ZN(new_n724));
  INV_X1    g538(.A(new_n318), .ZN(new_n725));
  AOI21_X1  g539(.A(G902), .B1(new_n725), .B2(new_n193), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n194), .B1(new_n305), .B2(new_n291), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G472), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n302), .A2(new_n308), .A3(new_n336), .A4(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n535), .A2(new_n536), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n732), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n713), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n721), .A2(new_n724), .A3(new_n730), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G143), .ZN(G45));
  NAND3_X1  g552(.A1(new_n672), .A2(new_n676), .A3(new_n706), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n703), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n337), .A2(new_n740), .A3(new_n698), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G146), .ZN(G48));
  NAND2_X1  g556(.A1(new_n627), .A2(new_n628), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n636), .B1(new_n620), .B2(new_n602), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n745), .A2(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n746));
  OAI21_X1  g560(.A(G469), .B1(new_n746), .B2(G902), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n650), .A3(new_n644), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n678), .A2(new_n337), .A3(new_n598), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT41), .B(G113), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(G15));
  NAND4_X1  g566(.A1(new_n689), .A2(new_n337), .A3(new_n598), .A4(new_n749), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G116), .ZN(G18));
  INV_X1    g568(.A(new_n659), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n464), .B1(new_n755), .B2(new_n696), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n335), .B1(new_n657), .B2(new_n187), .ZN(new_n757));
  AOI211_X1 g571(.A(KEYINPUT71), .B(KEYINPUT32), .C1(new_n307), .C2(new_n299), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n334), .A2(new_n308), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n756), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT108), .B1(new_n703), .B2(new_n748), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n713), .A2(new_n749), .A3(new_n763), .A4(new_n465), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G119), .ZN(G21));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n768));
  AND4_X1   g582(.A1(new_n456), .A2(new_n747), .A3(new_n650), .A4(new_n644), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n323), .A2(new_n193), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n304), .B2(new_n306), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n299), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n769), .A2(new_n598), .A3(new_n656), .A4(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n722), .B(new_n465), .C1(new_n535), .C2(new_n536), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n768), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n774), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n598), .A2(new_n656), .A3(new_n772), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n776), .A2(new_n777), .A3(KEYINPUT109), .A4(new_n769), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G122), .ZN(G24));
  NAND2_X1  g594(.A1(new_n656), .A2(new_n772), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n739), .A3(new_n697), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n765), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G125), .ZN(G27));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n645), .B1(new_n632), .B2(G469), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n649), .B1(new_n644), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n731), .A2(new_n785), .A3(new_n465), .A4(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n711), .A2(new_n787), .A3(new_n465), .A4(new_n712), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT110), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n739), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n337), .A3(new_n598), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT42), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n660), .B1(new_n759), .B2(new_n760), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(KEYINPUT111), .A3(new_n792), .A4(new_n791), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n760), .A2(new_n301), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n739), .A2(new_n796), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n791), .A2(new_n598), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G131), .ZN(G33));
  NAND3_X1  g618(.A1(new_n797), .A2(new_n714), .A3(new_n791), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  NAND2_X1  g620(.A1(new_n731), .A2(new_n465), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n391), .A2(new_n463), .ZN(new_n808));
  NOR2_X1   g622(.A1(KEYINPUT113), .A2(KEYINPUT43), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT113), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT43), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n672), .B(new_n808), .C1(new_n809), .C2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n669), .A2(new_n670), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n669), .A2(new_n670), .ZN(new_n815));
  OAI21_X1  g629(.A(G478), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n664), .ZN(new_n817));
  OAI22_X1  g631(.A1(new_n817), .A2(new_n676), .B1(new_n810), .B2(new_n811), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n819), .B(new_n658), .C1(new_n755), .C2(new_n696), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT44), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n807), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT46), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n625), .A2(new_n633), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT45), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n643), .B1(new_n632), .B2(KEYINPUT45), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n824), .B(new_n825), .C1(new_n830), .C2(new_n645), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n645), .B1(new_n828), .B2(new_n829), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT112), .B1(new_n832), .B2(KEYINPUT46), .ZN(new_n833));
  INV_X1    g647(.A(new_n644), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n832), .B2(KEYINPUT46), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n650), .A3(new_n719), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n823), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(KEYINPUT114), .B(G137), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n838), .B(new_n839), .ZN(G39));
  NAND2_X1  g654(.A1(new_n836), .A2(new_n650), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT47), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n836), .A2(KEYINPUT47), .A3(new_n650), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n337), .A2(new_n807), .A3(new_n598), .A4(new_n739), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G140), .ZN(G42));
  INV_X1    g662(.A(new_n465), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n817), .A2(new_n676), .A3(new_n849), .A4(new_n649), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n747), .A2(new_n644), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n850), .B1(KEYINPUT49), .B2(new_n851), .ZN(new_n852));
  AOI211_X1 g666(.A(new_n852), .B(new_n736), .C1(KEYINPUT49), .C2(new_n851), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n730), .A2(new_n660), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n775), .A2(new_n778), .B1(new_n761), .B2(new_n765), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n651), .A2(new_n660), .ZN(new_n857));
  INV_X1    g671(.A(new_n662), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n808), .A2(new_n687), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n677), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n857), .A2(new_n858), .A3(new_n699), .A4(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n653), .A2(new_n861), .A3(new_n700), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n750), .A2(new_n753), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n856), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n686), .A2(new_n462), .A3(new_n682), .A4(new_n706), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n535), .A2(new_n536), .A3(new_n865), .A4(new_n849), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n337), .A2(new_n698), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n337), .A2(new_n698), .A3(new_n866), .A4(KEYINPUT115), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n791), .A2(new_n782), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n805), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n864), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n717), .A2(new_n741), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT52), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n697), .A2(new_n706), .A3(new_n787), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n730), .A3(new_n776), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n875), .A2(new_n876), .A3(new_n783), .A4(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n783), .A2(new_n878), .A3(new_n717), .A4(new_n741), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT52), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n874), .A2(new_n803), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT116), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n779), .A2(new_n766), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n653), .A2(new_n861), .A3(new_n700), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n750), .A2(new_n753), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n871), .A2(new_n805), .A3(new_n872), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n879), .A2(new_n888), .A3(new_n889), .A4(new_n881), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT53), .A4(new_n803), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n882), .A2(new_n883), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n884), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(KEYINPUT117), .A3(KEYINPUT54), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT117), .B1(new_n894), .B2(KEYINPUT54), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n890), .A2(KEYINPUT53), .A3(new_n803), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n893), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n896), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n749), .A2(new_n849), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT118), .B1(new_n736), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n903), .B1(new_n733), .B2(new_n735), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n819), .A2(new_n777), .A3(new_n452), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n904), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n909), .A2(KEYINPUT119), .A3(KEYINPUT50), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT50), .B1(new_n909), .B2(KEYINPUT119), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n902), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n908), .B1(new_n905), .B2(new_n906), .ZN(new_n913));
  INV_X1    g727(.A(new_n907), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT119), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT50), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n909), .A2(KEYINPUT119), .A3(KEYINPUT50), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(KEYINPUT120), .A3(new_n918), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n807), .A2(new_n451), .A3(new_n748), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n854), .A2(new_n920), .A3(new_n808), .A4(new_n817), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n781), .A2(new_n697), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n920), .A2(new_n819), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n843), .B(new_n844), .C1(new_n650), .C2(new_n851), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n908), .A2(new_n465), .A3(new_n731), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n912), .A2(new_n919), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT51), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n800), .A2(new_n598), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n924), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT48), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n854), .A2(new_n920), .A3(new_n676), .A4(new_n672), .ZN(new_n937));
  INV_X1    g751(.A(G952), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n938), .B(G953), .C1(new_n908), .C2(new_n765), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  AOI211_X1 g754(.A(new_n930), .B(new_n925), .C1(new_n926), .C2(new_n927), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n910), .A2(new_n911), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n931), .A2(new_n932), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n932), .B1(new_n931), .B2(new_n943), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT122), .B1(new_n901), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n894), .A2(KEYINPUT54), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT117), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n900), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n950), .A2(KEYINPUT122), .A3(new_n895), .A4(new_n946), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n938), .A2(new_n345), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n855), .B1(new_n947), .B2(new_n953), .ZN(G75));
  NOR2_X1   g768(.A1(new_n345), .A2(G952), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n321), .B1(new_n898), .B2(new_n893), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT56), .B1(new_n957), .B2(G210), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n515), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT55), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n956), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n899), .A2(G902), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT123), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n957), .A2(KEYINPUT123), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n710), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT56), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n961), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n962), .B1(new_n968), .B2(new_n970), .ZN(G51));
  XNOR2_X1  g785(.A(new_n899), .B(KEYINPUT54), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n645), .B(KEYINPUT57), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n642), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n967), .A2(new_n830), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n955), .B1(new_n975), .B2(new_n976), .ZN(G54));
  NAND4_X1  g791(.A1(new_n965), .A2(KEYINPUT58), .A3(G475), .A4(new_n966), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n377), .A2(new_n384), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n978), .A2(KEYINPUT124), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n956), .B1(new_n978), .B2(new_n980), .ZN(new_n982));
  AOI21_X1  g796(.A(KEYINPUT124), .B1(new_n978), .B2(new_n980), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(G60));
  INV_X1    g798(.A(new_n671), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n950), .A2(new_n895), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n663), .B(KEYINPUT59), .Z(new_n987));
  AOI21_X1  g801(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n972), .A2(new_n985), .A3(new_n987), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n988), .A2(new_n955), .A3(new_n989), .ZN(G63));
  NAND2_X1  g804(.A1(G217), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT60), .Z(new_n992));
  NAND2_X1  g806(.A1(new_n899), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n578), .A2(new_n583), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n955), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n695), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n995), .B1(new_n996), .B2(new_n993), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT61), .Z(G66));
  NAND2_X1  g812(.A1(G224), .A2(G953), .ZN(new_n999));
  OAI22_X1  g813(.A1(new_n864), .A2(G953), .B1(new_n454), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n959), .B1(G898), .B2(new_n345), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1000), .B(new_n1001), .Z(G69));
  NAND3_X1  g816(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n295), .B(new_n379), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n875), .A2(new_n783), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n737), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n1006), .A2(KEYINPUT62), .ZN(new_n1007));
  AOI211_X1 g821(.A(new_n807), .B(new_n720), .C1(new_n677), .C2(new_n859), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n838), .B1(new_n797), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1006), .A2(KEYINPUT62), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1007), .A2(new_n847), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1003), .B(new_n1004), .C1(new_n1011), .C2(G953), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n838), .B1(new_n845), .B2(new_n846), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n837), .A2(new_n774), .A3(new_n933), .ZN(new_n1014));
  INV_X1    g828(.A(new_n805), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1013), .A2(new_n803), .A3(new_n1016), .A4(new_n1005), .ZN(new_n1017));
  OR2_X1    g831(.A1(new_n1017), .A2(KEYINPUT125), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(KEYINPUT125), .ZN(new_n1019));
  AOI21_X1  g833(.A(G953), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n704), .A2(new_n345), .A3(G227), .ZN(new_n1021));
  OR2_X1    g835(.A1(new_n1004), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1012), .B1(new_n1020), .B2(new_n1022), .ZN(G72));
  NAND3_X1  g837(.A1(new_n1018), .A2(new_n888), .A3(new_n1019), .ZN(new_n1024));
  NAND2_X1  g838(.A1(G472), .A2(G902), .ZN(new_n1025));
  XOR2_X1   g839(.A(new_n1025), .B(KEYINPUT63), .Z(new_n1026));
  NAND2_X1  g840(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g841(.A1(new_n305), .A2(new_n194), .A3(new_n291), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1026), .B1(new_n1011), .B2(new_n864), .ZN(new_n1030));
  INV_X1    g844(.A(new_n727), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1029), .A2(new_n956), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g847(.A(KEYINPUT126), .B1(new_n1031), .B2(new_n1028), .ZN(new_n1034));
  OAI211_X1 g848(.A(new_n1034), .B(new_n1026), .C1(KEYINPUT126), .C2(new_n331), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1035), .B(KEYINPUT127), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1033), .B1(new_n894), .B2(new_n1036), .ZN(G57));
endmodule


