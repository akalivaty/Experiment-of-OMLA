

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575;

  XNOR2_X1 U319 ( .A(n313), .B(n312), .ZN(n512) );
  XOR2_X1 U320 ( .A(n333), .B(n332), .Z(n287) );
  XOR2_X1 U321 ( .A(KEYINPUT33), .B(n413), .Z(n288) );
  XNOR2_X1 U322 ( .A(KEYINPUT54), .B(KEYINPUT116), .ZN(n403) );
  XNOR2_X1 U323 ( .A(n334), .B(n287), .ZN(n335) );
  XNOR2_X1 U324 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U325 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U326 ( .A(n439), .B(G190GAT), .ZN(n440) );
  XNOR2_X1 U327 ( .A(n441), .B(n440), .ZN(G1351GAT) );
  XOR2_X1 U328 ( .A(KEYINPUT1), .B(KEYINPUT88), .Z(n290) );
  XNOR2_X1 U329 ( .A(G148GAT), .B(G85GAT), .ZN(n289) );
  XNOR2_X1 U330 ( .A(n290), .B(n289), .ZN(n292) );
  XOR2_X1 U331 ( .A(G29GAT), .B(G162GAT), .Z(n291) );
  XNOR2_X1 U332 ( .A(n292), .B(n291), .ZN(n311) );
  XOR2_X1 U333 ( .A(KEYINPUT0), .B(KEYINPUT79), .Z(n294) );
  XNOR2_X1 U334 ( .A(G134GAT), .B(KEYINPUT80), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U336 ( .A(n295), .B(G127GAT), .Z(n297) );
  XNOR2_X1 U337 ( .A(G113GAT), .B(G120GAT), .ZN(n296) );
  XNOR2_X1 U338 ( .A(n297), .B(n296), .ZN(n437) );
  XOR2_X1 U339 ( .A(KEYINPUT92), .B(KEYINPUT90), .Z(n299) );
  XNOR2_X1 U340 ( .A(KEYINPUT89), .B(KEYINPUT91), .ZN(n298) );
  XNOR2_X1 U341 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U342 ( .A(n437), .B(n300), .ZN(n304) );
  XOR2_X1 U343 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n302) );
  XNOR2_X1 U344 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U346 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U347 ( .A(n305), .B(G57GAT), .Z(n309) );
  XOR2_X1 U348 ( .A(G155GAT), .B(KEYINPUT2), .Z(n307) );
  XNOR2_X1 U349 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n306) );
  XNOR2_X1 U350 ( .A(n307), .B(n306), .ZN(n409) );
  XNOR2_X1 U351 ( .A(n409), .B(KEYINPUT6), .ZN(n308) );
  XNOR2_X1 U352 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U353 ( .A(n311), .B(n310), .ZN(n313) );
  NAND2_X1 U354 ( .A1(G225GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U355 ( .A(G211GAT), .B(G218GAT), .ZN(n314) );
  XNOR2_X1 U356 ( .A(n314), .B(KEYINPUT21), .ZN(n315) );
  XOR2_X1 U357 ( .A(n315), .B(KEYINPUT86), .Z(n317) );
  XNOR2_X1 U358 ( .A(G197GAT), .B(G204GAT), .ZN(n316) );
  XNOR2_X1 U359 ( .A(n317), .B(n316), .ZN(n418) );
  XOR2_X1 U360 ( .A(G183GAT), .B(KEYINPUT19), .Z(n319) );
  XNOR2_X1 U361 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n318) );
  XNOR2_X1 U362 ( .A(n319), .B(n318), .ZN(n433) );
  XOR2_X1 U363 ( .A(n433), .B(KEYINPUT94), .Z(n321) );
  NAND2_X1 U364 ( .A1(G226GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U365 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U366 ( .A(G36GAT), .B(G190GAT), .Z(n342) );
  XOR2_X1 U367 ( .A(n322), .B(n342), .Z(n325) );
  XOR2_X1 U368 ( .A(G169GAT), .B(G8GAT), .Z(n388) );
  XNOR2_X1 U369 ( .A(G176GAT), .B(G92GAT), .ZN(n323) );
  XNOR2_X1 U370 ( .A(n323), .B(G64GAT), .ZN(n331) );
  XNOR2_X1 U371 ( .A(n388), .B(n331), .ZN(n324) );
  XNOR2_X1 U372 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U373 ( .A(n418), .B(n326), .ZN(n501) );
  XNOR2_X1 U374 ( .A(G120GAT), .B(G204GAT), .ZN(n327) );
  XOR2_X1 U375 ( .A(G99GAT), .B(G85GAT), .Z(n350) );
  XNOR2_X1 U376 ( .A(n327), .B(n350), .ZN(n338) );
  XNOR2_X1 U377 ( .A(G106GAT), .B(G78GAT), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n328), .B(G148GAT), .ZN(n413) );
  NAND2_X1 U379 ( .A1(G230GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n288), .B(n329), .ZN(n336) );
  XNOR2_X1 U381 ( .A(G71GAT), .B(G57GAT), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n330), .B(KEYINPUT13), .ZN(n360) );
  XNOR2_X1 U383 ( .A(n331), .B(n360), .ZN(n334) );
  XOR2_X1 U384 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n333) );
  XNOR2_X1 U385 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n332) );
  XOR2_X1 U386 ( .A(n338), .B(n337), .Z(n563) );
  XOR2_X1 U387 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n340) );
  XNOR2_X1 U388 ( .A(KEYINPUT74), .B(KEYINPUT10), .ZN(n339) );
  XNOR2_X1 U389 ( .A(n340), .B(n339), .ZN(n346) );
  XNOR2_X1 U390 ( .A(G50GAT), .B(KEYINPUT71), .ZN(n341) );
  XNOR2_X1 U391 ( .A(n341), .B(G162GAT), .ZN(n410) );
  XOR2_X1 U392 ( .A(n342), .B(n410), .Z(n344) );
  NAND2_X1 U393 ( .A1(G232GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U394 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U395 ( .A(n346), .B(n345), .ZN(n359) );
  XOR2_X1 U396 ( .A(KEYINPUT76), .B(G92GAT), .Z(n348) );
  XNOR2_X1 U397 ( .A(G218GAT), .B(G106GAT), .ZN(n347) );
  XNOR2_X1 U398 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U399 ( .A(n349), .B(KEYINPUT72), .Z(n352) );
  XNOR2_X1 U400 ( .A(G134GAT), .B(n350), .ZN(n351) );
  XNOR2_X1 U401 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U402 ( .A(n353), .B(KEYINPUT75), .Z(n357) );
  XOR2_X1 U403 ( .A(G29GAT), .B(G43GAT), .Z(n355) );
  XNOR2_X1 U404 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n354) );
  XNOR2_X1 U405 ( .A(n355), .B(n354), .ZN(n385) );
  XNOR2_X1 U406 ( .A(n385), .B(KEYINPUT73), .ZN(n356) );
  XNOR2_X1 U407 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U408 ( .A(n359), .B(n358), .Z(n538) );
  XOR2_X1 U409 ( .A(KEYINPUT36), .B(n538), .Z(n572) );
  XOR2_X1 U410 ( .A(n360), .B(G155GAT), .Z(n362) );
  NAND2_X1 U411 ( .A1(G231GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U412 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U413 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n364) );
  XNOR2_X1 U414 ( .A(G8GAT), .B(KEYINPUT14), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U416 ( .A(n366), .B(n365), .Z(n371) );
  XOR2_X1 U417 ( .A(G64GAT), .B(G78GAT), .Z(n368) );
  XNOR2_X1 U418 ( .A(G127GAT), .B(G183GAT), .ZN(n367) );
  XNOR2_X1 U419 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U420 ( .A(G211GAT), .B(n369), .ZN(n370) );
  XNOR2_X1 U421 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U422 ( .A(n372), .B(KEYINPUT12), .Z(n376) );
  XOR2_X1 U423 ( .A(KEYINPUT66), .B(G1GAT), .Z(n374) );
  XNOR2_X1 U424 ( .A(G22GAT), .B(G15GAT), .ZN(n373) );
  XNOR2_X1 U425 ( .A(n374), .B(n373), .ZN(n384) );
  XNOR2_X1 U426 ( .A(n384), .B(KEYINPUT77), .ZN(n375) );
  XOR2_X1 U427 ( .A(n376), .B(n375), .Z(n569) );
  NOR2_X1 U428 ( .A1(n572), .A2(n569), .ZN(n377) );
  XOR2_X1 U429 ( .A(KEYINPUT45), .B(n377), .Z(n378) );
  NOR2_X1 U430 ( .A1(n563), .A2(n378), .ZN(n394) );
  XOR2_X1 U431 ( .A(KEYINPUT29), .B(G113GAT), .Z(n380) );
  XNOR2_X1 U432 ( .A(G197GAT), .B(G141GAT), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n380), .B(n379), .ZN(n393) );
  XOR2_X1 U434 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n382) );
  NAND2_X1 U435 ( .A1(G229GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U437 ( .A(n383), .B(KEYINPUT65), .Z(n387) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U439 ( .A(n387), .B(n386), .ZN(n389) );
  XOR2_X1 U440 ( .A(n389), .B(n388), .Z(n391) );
  XNOR2_X1 U441 ( .A(G50GAT), .B(G36GAT), .ZN(n390) );
  XNOR2_X1 U442 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U443 ( .A(n393), .B(n392), .Z(n557) );
  NAND2_X1 U444 ( .A1(n394), .A2(n557), .ZN(n401) );
  INV_X1 U445 ( .A(KEYINPUT46), .ZN(n396) );
  XOR2_X1 U446 ( .A(KEYINPUT41), .B(n563), .Z(n547) );
  INV_X1 U447 ( .A(n557), .ZN(n542) );
  NAND2_X1 U448 ( .A1(n547), .A2(n542), .ZN(n395) );
  XOR2_X1 U449 ( .A(n396), .B(n395), .Z(n398) );
  INV_X1 U450 ( .A(n569), .ZN(n550) );
  NOR2_X1 U451 ( .A1(n550), .A2(n538), .ZN(n397) );
  AND2_X1 U452 ( .A1(n398), .A2(n397), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n399), .B(KEYINPUT47), .ZN(n400) );
  NAND2_X1 U454 ( .A1(n401), .A2(n400), .ZN(n402) );
  XNOR2_X1 U455 ( .A(KEYINPUT48), .B(n402), .ZN(n511) );
  NAND2_X1 U456 ( .A1(n501), .A2(n511), .ZN(n404) );
  NOR2_X1 U457 ( .A1(n512), .A2(n405), .ZN(n556) );
  XOR2_X1 U458 ( .A(KEYINPUT84), .B(KEYINPUT23), .Z(n407) );
  NAND2_X1 U459 ( .A1(G228GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U460 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U461 ( .A(n408), .B(KEYINPUT24), .Z(n412) );
  XNOR2_X1 U462 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U463 ( .A(n412), .B(n411), .ZN(n417) );
  XOR2_X1 U464 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n415) );
  XNOR2_X1 U465 ( .A(KEYINPUT87), .B(n413), .ZN(n414) );
  XNOR2_X1 U466 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U467 ( .A(n417), .B(n416), .Z(n420) );
  XNOR2_X1 U468 ( .A(G22GAT), .B(n418), .ZN(n419) );
  XNOR2_X1 U469 ( .A(n420), .B(n419), .ZN(n448) );
  AND2_X1 U470 ( .A1(n556), .A2(n448), .ZN(n421) );
  XNOR2_X1 U471 ( .A(KEYINPUT55), .B(n421), .ZN(n438) );
  XOR2_X1 U472 ( .A(G71GAT), .B(KEYINPUT20), .Z(n423) );
  XNOR2_X1 U473 ( .A(G15GAT), .B(KEYINPUT81), .ZN(n422) );
  XNOR2_X1 U474 ( .A(n423), .B(n422), .ZN(n431) );
  NAND2_X1 U475 ( .A1(G227GAT), .A2(G233GAT), .ZN(n429) );
  XOR2_X1 U476 ( .A(KEYINPUT64), .B(KEYINPUT82), .Z(n425) );
  XNOR2_X1 U477 ( .A(G99GAT), .B(KEYINPUT83), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n427) );
  XOR2_X1 U479 ( .A(G43GAT), .B(G190GAT), .Z(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U481 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U482 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U483 ( .A(n432), .B(G176GAT), .Z(n435) );
  XNOR2_X1 U484 ( .A(G169GAT), .B(n433), .ZN(n434) );
  XNOR2_X1 U485 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X2 U486 ( .A(n437), .B(n436), .Z(n503) );
  INV_X1 U487 ( .A(n503), .ZN(n518) );
  NOR2_X2 U488 ( .A1(n438), .A2(n518), .ZN(n551) );
  NAND2_X1 U489 ( .A1(n551), .A2(n538), .ZN(n441) );
  XOR2_X1 U490 ( .A(KEYINPUT58), .B(KEYINPUT121), .Z(n439) );
  NOR2_X1 U491 ( .A1(n563), .A2(n557), .ZN(n442) );
  XOR2_X1 U492 ( .A(n442), .B(KEYINPUT70), .Z(n470) );
  NOR2_X1 U493 ( .A1(n538), .A2(n569), .ZN(n443) );
  XNOR2_X1 U494 ( .A(KEYINPUT16), .B(n443), .ZN(n458) );
  XOR2_X1 U495 ( .A(n448), .B(KEYINPUT28), .Z(n505) );
  INV_X1 U496 ( .A(n505), .ZN(n516) );
  XOR2_X1 U497 ( .A(KEYINPUT27), .B(n501), .Z(n514) );
  NOR2_X1 U498 ( .A1(n503), .A2(n514), .ZN(n444) );
  NAND2_X1 U499 ( .A1(n516), .A2(n444), .ZN(n445) );
  NAND2_X1 U500 ( .A1(n445), .A2(n512), .ZN(n456) );
  NAND2_X1 U501 ( .A1(n503), .A2(n501), .ZN(n446) );
  NAND2_X1 U502 ( .A1(n448), .A2(n446), .ZN(n447) );
  XOR2_X1 U503 ( .A(KEYINPUT25), .B(n447), .Z(n454) );
  XNOR2_X1 U504 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n450) );
  NOR2_X1 U505 ( .A1(n503), .A2(n448), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U507 ( .A(KEYINPUT95), .B(n451), .ZN(n527) );
  NOR2_X1 U508 ( .A1(n527), .A2(n514), .ZN(n452) );
  NOR2_X1 U509 ( .A1(n512), .A2(n452), .ZN(n453) );
  NAND2_X1 U510 ( .A1(n454), .A2(n453), .ZN(n455) );
  NAND2_X1 U511 ( .A1(n456), .A2(n455), .ZN(n457) );
  XNOR2_X1 U512 ( .A(KEYINPUT97), .B(n457), .ZN(n468) );
  NAND2_X1 U513 ( .A1(n458), .A2(n468), .ZN(n484) );
  NOR2_X1 U514 ( .A1(n470), .A2(n484), .ZN(n465) );
  NAND2_X1 U515 ( .A1(n465), .A2(n512), .ZN(n461) );
  XNOR2_X1 U516 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n459), .B(KEYINPUT34), .ZN(n460) );
  XNOR2_X1 U518 ( .A(n461), .B(n460), .ZN(G1324GAT) );
  NAND2_X1 U519 ( .A1(n501), .A2(n465), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n462), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U521 ( .A(G15GAT), .B(KEYINPUT35), .Z(n464) );
  NAND2_X1 U522 ( .A1(n465), .A2(n503), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n464), .B(n463), .ZN(G1326GAT) );
  NAND2_X1 U524 ( .A1(n465), .A2(n505), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n466), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U526 ( .A1(n572), .A2(n550), .ZN(n467) );
  NAND2_X1 U527 ( .A1(n468), .A2(n467), .ZN(n469) );
  XOR2_X1 U528 ( .A(KEYINPUT37), .B(n469), .Z(n499) );
  OR2_X1 U529 ( .A1(n499), .A2(n470), .ZN(n471) );
  XOR2_X1 U530 ( .A(KEYINPUT38), .B(n471), .Z(n481) );
  NAND2_X1 U531 ( .A1(n481), .A2(n512), .ZN(n474) );
  XNOR2_X1 U532 ( .A(G29GAT), .B(KEYINPUT99), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n472), .B(KEYINPUT39), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(G1328GAT) );
  NAND2_X1 U535 ( .A1(n481), .A2(n501), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n475), .B(KEYINPUT100), .ZN(n476) );
  XNOR2_X1 U537 ( .A(G36GAT), .B(n476), .ZN(G1329GAT) );
  XNOR2_X1 U538 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n480) );
  XOR2_X1 U539 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n478) );
  NAND2_X1 U540 ( .A1(n503), .A2(n481), .ZN(n477) );
  XNOR2_X1 U541 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n480), .B(n479), .ZN(G1330GAT) );
  NAND2_X1 U543 ( .A1(n505), .A2(n481), .ZN(n482) );
  XNOR2_X1 U544 ( .A(G50GAT), .B(n482), .ZN(G1331GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT42), .B(KEYINPUT105), .Z(n487) );
  INV_X1 U546 ( .A(n547), .ZN(n533) );
  NOR2_X1 U547 ( .A1(n533), .A2(n542), .ZN(n483) );
  XNOR2_X1 U548 ( .A(n483), .B(KEYINPUT103), .ZN(n498) );
  NOR2_X1 U549 ( .A1(n484), .A2(n498), .ZN(n485) );
  XNOR2_X1 U550 ( .A(n485), .B(KEYINPUT104), .ZN(n494) );
  NAND2_X1 U551 ( .A1(n512), .A2(n494), .ZN(n486) );
  XNOR2_X1 U552 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U553 ( .A(G57GAT), .B(n488), .ZN(G1332GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n490) );
  NAND2_X1 U555 ( .A1(n494), .A2(n501), .ZN(n489) );
  XNOR2_X1 U556 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U557 ( .A(G64GAT), .B(n491), .ZN(G1333GAT) );
  NAND2_X1 U558 ( .A1(n494), .A2(n503), .ZN(n492) );
  XNOR2_X1 U559 ( .A(n492), .B(KEYINPUT108), .ZN(n493) );
  XNOR2_X1 U560 ( .A(G71GAT), .B(n493), .ZN(G1334GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n496) );
  NAND2_X1 U562 ( .A1(n505), .A2(n494), .ZN(n495) );
  XNOR2_X1 U563 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U564 ( .A(G78GAT), .B(n497), .Z(G1335GAT) );
  NOR2_X1 U565 ( .A1(n499), .A2(n498), .ZN(n506) );
  NAND2_X1 U566 ( .A1(n512), .A2(n506), .ZN(n500) );
  XNOR2_X1 U567 ( .A(G85GAT), .B(n500), .ZN(G1336GAT) );
  NAND2_X1 U568 ( .A1(n501), .A2(n506), .ZN(n502) );
  XNOR2_X1 U569 ( .A(n502), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U570 ( .A1(n506), .A2(n503), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n504), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U572 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n510) );
  XOR2_X1 U573 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n508) );
  NAND2_X1 U574 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1339GAT) );
  NAND2_X1 U577 ( .A1(n512), .A2(n511), .ZN(n513) );
  NOR2_X1 U578 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U579 ( .A(KEYINPUT112), .B(n515), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n528), .A2(n516), .ZN(n517) );
  NOR2_X1 U581 ( .A1(n518), .A2(n517), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n524), .A2(n542), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G113GAT), .B(n519), .ZN(G1340GAT) );
  XOR2_X1 U584 ( .A(G120GAT), .B(KEYINPUT49), .Z(n521) );
  NAND2_X1 U585 ( .A1(n524), .A2(n547), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n521), .B(n520), .ZN(G1341GAT) );
  NAND2_X1 U587 ( .A1(n524), .A2(n550), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(KEYINPUT50), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G127GAT), .B(n523), .ZN(G1342GAT) );
  XOR2_X1 U590 ( .A(G134GAT), .B(KEYINPUT51), .Z(n526) );
  NAND2_X1 U591 ( .A1(n524), .A2(n538), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(G1343GAT) );
  INV_X1 U593 ( .A(n527), .ZN(n555) );
  NAND2_X1 U594 ( .A1(n555), .A2(n528), .ZN(n539) );
  NOR2_X1 U595 ( .A1(n557), .A2(n539), .ZN(n530) );
  XNOR2_X1 U596 ( .A(G141GAT), .B(KEYINPUT113), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(G1344GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n532) );
  XNOR2_X1 U599 ( .A(G148GAT), .B(KEYINPUT114), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n532), .B(n531), .ZN(n535) );
  NOR2_X1 U601 ( .A1(n533), .A2(n539), .ZN(n534) );
  XOR2_X1 U602 ( .A(n535), .B(n534), .Z(G1345GAT) );
  NOR2_X1 U603 ( .A1(n569), .A2(n539), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G155GAT), .B(KEYINPUT115), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(G1346GAT) );
  INV_X1 U606 ( .A(n538), .ZN(n540) );
  NOR2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U608 ( .A(G162GAT), .B(n541), .Z(G1347GAT) );
  NAND2_X1 U609 ( .A1(n542), .A2(n551), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n543), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT57), .B(KEYINPUT118), .Z(n545) );
  XNOR2_X1 U612 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U614 ( .A(KEYINPUT117), .B(n546), .Z(n549) );
  NAND2_X1 U615 ( .A1(n547), .A2(n551), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1349GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n553) );
  NAND2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G183GAT), .B(n554), .ZN(G1350GAT) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n571) );
  NOR2_X1 U622 ( .A1(n557), .A2(n571), .ZN(n562) );
  XOR2_X1 U623 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n559) );
  XNOR2_X1 U624 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(KEYINPUT60), .B(n560), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1352GAT) );
  INV_X1 U628 ( .A(n563), .ZN(n564) );
  NOR2_X1 U629 ( .A1(n571), .A2(n564), .ZN(n568) );
  XOR2_X1 U630 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n566) );
  XNOR2_X1 U631 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1353GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n571), .ZN(n570) );
  XOR2_X1 U635 ( .A(G211GAT), .B(n570), .Z(G1354GAT) );
  NOR2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n574) );
  XNOR2_X1 U637 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U639 ( .A(G218GAT), .B(n575), .Z(G1355GAT) );
endmodule

