//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G107), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT77), .ZN(new_n194));
  AOI21_X1  g008(.A(KEYINPUT3), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n194), .A2(new_n189), .A3(KEYINPUT3), .A4(G104), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n191), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G101), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n189), .A2(G104), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(KEYINPUT77), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(new_n196), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(new_n189), .B2(G104), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT78), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT78), .ZN(new_n208));
  AOI211_X1 g022(.A(new_n208), .B(new_n205), .C1(new_n202), .C2(new_n196), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n199), .B(KEYINPUT4), .C1(new_n207), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT0), .A4(G128), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT0), .B(G128), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n190), .B1(new_n202), .B2(new_n196), .ZN(new_n220));
  OR2_X1    g034(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n204), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT80), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT80), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n198), .A2(new_n226), .A3(new_n223), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n210), .A2(new_n219), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G137), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT11), .A3(G134), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(G137), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G131), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(KEYINPUT64), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n236), .B(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n206), .B1(new_n195), .B2(new_n197), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n208), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n203), .A2(KEYINPUT78), .A3(new_n206), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT10), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n204), .B1(new_n191), .B2(new_n201), .ZN(new_n246));
  INV_X1    g060(.A(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT1), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n212), .A3(new_n214), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT65), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n216), .A2(new_n251), .A3(new_n248), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  OAI22_X1  g067(.A1(new_n248), .A2(new_n214), .B1(new_n212), .B2(G128), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n246), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n244), .A2(new_n245), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n245), .B1(new_n244), .B2(new_n256), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n229), .B(new_n240), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT81), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n251), .B1(new_n216), .B2(new_n248), .ZN(new_n261));
  AND4_X1   g075(.A1(new_n251), .A2(new_n248), .A3(new_n212), .A4(new_n214), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n255), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n246), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n263), .B(new_n264), .C1(new_n207), .C2(new_n209), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT10), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n244), .A2(new_n245), .A3(new_n256), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT81), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n268), .A2(new_n269), .A3(new_n240), .A4(new_n229), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n260), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G227), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n273), .B(KEYINPUT76), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G140), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n246), .B1(new_n242), .B2(new_n243), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n265), .B1(new_n278), .B2(new_n263), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n239), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT12), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(KEYINPUT12), .A3(new_n239), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n271), .A2(new_n277), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n268), .A2(new_n229), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n239), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n277), .B1(new_n271), .B2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n187), .B(new_n188), .C1(new_n285), .C2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n187), .A2(new_n188), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n271), .A2(new_n284), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n276), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n276), .B1(new_n260), .B2(new_n270), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n287), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(G469), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n289), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G221), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT9), .B(G234), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n298), .B1(new_n300), .B2(new_n188), .ZN(new_n301));
  XOR2_X1   g115(.A(new_n301), .B(KEYINPUT75), .Z(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT82), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT82), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n297), .A2(new_n306), .A3(new_n303), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT25), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n247), .A2(G119), .ZN(new_n310));
  INV_X1    g124(.A(G119), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G128), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n313), .B1(new_n310), .B2(new_n312), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT24), .B(G110), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n312), .A2(KEYINPUT23), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n321));
  OAI22_X1  g135(.A1(new_n318), .A2(new_n320), .B1(new_n310), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n317), .B1(G110), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT16), .ZN(new_n324));
  INV_X1    g138(.A(G140), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(G125), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n326), .B1(new_n330), .B2(new_n324), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n211), .ZN(new_n332));
  OAI211_X1 g146(.A(G146), .B(new_n326), .C1(new_n330), .C2(new_n324), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n323), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n316), .B1(new_n314), .B2(new_n315), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n322), .B2(G110), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n338));
  INV_X1    g152(.A(new_n330), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n211), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n340), .A2(new_n333), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n337), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n338), .B1(new_n337), .B2(new_n341), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n335), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT22), .B(G137), .ZN(new_n345));
  INV_X1    g159(.A(G234), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n298), .A2(new_n346), .A3(G953), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n345), .B(new_n347), .Z(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n335), .B(new_n348), .C1(new_n342), .C2(new_n343), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n309), .B1(new_n352), .B2(G902), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n350), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n351), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G217), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(G234), .B2(new_n188), .ZN(new_n357));
  INV_X1    g171(.A(new_n352), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(G902), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n355), .A2(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n254), .B1(new_n250), .B2(new_n252), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n237), .B1(G134), .B2(new_n233), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n236), .A2(new_n237), .B1(new_n235), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT66), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT66), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n236), .A2(new_n237), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n363), .A2(new_n235), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n263), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n239), .A2(new_n219), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n365), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT30), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT69), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT68), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n311), .A2(G116), .ZN(new_n377));
  INV_X1    g191(.A(G116), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G119), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT2), .B(G113), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n376), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n380), .B1(new_n381), .B2(KEYINPUT67), .ZN(new_n383));
  INV_X1    g197(.A(G113), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT2), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT2), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G113), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT67), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n382), .B1(new_n383), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n389), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n381), .A2(KEYINPUT67), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n392), .A2(new_n393), .A3(new_n376), .A4(new_n380), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n375), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n391), .A2(new_n375), .A3(new_n394), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n369), .A2(KEYINPUT70), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT70), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n364), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n263), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT30), .A3(new_n371), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n374), .A2(new_n398), .A3(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n396), .A2(new_n402), .A3(new_n397), .A4(new_n371), .ZN(new_n405));
  XOR2_X1   g219(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n406));
  NOR2_X1   g220(.A1(G237), .A2(G953), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G210), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n406), .B(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT26), .B(G101), .ZN(new_n410));
  XOR2_X1   g224(.A(new_n409), .B(new_n410), .Z(new_n411));
  NAND3_X1  g225(.A1(new_n404), .A2(new_n405), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT31), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n404), .A2(KEYINPUT31), .A3(new_n405), .A4(new_n411), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n405), .A2(KEYINPUT28), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n391), .A2(new_n375), .A3(new_n394), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(new_n395), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT28), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n371), .A4(new_n402), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n398), .A2(new_n372), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n411), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n414), .A2(new_n415), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G472), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n188), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT32), .ZN(new_n429));
  NOR4_X1   g243(.A1(new_n425), .A2(KEYINPUT32), .A3(G472), .A4(G902), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n423), .A2(new_n424), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n411), .B1(new_n404), .B2(new_n405), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT29), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n402), .A2(new_n371), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n398), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n421), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n411), .A2(KEYINPUT29), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n188), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(G472), .B1(new_n435), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n361), .B1(new_n432), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n443));
  OAI21_X1  g257(.A(G210), .B1(G237), .B2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT85), .B1(new_n219), .B2(new_n328), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n362), .A2(new_n328), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT85), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n218), .A2(new_n448), .A3(G125), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n272), .A2(G224), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n210), .B(new_n228), .C1(new_n417), .C2(new_n395), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n380), .A2(new_n381), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n377), .A2(new_n379), .A3(KEYINPUT5), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n377), .A2(KEYINPUT5), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(new_n384), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n454), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n278), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G110), .B(G122), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n453), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT84), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT6), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n453), .A2(new_n459), .ZN(new_n466));
  INV_X1    g280(.A(new_n460), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  AOI211_X1 g283(.A(new_n460), .B(new_n463), .C1(new_n453), .C2(new_n459), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n452), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n451), .A2(KEYINPUT7), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n450), .B(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n460), .B(KEYINPUT8), .ZN(new_n475));
  INV_X1    g289(.A(new_n459), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n278), .A2(new_n458), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n474), .A2(new_n478), .A3(new_n461), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n188), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n445), .B1(new_n472), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n452), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n460), .B1(new_n453), .B2(new_n459), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n461), .B2(new_n464), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n482), .B1(new_n484), .B2(new_n470), .ZN(new_n485));
  INV_X1    g299(.A(new_n480), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n444), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(G214), .B1(G237), .B2(G902), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n489), .B(KEYINPUT83), .Z(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n443), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  AOI211_X1 g306(.A(KEYINPUT86), .B(new_n490), .C1(new_n481), .C2(new_n487), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n407), .A2(G143), .A3(G214), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(G143), .B1(new_n407), .B2(G214), .ZN(new_n496));
  OAI211_X1 g310(.A(KEYINPUT17), .B(G131), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n332), .A2(new_n497), .A3(new_n333), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G131), .B1(new_n495), .B2(new_n496), .ZN(new_n501));
  INV_X1    g315(.A(new_n496), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n237), .A3(new_n494), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n332), .A2(new_n497), .A3(KEYINPUT90), .A4(new_n333), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n500), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n330), .B(G146), .ZN(new_n508));
  OAI211_X1 g322(.A(KEYINPUT18), .B(G131), .C1(new_n495), .C2(new_n496), .ZN(new_n509));
  NAND2_X1  g323(.A1(KEYINPUT18), .A2(G131), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n502), .A2(new_n494), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G113), .B(G122), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT88), .B(G104), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n514), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT89), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n507), .A2(new_n512), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n517), .B1(new_n507), .B2(new_n512), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n188), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT91), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT91), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n524), .B(new_n188), .C1(new_n520), .C2(new_n521), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(G475), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n501), .A2(new_n503), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT87), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT87), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n501), .A2(new_n503), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n339), .A2(KEYINPUT19), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT19), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n211), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n528), .A2(new_n333), .A3(new_n530), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n512), .ZN(new_n535));
  INV_X1    g349(.A(new_n517), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n537), .A2(new_n519), .ZN(new_n538));
  INV_X1    g352(.A(G475), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n188), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT20), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n519), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n542), .A2(new_n543), .A3(new_n539), .A4(new_n188), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n526), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n213), .A2(G128), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n213), .A2(G128), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n231), .ZN(new_n551));
  XNOR2_X1  g365(.A(G116), .B(G122), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(new_n189), .ZN(new_n553));
  INV_X1    g367(.A(new_n549), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n548), .B2(KEYINPUT13), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(KEYINPUT13), .B2(new_n548), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n551), .B(new_n553), .C1(new_n556), .C2(new_n231), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n378), .A2(KEYINPUT14), .A3(G122), .ZN(new_n558));
  INV_X1    g372(.A(new_n552), .ZN(new_n559));
  OAI211_X1 g373(.A(G107), .B(new_n558), .C1(new_n559), .C2(KEYINPUT14), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n548), .A2(new_n549), .A3(G134), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n550), .A2(new_n231), .ZN(new_n562));
  OAI221_X1 g376(.A(new_n560), .B1(G107), .B2(new_n559), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n299), .A2(new_n356), .A3(G953), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n557), .A2(new_n563), .A3(new_n565), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n188), .ZN(new_n570));
  INV_X1    g384(.A(G478), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(KEYINPUT15), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n570), .B(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n546), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n272), .A2(G952), .ZN(new_n575));
  INV_X1    g389(.A(G237), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n575), .B1(new_n346), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  AOI211_X1 g392(.A(new_n188), .B(new_n272), .C1(G234), .C2(G237), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT21), .B(G898), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n574), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n492), .A2(new_n493), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n308), .A2(new_n442), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  OAI21_X1  g400(.A(G472), .B1(new_n425), .B2(G902), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n428), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n308), .A2(new_n360), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT93), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT33), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(KEYINPUT93), .A2(KEYINPUT33), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n569), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n567), .A2(new_n592), .A3(new_n593), .A4(new_n568), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n571), .A2(G902), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n598), .A2(new_n599), .B1(new_n571), .B2(new_n570), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n526), .B2(new_n545), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n582), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n472), .A2(new_n445), .A3(new_n480), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n444), .B1(new_n485), .B2(new_n486), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n491), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT92), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT92), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n488), .A2(new_n607), .A3(new_n491), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n602), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n591), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT94), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT95), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT34), .B(G104), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  AND3_X1   g428(.A1(new_n526), .A2(new_n545), .A3(new_n573), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n615), .A2(new_n582), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n607), .B1(new_n488), .B2(new_n491), .ZN(new_n617));
  AOI211_X1 g431(.A(KEYINPUT92), .B(new_n490), .C1(new_n481), .C2(new_n487), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n590), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT96), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT35), .B(G107), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  NAND2_X1  g437(.A1(new_n355), .A2(new_n357), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n349), .A2(KEYINPUT36), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n344), .B(new_n625), .Z(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n359), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT97), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n624), .A2(new_n630), .A3(new_n627), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n308), .A2(new_n584), .A3(new_n589), .A4(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT37), .B(G110), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G12));
  NAND2_X1  g450(.A1(new_n606), .A2(new_n608), .ZN(new_n637));
  INV_X1    g451(.A(new_n307), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n306), .B1(new_n297), .B2(new_n303), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n578), .B1(new_n579), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n526), .A2(new_n545), .A3(new_n573), .A4(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT98), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n539), .B1(new_n522), .B2(KEYINPUT91), .ZN(new_n646));
  AOI22_X1  g460(.A1(new_n646), .A2(new_n525), .B1(new_n541), .B2(new_n544), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n647), .A2(new_n648), .A3(new_n573), .A4(new_n643), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT32), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n425), .A2(G902), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(new_n652), .B2(new_n427), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n441), .B1(new_n653), .B2(new_n430), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n633), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n640), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(new_n247), .ZN(G30));
  XOR2_X1   g471(.A(new_n642), .B(KEYINPUT39), .Z(new_n658));
  NAND2_X1  g472(.A1(new_n308), .A2(new_n658), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n659), .A2(KEYINPUT40), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n404), .A2(new_n405), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n411), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n437), .A2(new_n424), .A3(new_n405), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n188), .A3(new_n663), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n429), .A2(new_n431), .B1(G472), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n628), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n488), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n546), .A2(new_n573), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n490), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n666), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n659), .A2(KEYINPUT40), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n660), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n213), .ZN(G45));
  INV_X1    g488(.A(new_n655), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n601), .A2(new_n643), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n308), .A2(new_n675), .A3(new_n637), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  NAND2_X1  g493(.A1(new_n271), .A2(new_n287), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n680), .A2(new_n276), .B1(new_n294), .B2(new_n284), .ZN(new_n681));
  OAI21_X1  g495(.A(G469), .B1(new_n681), .B2(G902), .ZN(new_n682));
  INV_X1    g496(.A(new_n301), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n683), .A3(new_n289), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT100), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n682), .A2(KEYINPUT100), .A3(new_n683), .A4(new_n289), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n687), .B1(new_n686), .B2(new_n688), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n691), .A2(KEYINPUT102), .A3(new_n442), .A4(new_n609), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n686), .A2(new_n688), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT101), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n694), .A2(new_n442), .A3(new_n609), .A4(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  NAND2_X1  g515(.A1(new_n654), .A2(new_n360), .ZN(new_n702));
  NOR4_X1   g516(.A1(new_n689), .A2(new_n690), .A3(new_n702), .A4(new_n619), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n378), .ZN(G18));
  NAND4_X1  g518(.A1(new_n633), .A2(new_n654), .A3(new_n582), .A4(new_n574), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n617), .A2(new_n618), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT103), .B1(new_n693), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n637), .A2(new_n708), .A3(new_n686), .A4(new_n688), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n705), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n311), .ZN(G21));
  XOR2_X1   g525(.A(KEYINPUT105), .B(G472), .Z(new_n712));
  OAI21_X1  g526(.A(new_n712), .B1(new_n425), .B2(G902), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n414), .A2(new_n415), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n438), .A2(new_n424), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n427), .A2(new_n188), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT104), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n713), .A2(new_n719), .A3(new_n360), .A4(new_n582), .ZN(new_n720));
  AOI211_X1 g534(.A(new_n669), .B(new_n720), .C1(new_n606), .C2(new_n608), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n694), .A2(new_n721), .A3(new_n695), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  AND2_X1   g537(.A1(new_n713), .A2(new_n719), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n677), .A2(new_n628), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n707), .B2(new_n709), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n328), .ZN(G27));
  AOI22_X1  g541(.A1(new_n292), .A2(new_n276), .B1(new_n294), .B2(new_n287), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n290), .B1(new_n728), .B2(G469), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n301), .B1(new_n729), .B2(new_n289), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n488), .A2(new_n490), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n442), .A2(new_n732), .A3(new_n677), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n442), .A2(new_n732), .A3(KEYINPUT42), .A4(new_n677), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  NAND2_X1  g552(.A1(new_n650), .A2(KEYINPUT106), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n645), .A2(new_n649), .A3(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n442), .A2(new_n732), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  OAI21_X1  g557(.A(G469), .B1(new_n728), .B2(KEYINPUT45), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT107), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n746), .B(G469), .C1(new_n728), .C2(KEYINPUT45), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n728), .A2(KEYINPUT45), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT108), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n745), .A2(new_n751), .A3(new_n747), .A4(new_n748), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n290), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n753), .A2(KEYINPUT46), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n289), .B1(new_n753), .B2(KEYINPUT46), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n600), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n647), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g572(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n647), .B(new_n757), .C1(new_n761), .C2(KEYINPUT43), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n588), .A3(new_n628), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  INV_X1    g581(.A(new_n731), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n756), .A2(new_n769), .A3(new_n683), .A4(new_n658), .ZN(new_n770));
  XOR2_X1   g584(.A(KEYINPUT110), .B(G137), .Z(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(G39));
  OAI21_X1  g586(.A(new_n683), .B1(new_n754), .B2(new_n755), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(KEYINPUT47), .B(new_n683), .C1(new_n754), .C2(new_n755), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n677), .A2(new_n731), .A3(new_n361), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n654), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT111), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n781));
  INV_X1    g595(.A(new_n779), .ZN(new_n782));
  AOI211_X1 g596(.A(new_n781), .B(new_n782), .C1(new_n775), .C2(new_n776), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n582), .B1(new_n615), .B2(new_n601), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n492), .A2(new_n493), .A3(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n308), .A2(new_n788), .A3(new_n360), .A4(new_n589), .ZN(new_n789));
  AND4_X1   g603(.A1(new_n585), .A2(new_n722), .A3(new_n634), .A4(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n703), .A2(new_n710), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n699), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n640), .A2(new_n655), .A3(new_n676), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n726), .A2(new_n656), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n706), .A2(new_n669), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n666), .A3(new_n643), .A4(new_n730), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n707), .A2(new_n709), .ZN(new_n799));
  INV_X1    g613(.A(new_n725), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n656), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n802), .A3(new_n678), .A4(new_n797), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT52), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n731), .A2(new_n574), .A3(new_n643), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n305), .B2(new_n307), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n675), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n800), .A2(new_n732), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n807), .A2(new_n742), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n737), .A2(new_n810), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n806), .A2(new_n675), .B1(new_n800), .B2(new_n732), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n808), .B1(new_n812), .B2(new_n742), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n792), .A2(new_n798), .A3(new_n804), .A4(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT52), .B1(new_n726), .B2(new_n656), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT53), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n815), .A2(KEYINPUT114), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT114), .B1(new_n815), .B2(new_n819), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n786), .B(new_n818), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n815), .A2(new_n819), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n816), .A2(new_n819), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n823), .B1(new_n815), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT54), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n724), .A2(new_n360), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n577), .B1(new_n760), .B2(new_n762), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n829), .A2(KEYINPUT115), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(KEYINPUT115), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n693), .A2(new_n491), .A3(new_n668), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n832), .A2(KEYINPUT50), .A3(new_n833), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n693), .A2(new_n768), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT116), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n665), .A2(new_n360), .A3(new_n578), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n840), .A2(new_n647), .A3(new_n600), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n830), .A2(new_n831), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n840), .A2(new_n628), .A3(new_n724), .A4(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n838), .A2(new_n843), .A3(new_n845), .A4(KEYINPUT51), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n682), .A2(new_n302), .A3(new_n289), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n775), .A2(KEYINPUT117), .A3(new_n776), .A4(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n832), .A2(new_n731), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n775), .A2(new_n776), .A3(new_n847), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n846), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n840), .A2(new_n601), .A3(new_n842), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n799), .A2(new_n832), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n575), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n840), .A2(new_n442), .A3(new_n844), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n858), .A2(KEYINPUT48), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(KEYINPUT48), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n838), .A2(new_n843), .A3(new_n845), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n851), .B2(new_n849), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n861), .B1(new_n863), .B2(KEYINPUT51), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n854), .A2(new_n864), .ZN(new_n865));
  OAI22_X1  g679(.A1(new_n827), .A2(new_n865), .B1(G952), .B2(G953), .ZN(new_n866));
  NOR4_X1   g680(.A1(new_n361), .A2(new_n758), .A3(new_n302), .A4(new_n490), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n682), .A2(new_n289), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n868), .A2(KEYINPUT112), .B1(KEYINPUT49), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT112), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n668), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n869), .A2(KEYINPUT49), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n870), .A2(new_n665), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n866), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT118), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n866), .A2(new_n877), .A3(new_n874), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(G75));
  NOR2_X1   g693(.A1(new_n272), .A2(G952), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n882), .A2(G210), .A3(G902), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n484), .A2(new_n470), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n452), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n485), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n881), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT56), .B1(new_n883), .B2(KEYINPUT119), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(KEYINPUT119), .B2(new_n883), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n890), .B1(new_n892), .B2(new_n888), .ZN(G51));
  XNOR2_X1  g707(.A(new_n882), .B(new_n786), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n290), .B(KEYINPUT57), .Z(new_n895));
  OAI22_X1  g709(.A1(new_n894), .A2(new_n895), .B1(new_n288), .B2(new_n285), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n750), .A2(new_n752), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT120), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n882), .A2(G902), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n880), .B1(new_n896), .B2(new_n899), .ZN(G54));
  AND4_X1   g714(.A1(KEYINPUT58), .A2(new_n882), .A3(G475), .A4(G902), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n881), .B1(new_n901), .B2(new_n542), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n542), .B2(new_n901), .ZN(G60));
  XOR2_X1   g717(.A(new_n598), .B(KEYINPUT121), .Z(new_n904));
  NAND2_X1  g718(.A1(G478), .A2(G902), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT59), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n881), .B1(new_n894), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n904), .B1(new_n827), .B2(new_n906), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(G63));
  NAND2_X1  g724(.A1(G217), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT60), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n882), .A2(new_n626), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT114), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n823), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n815), .A2(KEYINPUT114), .A3(new_n819), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n912), .B1(new_n918), .B2(new_n818), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n914), .B(new_n881), .C1(new_n919), .C2(new_n358), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(KEYINPUT122), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(KEYINPUT122), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT123), .Z(new_n924));
  AND3_X1   g738(.A1(new_n920), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n924), .B1(new_n920), .B2(new_n922), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(G66));
  INV_X1    g741(.A(new_n580), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n272), .B1(new_n928), .B2(G224), .ZN(new_n929));
  INV_X1    g743(.A(new_n792), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n930), .B2(new_n272), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n885), .B1(G898), .B2(new_n272), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT124), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n933), .ZN(G69));
  NOR2_X1   g748(.A1(new_n272), .A2(G900), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n702), .A2(new_n706), .A3(new_n669), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n756), .A2(new_n683), .A3(new_n658), .A4(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n737), .A2(new_n742), .ZN(new_n938));
  AND4_X1   g752(.A1(new_n770), .A2(new_n937), .A3(new_n794), .A4(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n780), .B2(new_n783), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n935), .B1(new_n940), .B2(new_n272), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(G227), .A2(G900), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n374), .A2(new_n403), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n531), .A2(new_n532), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n943), .A2(G953), .A3(new_n944), .A4(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n941), .A2(new_n942), .ZN(new_n949));
  AOI211_X1 g763(.A(KEYINPUT126), .B(new_n935), .C1(new_n940), .C2(new_n272), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n944), .A2(G953), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n442), .B(new_n731), .C1(new_n601), .C2(new_n615), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n770), .B1(new_n659), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT125), .Z(new_n955));
  INV_X1    g769(.A(new_n673), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n794), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT62), .Z(new_n958));
  NAND3_X1  g772(.A1(new_n955), .A2(new_n784), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n947), .A2(G953), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n951), .A2(new_n952), .A3(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n948), .A2(new_n962), .ZN(G72));
  INV_X1    g777(.A(new_n959), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n792), .ZN(new_n965));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  AOI21_X1  g781(.A(new_n662), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n940), .B2(new_n930), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n969), .A2(new_n405), .A3(new_n424), .A4(new_n404), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n412), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(new_n434), .Z(new_n973));
  AND2_X1   g787(.A1(new_n973), .A2(new_n967), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n880), .B1(new_n825), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n968), .A2(new_n976), .ZN(G57));
endmodule


