

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718;

  AND2_X1 U367 ( .A1(n366), .A2(n365), .ZN(n642) );
  XNOR2_X1 U368 ( .A(n407), .B(n353), .ZN(n697) );
  XNOR2_X1 U369 ( .A(KEYINPUT8), .B(KEYINPUT68), .ZN(n440) );
  XNOR2_X1 U370 ( .A(n697), .B(n380), .ZN(n379) );
  INV_X2 U371 ( .A(G143), .ZN(n371) );
  XNOR2_X1 U372 ( .A(n379), .B(n491), .ZN(n670) );
  XNOR2_X1 U373 ( .A(n494), .B(n493), .ZN(n570) );
  NOR2_X1 U374 ( .A1(n492), .A2(n670), .ZN(n494) );
  XNOR2_X1 U375 ( .A(n442), .B(n441), .ZN(n443) );
  INV_X1 U376 ( .A(G119), .ZN(n410) );
  NOR2_X2 U377 ( .A1(G953), .A2(G237), .ZN(n464) );
  NOR2_X1 U378 ( .A1(n582), .A2(n581), .ZN(n399) );
  XNOR2_X1 U379 ( .A(n607), .B(n385), .ZN(n618) );
  BUF_X1 U380 ( .A(n607), .Z(n370) );
  XNOR2_X1 U381 ( .A(n386), .B(n349), .ZN(n607) );
  XNOR2_X1 U382 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X1 U383 ( .A1(G902), .A2(n676), .ZN(n439) );
  XNOR2_X1 U384 ( .A(n482), .B(n484), .ZN(n485) );
  XNOR2_X1 U385 ( .A(n443), .B(n444), .ZN(n476) );
  XNOR2_X1 U386 ( .A(n410), .B(G110), .ZN(n488) );
  XNOR2_X1 U387 ( .A(n383), .B(G125), .ZN(n483) );
  INV_X4 U388 ( .A(G953), .ZN(n706) );
  BUF_X1 U389 ( .A(n688), .Z(n346) );
  INV_X1 U390 ( .A(n593), .ZN(n347) );
  XNOR2_X1 U391 ( .A(n399), .B(n583), .ZN(n611) );
  NAND2_X1 U392 ( .A1(n627), .A2(n692), .ZN(n637) );
  OR2_X1 U393 ( .A1(n604), .A2(n596), .ZN(n619) );
  XNOR2_X1 U394 ( .A(n483), .B(n382), .ZN(n461) );
  INV_X1 U395 ( .A(KEYINPUT10), .ZN(n382) );
  XNOR2_X1 U396 ( .A(n454), .B(n453), .ZN(n455) );
  INV_X1 U397 ( .A(KEYINPUT25), .ZN(n453) );
  OR2_X1 U398 ( .A1(n636), .A2(G902), .ZN(n386) );
  XOR2_X1 U399 ( .A(G104), .B(G122), .Z(n486) );
  XOR2_X1 U400 ( .A(KEYINPUT94), .B(KEYINPUT11), .Z(n466) );
  XOR2_X1 U401 ( .A(KEYINPUT95), .B(KEYINPUT12), .Z(n463) );
  INV_X1 U402 ( .A(KEYINPUT85), .ZN(n374) );
  XOR2_X1 U403 ( .A(KEYINPUT5), .B(KEYINPUT75), .Z(n426) );
  XNOR2_X1 U404 ( .A(G137), .B(G116), .ZN(n428) );
  XNOR2_X1 U405 ( .A(n408), .B(KEYINPUT3), .ZN(n487) );
  XNOR2_X1 U406 ( .A(G113), .B(G101), .ZN(n408) );
  XNOR2_X1 U407 ( .A(KEYINPUT73), .B(KEYINPUT16), .ZN(n490) );
  XNOR2_X1 U408 ( .A(n406), .B(G107), .ZN(n489) );
  INV_X1 U409 ( .A(G116), .ZN(n406) );
  XNOR2_X1 U410 ( .A(n489), .B(n478), .ZN(n394) );
  XNOR2_X1 U411 ( .A(G134), .B(G122), .ZN(n478) );
  XNOR2_X1 U412 ( .A(n472), .B(n471), .ZN(n681) );
  XNOR2_X1 U413 ( .A(n437), .B(G101), .ZN(n418) );
  XOR2_X1 U414 ( .A(G110), .B(G107), .Z(n437) );
  XNOR2_X1 U415 ( .A(n433), .B(n432), .ZN(n435) );
  INV_X1 U416 ( .A(G104), .ZN(n432) );
  AND2_X1 U417 ( .A1(n659), .A2(n387), .ZN(n568) );
  NOR2_X1 U418 ( .A1(n618), .A2(n388), .ZN(n387) );
  INV_X1 U419 ( .A(n549), .ZN(n389) );
  BUF_X1 U420 ( .A(n570), .Z(n372) );
  XNOR2_X1 U421 ( .A(n401), .B(n400), .ZN(n582) );
  INV_X1 U422 ( .A(KEYINPUT19), .ZN(n400) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n563) );
  INV_X1 U424 ( .A(KEYINPUT107), .ZN(n367) );
  XNOR2_X1 U425 ( .A(n480), .B(G478), .ZN(n544) );
  XNOR2_X1 U426 ( .A(n504), .B(n360), .ZN(n559) );
  INV_X1 U427 ( .A(KEYINPUT98), .ZN(n360) );
  NAND2_X1 U428 ( .A1(n546), .A2(n544), .ZN(n504) );
  BUF_X1 U429 ( .A(n621), .Z(n363) );
  INV_X1 U430 ( .A(KEYINPUT121), .ZN(n391) );
  AND2_X2 U431 ( .A1(n384), .A2(n492), .ZN(n688) );
  XNOR2_X1 U432 ( .A(n637), .B(KEYINPUT2), .ZN(n384) );
  XNOR2_X1 U433 ( .A(n589), .B(KEYINPUT35), .ZN(n405) );
  XNOR2_X1 U434 ( .A(n559), .B(KEYINPUT102), .ZN(n659) );
  INV_X1 U435 ( .A(n654), .ZN(n413) );
  NOR2_X1 U436 ( .A1(n615), .A2(n656), .ZN(n564) );
  XOR2_X1 U437 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n452) );
  OR2_X1 U438 ( .A1(G237), .A2(G902), .ZN(n495) );
  INV_X1 U439 ( .A(KEYINPUT69), .ZN(n441) );
  XNOR2_X1 U440 ( .A(G113), .B(G140), .ZN(n462) );
  INV_X1 U441 ( .A(G146), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n499), .B(n369), .ZN(n528) );
  XOR2_X1 U443 ( .A(KEYINPUT87), .B(KEYINPUT14), .Z(n499) );
  XNOR2_X1 U444 ( .A(n498), .B(KEYINPUT74), .ZN(n369) );
  NAND2_X1 U445 ( .A1(G234), .A2(G237), .ZN(n498) );
  NOR2_X1 U446 ( .A1(n370), .A2(n549), .ZN(n551) );
  XNOR2_X1 U447 ( .A(n430), .B(n424), .ZN(n361) );
  INV_X1 U448 ( .A(KEYINPUT84), .ZN(n624) );
  INV_X1 U449 ( .A(KEYINPUT4), .ZN(n421) );
  INV_X1 U450 ( .A(KEYINPUT17), .ZN(n380) );
  XNOR2_X1 U451 ( .A(n473), .B(n359), .ZN(n546) );
  XNOR2_X1 U452 ( .A(n474), .B(G475), .ZN(n359) );
  INV_X1 U453 ( .A(KEYINPUT6), .ZN(n385) );
  XNOR2_X1 U454 ( .A(n409), .B(n487), .ZN(n407) );
  XNOR2_X1 U455 ( .A(n488), .B(n490), .ZN(n409) );
  XNOR2_X1 U456 ( .A(n395), .B(n393), .ZN(n684) );
  XNOR2_X1 U457 ( .A(n394), .B(n479), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n477), .B(n348), .ZN(n395) );
  XNOR2_X1 U459 ( .A(n417), .B(n436), .ZN(n676) );
  XNOR2_X1 U460 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U461 ( .A(n431), .B(n418), .ZN(n417) );
  XNOR2_X1 U462 ( .A(n415), .B(KEYINPUT40), .ZN(n414) );
  INV_X1 U463 ( .A(KEYINPUT108), .ZN(n415) );
  XNOR2_X1 U464 ( .A(n375), .B(KEYINPUT36), .ZN(n534) );
  NAND2_X1 U465 ( .A1(n568), .A2(n561), .ZN(n375) );
  NOR2_X1 U466 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U467 ( .A1(n619), .A2(n363), .ZN(n597) );
  XNOR2_X1 U468 ( .A(n392), .B(n390), .ZN(n690) );
  XNOR2_X1 U469 ( .A(n689), .B(n391), .ZN(n390) );
  XNOR2_X1 U470 ( .A(n397), .B(n396), .ZN(G60) );
  INV_X1 U471 ( .A(KEYINPUT60), .ZN(n396) );
  NAND2_X1 U472 ( .A1(n398), .A2(n365), .ZN(n397) );
  XNOR2_X1 U473 ( .A(n683), .B(n682), .ZN(n398) );
  NAND2_X1 U474 ( .A1(n350), .A2(n634), .ZN(n358) );
  XNOR2_X1 U475 ( .A(n405), .B(n357), .ZN(G24) );
  INV_X1 U476 ( .A(n659), .ZN(n657) );
  AND2_X1 U477 ( .A1(n575), .A2(n574), .ZN(n627) );
  XNOR2_X1 U478 ( .A(n475), .B(KEYINPUT9), .ZN(n348) );
  XOR2_X1 U479 ( .A(G472), .B(KEYINPUT72), .Z(n349) );
  OR2_X1 U480 ( .A1(n527), .A2(n526), .ZN(n350) );
  XOR2_X1 U481 ( .A(n592), .B(KEYINPUT99), .Z(n351) );
  AND2_X1 U482 ( .A1(n623), .A2(n643), .ZN(n352) );
  XOR2_X1 U483 ( .A(n486), .B(n489), .Z(n353) );
  XNOR2_X1 U484 ( .A(KEYINPUT64), .B(KEYINPUT1), .ZN(n354) );
  XOR2_X1 U485 ( .A(n636), .B(KEYINPUT62), .Z(n355) );
  XOR2_X1 U486 ( .A(n624), .B(KEYINPUT45), .Z(n356) );
  XOR2_X1 U487 ( .A(G902), .B(KEYINPUT15), .Z(n492) );
  NOR2_X1 U488 ( .A1(G952), .A2(n706), .ZN(n691) );
  INV_X1 U489 ( .A(n691), .ZN(n365) );
  XOR2_X1 U490 ( .A(G122), .B(KEYINPUT126), .Z(n357) );
  NAND2_X1 U491 ( .A1(n389), .A2(n562), .ZN(n388) );
  NOR2_X1 U492 ( .A1(n593), .A2(n584), .ZN(n586) );
  NOR2_X2 U493 ( .A1(n510), .A2(n618), .ZN(n364) );
  OR2_X2 U494 ( .A1(n633), .A2(n358), .ZN(n376) );
  NAND2_X1 U495 ( .A1(n378), .A2(n562), .ZN(n401) );
  INV_X1 U496 ( .A(n611), .ZN(n593) );
  AND2_X1 U497 ( .A1(n611), .A2(n351), .ZN(n595) );
  INV_X1 U498 ( .A(n596), .ZN(n601) );
  NAND2_X1 U499 ( .A1(n514), .A2(n596), .ZN(n510) );
  XNOR2_X2 U500 ( .A(n553), .B(n354), .ZN(n596) );
  XNOR2_X1 U501 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U502 ( .A(n666), .B(n374), .ZN(n373) );
  XNOR2_X1 U503 ( .A(n416), .B(n414), .ZN(n715) );
  INV_X1 U504 ( .A(n598), .ZN(n621) );
  NOR2_X2 U505 ( .A1(n689), .A2(G902), .ZN(n456) );
  XNOR2_X1 U506 ( .A(n361), .B(n431), .ZN(n636) );
  NAND2_X1 U507 ( .A1(n362), .A2(n412), .ZN(n411) );
  XNOR2_X1 U508 ( .A(n560), .B(KEYINPUT46), .ZN(n362) );
  NAND2_X1 U509 ( .A1(n476), .A2(G221), .ZN(n448) );
  XNOR2_X1 U510 ( .A(n459), .B(KEYINPUT67), .ZN(n538) );
  XNOR2_X1 U511 ( .A(n364), .B(n460), .ZN(n584) );
  XNOR2_X1 U512 ( .A(n639), .B(n355), .ZN(n366) );
  NAND2_X1 U513 ( .A1(n552), .A2(n553), .ZN(n368) );
  AND2_X1 U514 ( .A1(n565), .A2(n413), .ZN(n412) );
  NOR2_X1 U515 ( .A1(n717), .A2(n405), .ZN(n404) );
  XNOR2_X1 U516 ( .A(n605), .B(KEYINPUT32), .ZN(n717) );
  XNOR2_X2 U517 ( .A(n475), .B(n421), .ZN(n482) );
  XNOR2_X2 U518 ( .A(n371), .B(G128), .ZN(n475) );
  NOR2_X2 U519 ( .A1(n411), .A2(n373), .ZN(n566) );
  XNOR2_X1 U520 ( .A(n376), .B(n635), .ZN(G75) );
  XNOR2_X2 U521 ( .A(n377), .B(n356), .ZN(n692) );
  NAND2_X1 U522 ( .A1(n402), .A2(n352), .ZN(n377) );
  INV_X1 U523 ( .A(n570), .ZN(n378) );
  XNOR2_X1 U524 ( .A(n403), .B(n606), .ZN(n402) );
  NOR2_X2 U525 ( .A1(n715), .A2(n718), .ZN(n560) );
  NAND2_X1 U526 ( .A1(n538), .A2(n553), .ZN(n609) );
  XNOR2_X1 U527 ( .A(n381), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U528 ( .A1(n673), .A2(n691), .ZN(n381) );
  NAND2_X1 U529 ( .A1(n688), .A2(G210), .ZN(n672) );
  NAND2_X1 U530 ( .A1(n346), .A2(G217), .ZN(n392) );
  NAND2_X1 U531 ( .A1(n404), .A2(n649), .ZN(n403) );
  NAND2_X1 U532 ( .A1(n567), .A2(n559), .ZN(n416) );
  XNOR2_X2 U533 ( .A(n704), .B(G146), .ZN(n431) );
  XNOR2_X1 U534 ( .A(n625), .B(KEYINPUT2), .ZN(n626) );
  XNOR2_X1 U535 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X2 U536 ( .A1(n543), .A2(n542), .ZN(n557) );
  XOR2_X1 U537 ( .A(n675), .B(n674), .Z(n419) );
  AND2_X1 U538 ( .A1(G224), .A2(n706), .ZN(n420) );
  XNOR2_X1 U539 ( .A(n483), .B(n420), .ZN(n484) );
  XNOR2_X1 U540 ( .A(KEYINPUT0), .B(KEYINPUT66), .ZN(n583) );
  XNOR2_X1 U541 ( .A(n681), .B(n680), .ZN(n682) );
  INV_X1 U542 ( .A(KEYINPUT22), .ZN(n594) );
  INV_X1 U543 ( .A(KEYINPUT63), .ZN(n640) );
  XNOR2_X1 U544 ( .A(n640), .B(KEYINPUT86), .ZN(n641) );
  XNOR2_X1 U545 ( .A(n642), .B(n641), .ZN(G57) );
  XNOR2_X1 U546 ( .A(G134), .B(KEYINPUT70), .ZN(n422) );
  XNOR2_X1 U547 ( .A(n422), .B(G131), .ZN(n423) );
  XNOR2_X2 U548 ( .A(n482), .B(n423), .ZN(n704) );
  INV_X1 U549 ( .A(n487), .ZN(n424) );
  NAND2_X1 U550 ( .A1(n464), .A2(G210), .ZN(n425) );
  XNOR2_X1 U551 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U552 ( .A(n427), .B(G119), .Z(n429) );
  XNOR2_X1 U553 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U554 ( .A(G137), .B(G140), .Z(n449) );
  XOR2_X1 U555 ( .A(KEYINPUT77), .B(n449), .Z(n433) );
  NAND2_X1 U556 ( .A1(G227), .A2(n706), .ZN(n434) );
  XNOR2_X1 U557 ( .A(KEYINPUT71), .B(G469), .ZN(n438) );
  XNOR2_X2 U558 ( .A(n439), .B(n438), .ZN(n553) );
  XNOR2_X1 U559 ( .A(n440), .B(KEYINPUT81), .ZN(n444) );
  NAND2_X1 U560 ( .A1(G234), .A2(n706), .ZN(n442) );
  XOR2_X1 U561 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n446) );
  XNOR2_X1 U562 ( .A(n488), .B(G128), .ZN(n445) );
  XNOR2_X1 U563 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U564 ( .A(n448), .B(n447), .ZN(n450) );
  XOR2_X1 U565 ( .A(n449), .B(n461), .Z(n702) );
  XNOR2_X1 U566 ( .A(n450), .B(n702), .ZN(n689) );
  INV_X1 U567 ( .A(n492), .ZN(n638) );
  NAND2_X1 U568 ( .A1(G234), .A2(n638), .ZN(n451) );
  XNOR2_X1 U569 ( .A(n452), .B(n451), .ZN(n457) );
  NAND2_X1 U570 ( .A1(n457), .A2(G217), .ZN(n454) );
  XNOR2_X2 U571 ( .A(n456), .B(n455), .ZN(n598) );
  NAND2_X1 U572 ( .A1(n457), .A2(G221), .ZN(n458) );
  XNOR2_X1 U573 ( .A(n458), .B(KEYINPUT21), .ZN(n591) );
  INV_X1 U574 ( .A(n591), .ZN(n511) );
  NAND2_X1 U575 ( .A1(n621), .A2(n511), .ZN(n459) );
  BUF_X1 U576 ( .A(n538), .Z(n514) );
  XNOR2_X1 U577 ( .A(KEYINPUT100), .B(KEYINPUT33), .ZN(n460) );
  XNOR2_X1 U578 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n474) );
  XOR2_X1 U579 ( .A(n461), .B(n486), .Z(n472) );
  XNOR2_X1 U580 ( .A(n463), .B(n462), .ZN(n468) );
  NAND2_X1 U581 ( .A1(G214), .A2(n464), .ZN(n465) );
  XNOR2_X1 U582 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U583 ( .A(n468), .B(n467), .ZN(n470) );
  XNOR2_X1 U584 ( .A(G143), .B(G131), .ZN(n469) );
  NOR2_X1 U585 ( .A1(G902), .A2(n681), .ZN(n473) );
  INV_X1 U586 ( .A(n546), .ZN(n481) );
  NAND2_X1 U587 ( .A1(G217), .A2(n476), .ZN(n477) );
  XOR2_X1 U588 ( .A(KEYINPUT97), .B(KEYINPUT7), .Z(n479) );
  NOR2_X1 U589 ( .A1(n684), .A2(G902), .ZN(n480) );
  NAND2_X1 U590 ( .A1(n481), .A2(n544), .ZN(n590) );
  XNOR2_X1 U591 ( .A(n485), .B(KEYINPUT18), .ZN(n491) );
  AND2_X1 U592 ( .A1(G210), .A2(n495), .ZN(n493) );
  XNOR2_X1 U593 ( .A(KEYINPUT38), .B(n570), .ZN(n556) );
  NAND2_X1 U594 ( .A1(G214), .A2(n495), .ZN(n562) );
  NAND2_X1 U595 ( .A1(n556), .A2(n562), .ZN(n505) );
  NOR2_X1 U596 ( .A1(n590), .A2(n505), .ZN(n496) );
  XNOR2_X1 U597 ( .A(n496), .B(KEYINPUT41), .ZN(n554) );
  NOR2_X1 U598 ( .A1(n584), .A2(n554), .ZN(n497) );
  NOR2_X1 U599 ( .A1(G953), .A2(n497), .ZN(n634) );
  NAND2_X1 U600 ( .A1(n528), .A2(G952), .ZN(n500) );
  XNOR2_X1 U601 ( .A(n500), .B(KEYINPUT88), .ZN(n527) );
  NOR2_X1 U602 ( .A1(n556), .A2(n562), .ZN(n501) );
  XOR2_X1 U603 ( .A(KEYINPUT115), .B(n501), .Z(n502) );
  NOR2_X1 U604 ( .A1(n590), .A2(n502), .ZN(n503) );
  XNOR2_X1 U605 ( .A(n503), .B(KEYINPUT116), .ZN(n507) );
  NOR2_X1 U606 ( .A1(n544), .A2(n546), .ZN(n662) );
  NOR2_X1 U607 ( .A1(n662), .A2(n559), .ZN(n615) );
  NOR2_X1 U608 ( .A1(n505), .A2(n615), .ZN(n506) );
  NOR2_X1 U609 ( .A1(n507), .A2(n506), .ZN(n508) );
  XOR2_X1 U610 ( .A(KEYINPUT117), .B(n508), .Z(n509) );
  NOR2_X1 U611 ( .A1(n584), .A2(n509), .ZN(n524) );
  NOR2_X1 U612 ( .A1(n370), .A2(n510), .ZN(n610) );
  NOR2_X1 U613 ( .A1(n511), .A2(n363), .ZN(n512) );
  XNOR2_X1 U614 ( .A(n512), .B(KEYINPUT49), .ZN(n513) );
  NAND2_X1 U615 ( .A1(n370), .A2(n513), .ZN(n517) );
  NOR2_X1 U616 ( .A1(n596), .A2(n514), .ZN(n515) );
  XNOR2_X1 U617 ( .A(n515), .B(KEYINPUT50), .ZN(n516) );
  NOR2_X1 U618 ( .A1(n517), .A2(n516), .ZN(n518) );
  XOR2_X1 U619 ( .A(KEYINPUT113), .B(n518), .Z(n519) );
  NOR2_X1 U620 ( .A1(n610), .A2(n519), .ZN(n520) );
  XOR2_X1 U621 ( .A(KEYINPUT51), .B(n520), .Z(n521) );
  NOR2_X1 U622 ( .A1(n554), .A2(n521), .ZN(n522) );
  XNOR2_X1 U623 ( .A(n522), .B(KEYINPUT114), .ZN(n523) );
  NOR2_X1 U624 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U625 ( .A(n525), .B(KEYINPUT52), .ZN(n526) );
  INV_X1 U626 ( .A(n372), .ZN(n561) );
  NOR2_X1 U627 ( .A1(G953), .A2(n527), .ZN(n576) );
  NAND2_X1 U628 ( .A1(n528), .A2(G902), .ZN(n529) );
  XNOR2_X1 U629 ( .A(n529), .B(KEYINPUT89), .ZN(n577) );
  NAND2_X1 U630 ( .A1(G953), .A2(n577), .ZN(n530) );
  NOR2_X1 U631 ( .A1(G900), .A2(n530), .ZN(n531) );
  XOR2_X1 U632 ( .A(KEYINPUT103), .B(n531), .Z(n532) );
  NOR2_X1 U633 ( .A1(n576), .A2(n532), .ZN(n539) );
  NOR2_X1 U634 ( .A1(n539), .A2(n591), .ZN(n533) );
  NAND2_X1 U635 ( .A1(n598), .A2(n533), .ZN(n549) );
  NOR2_X1 U636 ( .A1(n601), .A2(n534), .ZN(n666) );
  INV_X1 U637 ( .A(n607), .ZN(n535) );
  NAND2_X1 U638 ( .A1(n562), .A2(n535), .ZN(n537) );
  XOR2_X1 U639 ( .A(KEYINPUT105), .B(KEYINPUT30), .Z(n536) );
  XNOR2_X1 U640 ( .A(n537), .B(n536), .ZN(n543) );
  NOR2_X2 U641 ( .A1(n609), .A2(n539), .ZN(n541) );
  INV_X1 U642 ( .A(KEYINPUT76), .ZN(n540) );
  XNOR2_X1 U643 ( .A(n541), .B(n540), .ZN(n542) );
  INV_X1 U644 ( .A(n544), .ZN(n545) );
  NAND2_X1 U645 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U646 ( .A(n547), .B(KEYINPUT101), .ZN(n587) );
  NAND2_X1 U647 ( .A1(n557), .A2(n587), .ZN(n548) );
  NOR2_X1 U648 ( .A1(n372), .A2(n548), .ZN(n654) );
  XNOR2_X1 U649 ( .A(KEYINPUT28), .B(KEYINPUT106), .ZN(n550) );
  XNOR2_X1 U650 ( .A(n551), .B(n550), .ZN(n552) );
  NOR2_X1 U651 ( .A1(n563), .A2(n554), .ZN(n555) );
  XNOR2_X1 U652 ( .A(n555), .B(KEYINPUT42), .ZN(n718) );
  NAND2_X1 U653 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U654 ( .A(n558), .B(KEYINPUT39), .ZN(n567) );
  OR2_X1 U655 ( .A1(n563), .A2(n582), .ZN(n656) );
  XNOR2_X1 U656 ( .A(n564), .B(KEYINPUT47), .ZN(n565) );
  XNOR2_X1 U657 ( .A(n566), .B(KEYINPUT48), .ZN(n575) );
  NAND2_X1 U658 ( .A1(n567), .A2(n662), .ZN(n668) );
  NAND2_X1 U659 ( .A1(n568), .A2(n601), .ZN(n569) );
  XNOR2_X1 U660 ( .A(n569), .B(KEYINPUT43), .ZN(n571) );
  NAND2_X1 U661 ( .A1(n571), .A2(n372), .ZN(n572) );
  XOR2_X1 U662 ( .A(KEYINPUT104), .B(n572), .Z(n716) );
  INV_X1 U663 ( .A(n716), .ZN(n573) );
  AND2_X1 U664 ( .A1(n668), .A2(n573), .ZN(n574) );
  INV_X1 U665 ( .A(n576), .ZN(n579) );
  NOR2_X1 U666 ( .A1(G898), .A2(n706), .ZN(n699) );
  NAND2_X1 U667 ( .A1(n577), .A2(n699), .ZN(n578) );
  NAND2_X1 U668 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U669 ( .A(KEYINPUT90), .B(n580), .Z(n581) );
  XNOR2_X1 U670 ( .A(KEYINPUT34), .B(KEYINPUT78), .ZN(n585) );
  XNOR2_X1 U671 ( .A(n586), .B(n585), .ZN(n588) );
  NAND2_X1 U672 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U673 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U674 ( .A(n595), .B(n594), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n370), .A2(n597), .ZN(n649) );
  XNOR2_X1 U676 ( .A(n618), .B(KEYINPUT80), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U678 ( .A(n602), .B(KEYINPUT79), .ZN(n603) );
  NOR2_X1 U679 ( .A1(n604), .A2(n603), .ZN(n605) );
  INV_X1 U680 ( .A(KEYINPUT44), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n370), .A2(n347), .ZN(n608) );
  NOR2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n645) );
  NAND2_X1 U683 ( .A1(n347), .A2(n610), .ZN(n613) );
  XNOR2_X1 U684 ( .A(KEYINPUT31), .B(KEYINPUT92), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n613), .B(n612), .ZN(n663) );
  NOR2_X1 U686 ( .A1(n645), .A2(n663), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n614), .B(KEYINPUT93), .ZN(n617) );
  INV_X1 U688 ( .A(n615), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n623) );
  INV_X1 U690 ( .A(n618), .ZN(n620) );
  NOR2_X1 U691 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U692 ( .A1(n622), .A2(n363), .ZN(n643) );
  NAND2_X1 U693 ( .A1(n637), .A2(KEYINPUT82), .ZN(n625) );
  INV_X1 U694 ( .A(n626), .ZN(n631) );
  INV_X1 U695 ( .A(KEYINPUT82), .ZN(n629) );
  INV_X1 U696 ( .A(n627), .ZN(n705) );
  NAND2_X1 U697 ( .A1(n705), .A2(n692), .ZN(n628) );
  NAND2_X1 U698 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U699 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U700 ( .A(KEYINPUT83), .B(n632), .ZN(n633) );
  INV_X1 U701 ( .A(KEYINPUT53), .ZN(n635) );
  NAND2_X1 U702 ( .A1(n688), .A2(G472), .ZN(n639) );
  XNOR2_X1 U703 ( .A(G101), .B(n643), .ZN(G3) );
  NAND2_X1 U704 ( .A1(n645), .A2(n659), .ZN(n644) );
  XNOR2_X1 U705 ( .A(n644), .B(G104), .ZN(G6) );
  XOR2_X1 U706 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n647) );
  NAND2_X1 U707 ( .A1(n645), .A2(n662), .ZN(n646) );
  XNOR2_X1 U708 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U709 ( .A(G107), .B(n648), .ZN(G9) );
  XNOR2_X1 U710 ( .A(G110), .B(n649), .ZN(G12) );
  INV_X1 U711 ( .A(n662), .ZN(n650) );
  NOR2_X1 U712 ( .A1(n650), .A2(n656), .ZN(n652) );
  XNOR2_X1 U713 ( .A(KEYINPUT109), .B(KEYINPUT29), .ZN(n651) );
  XNOR2_X1 U714 ( .A(n652), .B(n651), .ZN(n653) );
  XOR2_X1 U715 ( .A(G128), .B(n653), .Z(G30) );
  XOR2_X1 U716 ( .A(G143), .B(n654), .Z(n655) );
  XNOR2_X1 U717 ( .A(KEYINPUT110), .B(n655), .ZN(G45) );
  NOR2_X1 U718 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U719 ( .A(G146), .B(n658), .Z(G48) );
  XOR2_X1 U720 ( .A(G113), .B(KEYINPUT111), .Z(n661) );
  NAND2_X1 U721 ( .A1(n659), .A2(n663), .ZN(n660) );
  XNOR2_X1 U722 ( .A(n661), .B(n660), .ZN(G15) );
  NAND2_X1 U723 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U724 ( .A(n664), .B(KEYINPUT112), .ZN(n665) );
  XNOR2_X1 U725 ( .A(G116), .B(n665), .ZN(G18) );
  XNOR2_X1 U726 ( .A(G125), .B(n666), .ZN(n667) );
  XNOR2_X1 U727 ( .A(n667), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U728 ( .A(G134), .B(n668), .ZN(G36) );
  XOR2_X1 U729 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n669) );
  NAND2_X1 U730 ( .A1(n346), .A2(G469), .ZN(n678) );
  XOR2_X1 U731 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n675) );
  XNOR2_X1 U732 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n674) );
  XNOR2_X1 U733 ( .A(n676), .B(n419), .ZN(n677) );
  XNOR2_X1 U734 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X1 U735 ( .A1(n691), .A2(n679), .ZN(G54) );
  NAND2_X1 U736 ( .A1(n688), .A2(G475), .ZN(n683) );
  XOR2_X1 U737 ( .A(KEYINPUT59), .B(KEYINPUT65), .Z(n680) );
  XNOR2_X1 U738 ( .A(n684), .B(KEYINPUT120), .ZN(n686) );
  NAND2_X1 U739 ( .A1(G478), .A2(n688), .ZN(n685) );
  XNOR2_X1 U740 ( .A(n686), .B(n685), .ZN(n687) );
  NOR2_X1 U741 ( .A1(n691), .A2(n687), .ZN(G63) );
  NOR2_X1 U742 ( .A1(n691), .A2(n690), .ZN(G66) );
  NAND2_X1 U743 ( .A1(n706), .A2(n692), .ZN(n696) );
  NAND2_X1 U744 ( .A1(G953), .A2(G224), .ZN(n693) );
  XNOR2_X1 U745 ( .A(KEYINPUT61), .B(n693), .ZN(n694) );
  NAND2_X1 U746 ( .A1(n694), .A2(G898), .ZN(n695) );
  NAND2_X1 U747 ( .A1(n696), .A2(n695), .ZN(n701) );
  XOR2_X1 U748 ( .A(n697), .B(KEYINPUT122), .Z(n698) );
  NOR2_X1 U749 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U750 ( .A(n701), .B(n700), .ZN(G69) );
  XOR2_X1 U751 ( .A(n702), .B(KEYINPUT123), .Z(n703) );
  XOR2_X1 U752 ( .A(n704), .B(n703), .Z(n708) );
  XNOR2_X1 U753 ( .A(n705), .B(n708), .ZN(n707) );
  NAND2_X1 U754 ( .A1(n707), .A2(n706), .ZN(n714) );
  XNOR2_X1 U755 ( .A(KEYINPUT124), .B(n708), .ZN(n709) );
  XNOR2_X1 U756 ( .A(G227), .B(n709), .ZN(n710) );
  NAND2_X1 U757 ( .A1(G900), .A2(n710), .ZN(n711) );
  XOR2_X1 U758 ( .A(KEYINPUT125), .B(n711), .Z(n712) );
  NAND2_X1 U759 ( .A1(G953), .A2(n712), .ZN(n713) );
  NAND2_X1 U760 ( .A1(n714), .A2(n713), .ZN(G72) );
  XOR2_X1 U761 ( .A(G131), .B(n715), .Z(G33) );
  XOR2_X1 U762 ( .A(G140), .B(n716), .Z(G42) );
  XOR2_X1 U763 ( .A(G119), .B(n717), .Z(G21) );
  XOR2_X1 U764 ( .A(G137), .B(n718), .Z(G39) );
endmodule

