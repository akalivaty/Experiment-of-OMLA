//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1221, new_n1222, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT65), .B(G77), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G58), .A2(G232), .ZN(new_n227));
  NAND4_X1  g0027(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n211), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n214), .B1(new_n218), .B2(new_n219), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT68), .ZN(new_n248));
  AND2_X1   g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n248), .B1(new_n249), .B2(new_n215), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n251), .A2(KEYINPUT68), .A3(G1), .A4(G13), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(G274), .A3(new_n252), .ZN(new_n253));
  OR2_X1    g0053(.A1(KEYINPUT67), .A2(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT67), .A2(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OR2_X1    g0059(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G226), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n250), .A2(new_n252), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G223), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n267), .A2(new_n268), .B1(new_n221), .B2(new_n266), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1698), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n269), .B1(G222), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n249), .A2(new_n215), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n260), .B1(new_n261), .B2(new_n265), .C1(new_n274), .C2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G190), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n279), .B1(G200), .B2(new_n277), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT9), .ZN(new_n281));
  INV_X1    g0081(.A(G13), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G1), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G20), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT71), .ZN(new_n286));
  NAND4_X1  g0086(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n287), .A2(new_n215), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT69), .ZN(new_n289));
  INV_X1    g0089(.A(G33), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n289), .B1(new_n211), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(KEYINPUT70), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  AND4_X1   g0092(.A1(KEYINPUT70), .A2(new_n291), .A3(new_n215), .A4(new_n287), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n286), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(new_n215), .A3(new_n287), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT70), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n288), .A2(KEYINPUT70), .A3(new_n291), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT71), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n285), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n300), .B(G50), .C1(G1), .C2(new_n216), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n285), .A2(new_n202), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT72), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n301), .A2(KEYINPUT72), .A3(new_n302), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n294), .A2(new_n299), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n204), .A2(new_n216), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT8), .B(G58), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n216), .A2(G33), .ZN(new_n312));
  INV_X1    g0112(.A(G150), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n216), .A2(new_n290), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n311), .A2(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n309), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n281), .B1(new_n307), .B2(new_n316), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n301), .A2(KEYINPUT72), .A3(new_n302), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT72), .B1(new_n301), .B2(new_n302), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n281), .B(new_n316), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n280), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT10), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT9), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n320), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT10), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(new_n280), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT13), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n261), .A2(G1698), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n270), .B2(new_n271), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT74), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n266), .A2(KEYINPUT74), .A3(new_n331), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g0136(.A(G232), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n337), .A2(KEYINPUT75), .B1(G33), .B2(G97), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT75), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n266), .A2(new_n339), .A3(G232), .A4(G1698), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n336), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n275), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n250), .A2(G238), .A3(new_n252), .A4(new_n264), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n253), .B2(new_n259), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n330), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  AOI211_X1 g0146(.A(KEYINPUT13), .B(new_n344), .C1(new_n341), .C2(new_n275), .ZN(new_n347));
  OAI21_X1  g0147(.A(G169), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(KEYINPUT14), .ZN(new_n349));
  INV_X1    g0149(.A(G179), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n346), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n348), .A2(KEYINPUT78), .A3(KEYINPUT14), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT78), .B1(new_n348), .B2(KEYINPUT14), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G68), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G20), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n358), .B1(new_n312), .B2(new_n205), .C1(new_n202), .C2(new_n314), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n294), .A2(new_n299), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT11), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n294), .A2(KEYINPUT11), .A3(new_n299), .A4(new_n359), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n284), .A2(G68), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT12), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n285), .B1(new_n297), .B2(new_n298), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n216), .A2(G1), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n367), .A2(new_n357), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n365), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n362), .A2(new_n363), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n356), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n277), .A2(G179), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT73), .ZN(new_n373));
  INV_X1    g0173(.A(G169), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n277), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n324), .A3(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n260), .B1(new_n265), .B2(new_n222), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n273), .A2(G232), .ZN(new_n378));
  INV_X1    g0178(.A(G238), .ZN(new_n379));
  OAI221_X1 g0179(.A(new_n378), .B1(new_n208), .B2(new_n266), .C1(new_n379), .C2(new_n267), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n377), .B1(new_n275), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G190), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n292), .A2(new_n293), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n220), .A2(G20), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT15), .B(G87), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n384), .B1(new_n312), .B2(new_n385), .C1(new_n311), .C2(new_n314), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n220), .B2(new_n284), .ZN(new_n388));
  NOR4_X1   g0188(.A1(new_n383), .A2(new_n205), .A3(new_n285), .A4(new_n367), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G200), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n382), .B(new_n390), .C1(new_n391), .C2(new_n381), .ZN(new_n392));
  INV_X1    g0192(.A(new_n390), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n381), .A2(new_n350), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n393), .B(new_n394), .C1(G169), .C2(new_n381), .ZN(new_n395));
  AND4_X1   g0195(.A1(new_n371), .A2(new_n376), .A3(new_n392), .A4(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n311), .A2(new_n367), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n300), .A2(new_n397), .B1(new_n311), .B2(new_n285), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n266), .B2(G20), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n216), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n357), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  INV_X1    g0203(.A(G58), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(new_n357), .ZN(new_n405));
  OAI21_X1  g0205(.A(G20), .B1(new_n405), .B2(new_n201), .ZN(new_n406));
  INV_X1    g0206(.A(G159), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n406), .B1(new_n407), .B2(new_n314), .ZN(new_n408));
  OR3_X1    g0208(.A1(new_n402), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n403), .B1(new_n402), .B2(new_n408), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n383), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n398), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT79), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT80), .ZN(new_n415));
  INV_X1    g0215(.A(G1698), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n272), .A2(new_n416), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n273), .A2(G223), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n276), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n250), .A2(G232), .A3(new_n252), .A4(new_n264), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n253), .B2(new_n259), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n420), .A2(new_n350), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n266), .A2(G226), .A3(G1698), .ZN(new_n424));
  INV_X1    g0224(.A(G87), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n266), .A2(new_n416), .ZN(new_n426));
  OAI221_X1 g0226(.A(new_n424), .B1(new_n290), .B2(new_n425), .C1(new_n426), .C2(new_n268), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n275), .ZN(new_n428));
  INV_X1    g0228(.A(new_n422), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n374), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n415), .B1(new_n423), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(G169), .B1(new_n420), .B2(new_n422), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(G179), .A3(new_n429), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT80), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n398), .A2(KEYINPUT79), .A3(new_n411), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n414), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT18), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  OAI21_X1  g0239(.A(G200), .B1(new_n420), .B2(new_n422), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n428), .A2(G190), .A3(new_n429), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n439), .B1(new_n412), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n442), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n444), .A2(KEYINPUT17), .A3(new_n411), .A4(new_n398), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT18), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n414), .A2(new_n435), .A3(new_n447), .A4(new_n436), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n438), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT77), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT76), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n391), .B1(new_n346), .B2(new_n347), .ZN(new_n453));
  INV_X1    g0253(.A(new_n337), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n334), .A2(new_n335), .B1(new_n454), .B2(new_n339), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n276), .B1(new_n455), .B2(new_n338), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT13), .B1(new_n456), .B2(new_n344), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n342), .A2(new_n330), .A3(new_n345), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n278), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n370), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n452), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI211_X1 g0262(.A(KEYINPUT76), .B(new_n370), .C1(new_n453), .C2(new_n459), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n451), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n346), .A2(new_n347), .A3(G190), .ZN(new_n465));
  AOI21_X1  g0265(.A(G200), .B1(new_n457), .B2(new_n458), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT76), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n460), .A2(new_n452), .A3(new_n461), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(KEYINPUT77), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  AND4_X1   g0271(.A1(new_n329), .A2(new_n396), .A3(new_n450), .A4(new_n471), .ZN(new_n472));
  XNOR2_X1  g0272(.A(G97), .B(G107), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT81), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(KEYINPUT6), .ZN(new_n475));
  MUX2_X1   g0275(.A(new_n474), .B(G97), .S(KEYINPUT6), .Z(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n477), .A2(new_n216), .B1(new_n205), .B2(new_n314), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n208), .B1(new_n400), .B2(new_n401), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n383), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n285), .A2(new_n207), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n290), .A2(G1), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n300), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n482), .B1(new_n486), .B2(G97), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT5), .B1(new_n254), .B2(new_n256), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT5), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n258), .B(G45), .C1(new_n489), .C2(G41), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n253), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n254), .A2(new_n256), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n490), .B1(new_n492), .B2(new_n489), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(new_n262), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n491), .B1(G257), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n417), .A2(G250), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n266), .A2(G244), .A3(new_n416), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .A4(new_n416), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G283), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n496), .A2(new_n499), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n275), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n495), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT83), .B1(new_n504), .B2(new_n278), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT83), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n495), .A2(new_n503), .A3(new_n506), .A4(G190), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n502), .A2(KEYINPUT82), .A3(new_n275), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT82), .B1(new_n502), .B2(new_n275), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n495), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G200), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n487), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n300), .A2(G87), .A3(new_n484), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n266), .A2(new_n216), .A3(G68), .ZN(new_n515));
  NAND3_X1  g0315(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n216), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(G87), .B2(new_n209), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n312), .A2(new_n207), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n515), .B(new_n518), .C1(KEYINPUT19), .C2(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n383), .A2(new_n520), .B1(new_n285), .B2(new_n385), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n266), .A2(G244), .A3(G1698), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G116), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n523), .B(new_n524), .C1(new_n426), .C2(new_n379), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n275), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n258), .A2(G45), .ZN(new_n527));
  INV_X1    g0327(.A(G250), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n263), .B(new_n529), .C1(G274), .C2(new_n527), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G190), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n526), .A2(new_n530), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G200), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n521), .B1(new_n485), .B2(new_n385), .ZN(new_n536));
  AOI21_X1  g0336(.A(G169), .B1(new_n526), .B2(new_n530), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n350), .B2(new_n531), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n522), .A2(new_n535), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n481), .B(new_n480), .C1(new_n485), .C2(new_n207), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n504), .A2(new_n374), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n350), .B(new_n495), .C1(new_n509), .C2(new_n510), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n513), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n494), .A2(G270), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT84), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n263), .A2(G274), .A3(new_n493), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(G270), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n493), .A2(new_n262), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT84), .B1(new_n550), .B2(new_n491), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n417), .A2(G264), .ZN(new_n553));
  INV_X1    g0353(.A(G257), .ZN(new_n554));
  INV_X1    g0354(.A(G303), .ZN(new_n555));
  OAI221_X1 g0355(.A(new_n553), .B1(new_n554), .B2(new_n426), .C1(new_n555), .C2(new_n266), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n275), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(G20), .B1(new_n290), .B2(G97), .ZN(new_n559));
  INV_X1    g0359(.A(G116), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n559), .A2(new_n501), .B1(G20), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n295), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g0362(.A(new_n562), .B(KEYINPUT20), .Z(new_n563));
  NAND3_X1  g0363(.A1(new_n366), .A2(G116), .A3(new_n484), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n284), .A2(G116), .ZN(new_n565));
  XNOR2_X1  g0365(.A(new_n565), .B(KEYINPUT85), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n558), .A2(KEYINPUT21), .A3(G169), .A4(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n548), .A2(new_n551), .B1(new_n275), .B2(new_n556), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n567), .A3(G179), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n558), .A2(G169), .A3(new_n567), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n567), .B1(new_n558), .B2(G200), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n278), .B2(new_n558), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n571), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n266), .A2(new_n216), .A3(G87), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n578), .B(KEYINPUT22), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT24), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT23), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n216), .B2(G107), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n208), .A2(KEYINPUT23), .A3(G20), .ZN(new_n583));
  INV_X1    g0383(.A(new_n524), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n582), .A2(new_n583), .B1(new_n584), .B2(new_n216), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n579), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n580), .B1(new_n579), .B2(new_n585), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n383), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n300), .A2(G107), .A3(new_n484), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n285), .A2(KEYINPUT25), .A3(new_n208), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT86), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT25), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n284), .B2(G107), .ZN(new_n594));
  XOR2_X1   g0394(.A(new_n592), .B(new_n594), .Z(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n589), .A2(new_n590), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n494), .A2(G264), .ZN(new_n598));
  INV_X1    g0398(.A(G294), .ZN(new_n599));
  OAI22_X1  g0399(.A1(new_n426), .A2(new_n528), .B1(new_n290), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT87), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n417), .A2(new_n601), .A3(G257), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT87), .B1(new_n267), .B2(new_n554), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n547), .B(new_n598), .C1(new_n604), .C2(new_n276), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT88), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n606), .A3(G169), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n350), .B2(new_n605), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n606), .B1(new_n605), .B2(G169), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n597), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n579), .A2(new_n585), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT24), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n586), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n595), .B1(new_n613), .B2(new_n383), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n273), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n601), .B1(new_n417), .B2(G257), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n267), .A2(KEYINPUT87), .A3(new_n554), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n618), .A2(new_n275), .B1(G264), .B2(new_n494), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(G190), .A3(new_n547), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n605), .A2(G200), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n614), .A2(new_n590), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n610), .A2(new_n622), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n472), .A2(new_n544), .A3(new_n577), .A4(new_n623), .ZN(G372));
  INV_X1    g0424(.A(new_n376), .ZN(new_n625));
  INV_X1    g0425(.A(new_n371), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n395), .B1(new_n468), .B2(new_n469), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n446), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n432), .A2(new_n433), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n412), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n630), .B(KEYINPUT18), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n625), .B1(new_n633), .B2(new_n329), .ZN(new_n634));
  INV_X1    g0434(.A(new_n472), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n543), .A2(new_n513), .A3(new_n539), .A4(new_n622), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n610), .A2(new_n571), .A3(new_n574), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n536), .A2(new_n538), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT89), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n543), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n540), .A2(KEYINPUT89), .A3(new_n541), .A4(new_n542), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n642), .A2(new_n643), .A3(new_n539), .A4(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n514), .A2(new_n532), .A3(new_n521), .A4(new_n534), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT26), .B1(new_n647), .B2(new_n543), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n640), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n634), .B1(new_n635), .B2(new_n650), .ZN(G369));
  NAND2_X1  g0451(.A1(new_n283), .A2(new_n216), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  XOR2_X1   g0453(.A(new_n653), .B(KEYINPUT90), .Z(new_n654));
  INV_X1    g0454(.A(G213), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n652), .B2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n567), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n577), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n571), .A2(new_n574), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(new_n660), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G330), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n597), .A2(new_n659), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n623), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n659), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n667), .B1(new_n610), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n610), .A2(new_n659), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n662), .A2(new_n659), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n623), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n212), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(new_n492), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n209), .A2(G87), .A3(G116), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G1), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n219), .B2(new_n677), .ZN(new_n680));
  XOR2_X1   g0480(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n681));
  XNOR2_X1  g0481(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n577), .A2(new_n623), .A3(new_n544), .A4(new_n668), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n569), .A2(G179), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n619), .A2(new_n503), .A3(new_n495), .A4(new_n531), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT92), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT30), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  OAI211_X1 g0488(.A(KEYINPUT92), .B(new_n688), .C1(new_n684), .C2(new_n685), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n569), .A2(G179), .A3(new_n531), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(new_n511), .A3(new_n605), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n687), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT31), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n692), .A2(new_n693), .A3(new_n659), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n693), .B1(new_n692), .B2(new_n659), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n683), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G330), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n668), .B1(new_n640), .B2(new_n649), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT93), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n636), .A2(new_n637), .B1(new_n536), .B2(new_n538), .ZN(new_n704));
  INV_X1    g0504(.A(new_n649), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n659), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(KEYINPUT93), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n702), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n642), .A2(KEYINPUT26), .A3(new_n539), .A4(new_n644), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n643), .B1(new_n647), .B2(new_n543), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(KEYINPUT94), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n647), .B1(new_n641), .B2(new_n543), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT94), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n712), .A2(new_n713), .A3(KEYINPUT26), .A4(new_n644), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n638), .A2(new_n711), .A3(new_n714), .A4(new_n639), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(KEYINPUT29), .A3(new_n668), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n699), .B1(new_n708), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n682), .B1(new_n717), .B2(G1), .ZN(G364));
  NOR2_X1   g0518(.A1(new_n282), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n258), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n676), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n665), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(G330), .B2(new_n663), .ZN(new_n724));
  INV_X1    g0524(.A(new_n722), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n215), .B1(G20), .B2(new_n374), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n216), .A2(G179), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(new_n278), .A3(G200), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n208), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(G190), .A3(G200), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n730), .B1(G87), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n216), .A2(new_n350), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G200), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G190), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n733), .B1(new_n357), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(G190), .A3(new_n391), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n735), .A2(new_n278), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI221_X1 g0541(.A(new_n266), .B1(new_n404), .B2(new_n739), .C1(new_n741), .C2(new_n202), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n216), .A2(G190), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n744), .A2(new_n350), .A3(G200), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n746), .A2(KEYINPUT96), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(KEYINPUT96), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n738), .B(new_n742), .C1(new_n750), .C2(new_n220), .ZN(new_n751));
  OR3_X1    g0551(.A1(KEYINPUT97), .A2(G179), .A3(G200), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT97), .B1(G179), .B2(G200), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n278), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n216), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G97), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n744), .B1(new_n752), .B2(new_n753), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(KEYINPUT32), .B1(new_n759), .B2(new_n407), .ZN(new_n760));
  OR3_X1    g0560(.A1(new_n759), .A2(KEYINPUT32), .A3(new_n407), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n751), .A2(new_n757), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G283), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n729), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g0564(.A(KEYINPUT33), .B(G317), .Z(new_n765));
  OAI22_X1  g0565(.A1(new_n737), .A2(new_n765), .B1(new_n731), .B2(new_n555), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n764), .B(new_n766), .C1(G326), .C2(new_n740), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n756), .A2(G294), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n758), .A2(G329), .ZN(new_n769));
  INV_X1    g0569(.A(G322), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n272), .B1(new_n739), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(G311), .B2(new_n745), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n767), .A2(new_n768), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n727), .B1(new_n762), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n726), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n675), .A2(new_n272), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT95), .ZN(new_n780));
  INV_X1    g0580(.A(G355), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n780), .A2(new_n781), .B1(G116), .B2(new_n212), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n675), .A2(new_n266), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(G45), .B2(new_n219), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(G45), .B2(new_n246), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n725), .B(new_n774), .C1(new_n778), .C2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n777), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n663), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n724), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(G396));
  NAND2_X1  g0591(.A1(new_n393), .A2(new_n659), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT100), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(KEYINPUT100), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n793), .A2(new_n392), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n395), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n395), .A2(new_n659), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n702), .A2(new_n707), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(KEYINPUT101), .ZN(new_n800));
  INV_X1    g0600(.A(new_n798), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n706), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT101), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n702), .A2(new_n707), .A3(new_n803), .A4(new_n798), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n800), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n699), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n722), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n806), .B2(new_n805), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n726), .A2(new_n775), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n725), .B1(new_n205), .B2(new_n809), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n272), .B1(new_n599), .B2(new_n739), .C1(new_n741), .C2(new_n555), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n749), .A2(new_n560), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n811), .B(new_n812), .C1(G311), .C2(new_n758), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n732), .A2(G107), .ZN(new_n814));
  INV_X1    g0614(.A(new_n729), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n736), .A2(G283), .B1(new_n815), .B2(G87), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n813), .A2(new_n757), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT98), .Z(new_n818));
  NOR2_X1   g0618(.A1(new_n729), .A2(new_n357), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n272), .B(new_n819), .C1(G50), .C2(new_n732), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n758), .A2(G132), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(new_n404), .C2(new_n755), .ZN(new_n822));
  INV_X1    g0622(.A(new_n739), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G137), .A2(new_n740), .B1(new_n823), .B2(G143), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n313), .B2(new_n737), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n750), .B2(G159), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n822), .B1(new_n826), .B2(KEYINPUT34), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(KEYINPUT34), .B2(new_n826), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n818), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(KEYINPUT99), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n726), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n829), .A2(KEYINPUT99), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n810), .B1(new_n776), .B2(new_n801), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n808), .A2(new_n833), .ZN(G384));
  INV_X1    g0634(.A(KEYINPUT35), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n560), .B(new_n218), .C1(new_n477), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n477), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n836), .A2(KEYINPUT102), .B1(KEYINPUT35), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(KEYINPUT102), .B2(new_n836), .ZN(new_n839));
  XNOR2_X1  g0639(.A(KEYINPUT103), .B(KEYINPUT36), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n839), .B(new_n840), .ZN(new_n841));
  OR3_X1    g0641(.A1(new_n221), .A2(new_n219), .A3(new_n405), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n202), .A2(G68), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n258), .B(G13), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n472), .A2(new_n699), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n461), .A2(new_n668), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n462), .B2(new_n463), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n626), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT104), .ZN(new_n852));
  INV_X1    g0652(.A(new_n356), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n462), .A2(new_n463), .A3(new_n451), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT77), .B1(new_n468), .B2(new_n469), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n852), .B1(new_n856), .B2(new_n847), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n356), .B1(new_n464), .B2(new_n470), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n858), .A2(KEYINPUT104), .A3(new_n848), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n851), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n657), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n309), .A2(new_n410), .A3(new_n409), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n300), .A2(new_n397), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n285), .A2(new_n311), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n861), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n449), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n657), .B(KEYINPUT105), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n414), .A2(new_n436), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n412), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT37), .B1(new_n871), .B2(new_n444), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n437), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n629), .B1(new_n862), .B2(new_n865), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n444), .A2(new_n411), .A3(new_n398), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n866), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n878), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n414), .A2(new_n436), .A3(new_n869), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n875), .A2(new_n630), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n873), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n443), .A2(new_n445), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n880), .B1(new_n631), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n879), .B1(new_n886), .B2(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n696), .A2(new_n801), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n860), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n856), .A2(new_n852), .A3(new_n847), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT104), .B1(new_n858), .B2(new_n848), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n888), .B1(new_n893), .B2(new_n851), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n868), .A2(new_n878), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT40), .B1(new_n897), .B2(new_n879), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n890), .A2(KEYINPUT40), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n846), .B1(new_n899), .B2(new_n698), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT106), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n899), .A2(new_n635), .A3(new_n697), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n802), .A2(new_n797), .B1(new_n893), .B2(new_n851), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n897), .A2(new_n879), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n887), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n626), .A2(new_n668), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n908), .B(new_n910), .C1(new_n905), .C2(new_n907), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n632), .A2(new_n869), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n906), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n708), .A2(new_n472), .A3(new_n716), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n634), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n913), .B(new_n915), .Z(new_n916));
  OAI22_X1  g0716(.A1(new_n903), .A2(new_n916), .B1(new_n258), .B2(new_n719), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n903), .A2(new_n916), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n845), .B1(new_n917), .B2(new_n918), .ZN(G367));
  INV_X1    g0719(.A(new_n778), .ZN(new_n920));
  INV_X1    g0720(.A(new_n385), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n675), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n239), .A2(new_n783), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n725), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n522), .A2(new_n668), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n539), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n639), .B2(new_n925), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n750), .A2(G283), .B1(G317), .B2(new_n758), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n729), .A2(new_n207), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n266), .B(new_n929), .C1(G303), .C2(new_n823), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n736), .A2(G294), .B1(new_n740), .B2(G311), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n731), .A2(KEYINPUT46), .A3(new_n560), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT46), .B1(new_n731), .B2(new_n560), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n756), .A2(G107), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n928), .A2(new_n930), .A3(new_n931), .A4(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT109), .ZN(new_n936));
  XOR2_X1   g0736(.A(KEYINPUT111), .B(G137), .Z(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n750), .A2(G50), .B1(new_n758), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(G143), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n741), .A2(new_n940), .B1(new_n313), .B2(new_n739), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n737), .A2(new_n407), .B1(new_n731), .B2(new_n404), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n266), .B1(new_n221), .B2(new_n729), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT110), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n755), .A2(new_n357), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n945), .B2(new_n944), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n939), .A2(new_n943), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n936), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT113), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n950), .B(new_n952), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n924), .B1(new_n927), .B2(new_n788), .C1(new_n953), .C2(new_n727), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n513), .B(new_n543), .C1(new_n487), .C2(new_n668), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n543), .A2(new_n668), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n673), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT42), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n543), .B1(new_n955), .B2(new_n610), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n958), .A2(KEYINPUT42), .B1(new_n668), .B2(new_n960), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n959), .A2(new_n961), .B1(KEYINPUT43), .B2(new_n927), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n670), .A2(new_n957), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n964), .B(new_n965), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n673), .A2(new_n671), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(new_n957), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT45), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n957), .ZN(new_n970));
  XOR2_X1   g0770(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n670), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n969), .A2(new_n670), .A3(new_n972), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n673), .B1(new_n669), .B2(new_n672), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n664), .B2(KEYINPUT108), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n664), .A2(KEYINPUT108), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n979), .B(new_n980), .Z(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n717), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n717), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n676), .B(KEYINPUT41), .Z(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n721), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n954), .B1(new_n966), .B2(new_n986), .ZN(G387));
  OR2_X1    g0787(.A1(new_n669), .A2(new_n788), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n783), .B1(new_n236), .B2(new_n255), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n678), .B2(new_n780), .ZN(new_n990));
  OR3_X1    g0790(.A1(new_n311), .A2(KEYINPUT50), .A3(G50), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT50), .B1(new_n311), .B2(G50), .ZN(new_n992));
  AOI21_X1  g0792(.A(G45), .B1(G68), .B2(G77), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n991), .A2(new_n678), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n990), .A2(new_n994), .B1(new_n208), .B2(new_n675), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n722), .B1(new_n995), .B2(new_n920), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G311), .A2(new_n736), .B1(new_n823), .B2(G317), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n770), .B2(new_n741), .C1(new_n749), .C2(new_n555), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT48), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n999), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n756), .A2(G283), .B1(G294), .B2(new_n732), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT49), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n272), .B1(new_n729), .B2(new_n560), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G326), .B2(new_n758), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n732), .A2(new_n220), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n737), .B2(new_n311), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n929), .B(new_n1011), .C1(G159), .C2(new_n740), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n756), .A2(new_n921), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n266), .B1(new_n202), .B2(new_n739), .C1(new_n746), .C2(new_n357), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G150), .B2(new_n758), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1009), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n996), .B1(new_n1017), .B2(new_n726), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n981), .A2(new_n721), .B1(new_n988), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n982), .A2(new_n676), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n981), .A2(new_n717), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(G393));
  OR2_X1    g0822(.A1(new_n977), .A2(new_n982), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n977), .A2(new_n982), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n676), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n957), .A2(new_n777), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT114), .Z(new_n1027));
  OAI21_X1  g0827(.A(new_n778), .B1(new_n207), .B2(new_n212), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n243), .B2(new_n783), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n737), .A2(new_n202), .B1(new_n731), .B2(new_n357), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n272), .B(new_n1030), .C1(G87), .C2(new_n815), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n940), .B2(new_n759), .C1(new_n311), .C2(new_n749), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n741), .A2(new_n313), .B1(new_n407), .B2(new_n739), .ZN(new_n1033));
  XOR2_X1   g0833(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(new_n205), .C2(new_n755), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G317), .A2(new_n740), .B1(new_n823), .B2(G311), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT52), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n266), .B(new_n730), .C1(G294), .C2(new_n745), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n736), .A2(G303), .B1(new_n732), .B2(G283), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n560), .B2(new_n755), .C1(new_n770), .C2(new_n759), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1032), .A2(new_n1037), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n725), .B(new_n1029), .C1(new_n1044), .C2(new_n726), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1027), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1025), .B(new_n1046), .C1(new_n720), .C2(new_n977), .ZN(G390));
  NAND3_X1  g0847(.A1(new_n696), .A2(G330), .A3(new_n801), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n860), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n850), .B1(new_n891), .B2(new_n892), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n1048), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(KEYINPUT117), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT117), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1051), .A2(new_n1054), .A3(new_n1048), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n802), .A2(new_n797), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n715), .A2(new_n668), .A3(new_n796), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n797), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1050), .A2(new_n1060), .A3(new_n1052), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1057), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n914), .A2(new_n846), .A3(new_n634), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n908), .B1(new_n905), .B2(new_n907), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n904), .B2(new_n910), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1059), .A2(new_n860), .ZN(new_n1068));
  AOI221_X4 g0868(.A(new_n896), .B1(new_n873), .B2(new_n877), .C1(new_n449), .C2(new_n867), .ZN(new_n1069));
  AOI21_X1  g0869(.A(KEYINPUT38), .B1(new_n883), .B2(new_n885), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n909), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(KEYINPUT116), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT116), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1074), .B(new_n1071), .C1(new_n1059), .C2(new_n860), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1067), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1050), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n893), .A2(new_n851), .B1(new_n1058), .B2(new_n797), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1074), .B1(new_n1079), .B2(new_n1071), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1068), .A2(KEYINPUT116), .A3(new_n1072), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1050), .B1(new_n1082), .B2(new_n1067), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1065), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1063), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1082), .A2(new_n1067), .A3(new_n1050), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1084), .A2(new_n676), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n725), .B1(new_n311), .B2(new_n809), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n736), .A2(new_n938), .B1(new_n823), .B2(G132), .ZN(new_n1091));
  INV_X1    g0891(.A(G128), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1091), .B1(new_n1092), .B2(new_n741), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT54), .B(G143), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n749), .A2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(G125), .C2(new_n758), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n266), .B1(new_n729), .B2(new_n202), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT118), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n732), .A2(G150), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT53), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(G159), .C2(new_n756), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n759), .A2(new_n599), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n272), .B1(new_n731), .B2(new_n425), .C1(new_n560), .C2(new_n739), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(new_n750), .C2(G97), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n819), .B1(G107), .B2(new_n736), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n763), .B2(new_n741), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G77), .B2(new_n756), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1096), .A2(new_n1101), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1090), .B1(new_n1108), .B2(new_n727), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n1066), .B2(new_n775), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1078), .A2(new_n1083), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1110), .B1(new_n1111), .B2(new_n721), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1089), .A2(new_n1112), .ZN(G378));
  NAND2_X1  g0913(.A1(new_n1088), .A2(new_n1064), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n913), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n327), .B1(new_n326), .B2(new_n280), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n280), .ZN(new_n1117));
  AOI211_X1 g0917(.A(KEYINPUT10), .B(new_n1117), .C1(new_n325), .C2(new_n320), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n376), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n657), .B1(new_n307), .B2(new_n316), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1120), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n329), .A2(new_n376), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n899), .A2(new_n698), .A3(new_n1129), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1125), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n860), .A2(new_n898), .A3(new_n889), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1051), .A2(new_n1135), .A3(new_n888), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT40), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1133), .B1(new_n1138), .B2(G330), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1115), .B1(new_n1130), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT122), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1129), .B1(new_n899), .B2(new_n698), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1138), .A2(G330), .A3(new_n1133), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n913), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1140), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  OAI211_X1 g0945(.A(KEYINPUT122), .B(new_n1115), .C1(new_n1130), .C2(new_n1139), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1114), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT57), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n677), .B1(new_n1150), .B2(new_n1114), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1145), .A2(new_n721), .A3(new_n1146), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n809), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n722), .B1(G50), .B2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT121), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n745), .A2(G137), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1092), .B2(new_n739), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G132), .B2(new_n736), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1094), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n740), .A2(G125), .B1(new_n732), .B2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1159), .B(new_n1161), .C1(new_n313), .C2(new_n755), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT59), .Z(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(KEYINPUT120), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(KEYINPUT120), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n758), .A2(G124), .ZN(new_n1167));
  AOI211_X1 g0967(.A(G33), .B(G41), .C1(new_n815), .C2(G159), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n266), .B(new_n492), .C1(new_n823), .C2(G107), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n763), .B2(new_n759), .C1(new_n385), .C2(new_n746), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n729), .A2(new_n404), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G116), .B2(new_n740), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1173), .B(new_n1010), .C1(new_n207), .C2(new_n737), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n1171), .A2(new_n947), .A3(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT119), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(KEYINPUT58), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n202), .B1(G33), .B2(G41), .C1(new_n492), .C2(new_n266), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1176), .A2(KEYINPUT58), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1169), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1156), .B1(new_n1180), .B2(new_n726), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1129), .B2(new_n776), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1153), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1152), .A2(new_n1184), .ZN(G375));
  NAND2_X1  g0985(.A1(new_n1051), .A2(new_n775), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT123), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n722), .B1(G68), .B2(new_n1154), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n737), .A2(new_n1094), .B1(new_n731), .B2(new_n407), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1172), .B(new_n1189), .C1(G132), .C2(new_n740), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n756), .A2(G50), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n758), .A2(G128), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n266), .B1(new_n746), .B2(new_n313), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n823), .B2(new_n938), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n272), .B1(new_n739), .B2(new_n763), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n737), .A2(new_n560), .B1(new_n729), .B2(new_n205), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(G294), .C2(new_n740), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1198), .B(new_n1013), .C1(new_n208), .C2(new_n749), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n758), .A2(G303), .B1(new_n732), .B2(G97), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT124), .Z(new_n1201));
  OAI21_X1  g1001(.A(new_n1195), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1188), .B1(new_n1202), .B2(new_n726), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1062), .A2(new_n721), .B1(new_n1187), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1086), .A2(new_n984), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1050), .A2(new_n1060), .A3(new_n1052), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1054), .B1(new_n860), .B2(new_n1049), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1208), .A2(new_n1052), .B1(new_n797), .B2(new_n802), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1207), .B1(new_n1209), .B2(new_n1055), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1063), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1205), .B1(new_n1206), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(G381));
  OR2_X1    g1013(.A1(G393), .A2(G396), .ZN(new_n1214));
  OR3_X1    g1014(.A1(G390), .A2(G384), .A3(new_n1214), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1215), .A2(G387), .A3(G381), .ZN(new_n1216));
  INV_X1    g1016(.A(G378), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1183), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(G407));
  NOR2_X1   g1019(.A1(new_n655), .A2(G343), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1217), .A3(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G407), .A2(G213), .A3(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT125), .ZN(G409));
  NAND2_X1  g1023(.A1(new_n1220), .A2(G2897), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1057), .A2(new_n1063), .A3(KEYINPUT60), .A4(new_n1061), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n676), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT60), .B1(new_n1210), .B2(new_n1063), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1211), .B2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n833), .B(new_n808), .C1(new_n1229), .C2(new_n1205), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1228), .A2(new_n1211), .ZN(new_n1231));
  OAI211_X1 g1031(.A(G384), .B(new_n1204), .C1(new_n1231), .C2(new_n1227), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1225), .B1(new_n1233), .B2(KEYINPUT126), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT126), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1236), .A3(new_n1224), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1234), .A2(new_n1237), .B1(KEYINPUT126), .B2(new_n1233), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1152), .A2(G378), .A3(new_n1184), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1114), .A2(new_n1145), .A3(new_n985), .A4(new_n1146), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1182), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1242), .B2(new_n721), .ZN(new_n1243));
  AOI21_X1  g1043(.A(G378), .B1(new_n1240), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1239), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1220), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT61), .B1(new_n1238), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT63), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1248), .B2(new_n1235), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(G387), .B(G390), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(G393), .B(new_n790), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1252), .B(new_n1253), .Z(new_n1254));
  AOI21_X1  g1054(.A(new_n1220), .B1(new_n1239), .B2(new_n1245), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(KEYINPUT63), .A3(new_n1233), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1249), .A2(new_n1251), .A3(new_n1254), .A4(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1224), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1259));
  AOI211_X1 g1059(.A(KEYINPUT126), .B(new_n1225), .C1(new_n1230), .C2(new_n1232), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n1259), .A2(new_n1260), .B1(new_n1236), .B2(new_n1235), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1258), .B1(new_n1261), .B2(new_n1255), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT127), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(KEYINPUT62), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1255), .B2(new_n1233), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1244), .B1(new_n1218), .B2(G378), .ZN(new_n1266));
  XOR2_X1   g1066(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1267));
  NOR4_X1   g1067(.A1(new_n1266), .A2(new_n1220), .A3(new_n1235), .A4(new_n1267), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1262), .A2(new_n1265), .A3(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1257), .B1(new_n1269), .B2(new_n1254), .ZN(G405));
  INV_X1    g1070(.A(new_n1254), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G375), .A2(new_n1217), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1239), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1233), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1272), .A2(new_n1235), .A3(new_n1239), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1271), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1254), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(G402));
endmodule


