

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747;

  INV_X2 U367 ( .A(G953), .ZN(n733) );
  XNOR2_X1 U368 ( .A(n552), .B(KEYINPUT97), .ZN(n667) );
  XNOR2_X1 U369 ( .A(n399), .B(n398), .ZN(n643) );
  NAND2_X4 U370 ( .A1(n383), .A2(n380), .ZN(n394) );
  AND2_X2 U371 ( .A1(n385), .A2(n384), .ZN(n383) );
  XNOR2_X2 U372 ( .A(n583), .B(KEYINPUT1), .ZN(n688) );
  NOR2_X1 U373 ( .A1(n586), .A2(n351), .ZN(n397) );
  NOR2_X1 U374 ( .A1(n534), .A2(n486), .ZN(n395) );
  NAND2_X1 U375 ( .A1(n382), .A2(n381), .ZN(n380) );
  NOR2_X1 U376 ( .A1(n732), .A2(KEYINPUT2), .ZN(n381) );
  NAND2_X1 U377 ( .A1(n423), .A2(KEYINPUT100), .ZN(n390) );
  XNOR2_X1 U378 ( .A(n397), .B(n396), .ZN(n534) );
  XNOR2_X1 U379 ( .A(n566), .B(KEYINPUT19), .ZN(n586) );
  XNOR2_X1 U380 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U381 ( .A(n373), .B(n498), .ZN(n583) );
  XOR2_X1 U382 ( .A(KEYINPUT59), .B(n630), .Z(n631) );
  XNOR2_X1 U383 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U384 ( .A(G143), .B(G128), .ZN(n455) );
  INV_X1 U385 ( .A(n423), .ZN(n345) );
  XNOR2_X1 U386 ( .A(n395), .B(n363), .ZN(n527) );
  BUF_X1 U387 ( .A(n716), .Z(n346) );
  XNOR2_X1 U388 ( .A(n431), .B(n499), .ZN(n716) );
  XNOR2_X1 U389 ( .A(n427), .B(n426), .ZN(n499) );
  XNOR2_X1 U390 ( .A(n422), .B(G119), .ZN(n427) );
  BUF_X1 U391 ( .A(n695), .Z(n401) );
  INV_X1 U392 ( .A(KEYINPUT82), .ZN(n444) );
  INV_X1 U393 ( .A(KEYINPUT100), .ZN(n425) );
  XNOR2_X1 U394 ( .A(n510), .B(n509), .ZN(n695) );
  XNOR2_X1 U395 ( .A(n489), .B(n488), .ZN(n500) );
  XNOR2_X1 U396 ( .A(G134), .B(G131), .ZN(n488) );
  NOR2_X1 U397 ( .A1(n681), .A2(n484), .ZN(n485) );
  NOR2_X1 U398 ( .A1(G953), .A2(G237), .ZN(n501) );
  NAND2_X1 U399 ( .A1(n732), .A2(KEYINPUT2), .ZN(n384) );
  AND2_X1 U400 ( .A1(n741), .A2(n541), .ZN(n376) );
  INV_X1 U401 ( .A(KEYINPUT0), .ZN(n396) );
  NAND2_X1 U402 ( .A1(n695), .A2(n678), .ZN(n421) );
  INV_X1 U403 ( .A(KEYINPUT30), .ZN(n420) );
  OR2_X1 U404 ( .A1(n625), .A2(G902), .ZN(n373) );
  XOR2_X1 U405 ( .A(G101), .B(G110), .Z(n492) );
  XNOR2_X1 U406 ( .A(n500), .B(n490), .ZN(n730) );
  XNOR2_X1 U407 ( .A(n369), .B(KEYINPUT33), .ZN(n708) );
  NOR2_X1 U408 ( .A1(n372), .A2(n370), .ZN(n369) );
  INV_X1 U409 ( .A(n558), .ZN(n370) );
  NAND2_X1 U410 ( .A1(n443), .A2(G214), .ZN(n678) );
  NOR2_X1 U411 ( .A1(n535), .A2(n708), .ZN(n536) );
  INV_X1 U412 ( .A(n372), .ZN(n545) );
  AND2_X1 U413 ( .A1(n413), .A2(n543), .ZN(n393) );
  AND2_X1 U414 ( .A1(n359), .A2(n414), .ZN(n413) );
  INV_X1 U415 ( .A(KEYINPUT65), .ZN(n414) );
  XNOR2_X1 U416 ( .A(n480), .B(n479), .ZN(n553) );
  XNOR2_X1 U417 ( .A(G137), .B(G116), .ZN(n504) );
  XOR2_X1 U418 ( .A(KEYINPUT85), .B(KEYINPUT23), .Z(n516) );
  XNOR2_X1 U419 ( .A(G128), .B(KEYINPUT24), .ZN(n515) );
  XNOR2_X1 U420 ( .A(G119), .B(G110), .ZN(n514) );
  XOR2_X1 U421 ( .A(G137), .B(G140), .Z(n513) );
  XNOR2_X1 U422 ( .A(n455), .B(n436), .ZN(n489) );
  XNOR2_X1 U423 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n436) );
  NAND2_X1 U424 ( .A1(G234), .A2(G237), .ZN(n445) );
  INV_X1 U425 ( .A(G237), .ZN(n440) );
  OR2_X1 U426 ( .A1(n688), .A2(n689), .ZN(n372) );
  NAND2_X1 U427 ( .A1(n612), .A2(KEYINPUT100), .ZN(n424) );
  XNOR2_X1 U428 ( .A(n402), .B(n503), .ZN(n505) );
  XNOR2_X1 U429 ( .A(n502), .B(n403), .ZN(n402) );
  INV_X1 U430 ( .A(KEYINPUT88), .ZN(n403) );
  XOR2_X1 U431 ( .A(KEYINPUT95), .B(KEYINPUT7), .Z(n452) );
  XNOR2_X1 U432 ( .A(G134), .B(G122), .ZN(n450) );
  XOR2_X1 U433 ( .A(KEYINPUT66), .B(KEYINPUT8), .Z(n459) );
  XNOR2_X1 U434 ( .A(G140), .B(KEYINPUT91), .ZN(n464) );
  XOR2_X1 U435 ( .A(KEYINPUT12), .B(KEYINPUT92), .Z(n465) );
  INV_X1 U436 ( .A(KEYINPUT67), .ZN(n467) );
  XNOR2_X1 U437 ( .A(n417), .B(KEYINPUT48), .ZN(n416) );
  AND2_X1 U438 ( .A1(n609), .A2(n347), .ZN(n417) );
  BUF_X1 U439 ( .A(n573), .Z(n614) );
  AND2_X1 U440 ( .A1(n419), .A2(n418), .ZN(n572) );
  INV_X1 U441 ( .A(n571), .ZN(n418) );
  XNOR2_X1 U442 ( .A(n421), .B(n420), .ZN(n419) );
  XNOR2_X1 U443 ( .A(n695), .B(n371), .ZN(n558) );
  INV_X1 U444 ( .A(KEYINPUT6), .ZN(n371) );
  XNOR2_X1 U445 ( .A(n730), .B(n497), .ZN(n625) );
  NOR2_X1 U446 ( .A1(n688), .A2(n570), .ZN(n674) );
  XNOR2_X1 U447 ( .A(n374), .B(n538), .ZN(n741) );
  NAND2_X1 U448 ( .A1(n537), .A2(n575), .ZN(n374) );
  XNOR2_X1 U449 ( .A(n547), .B(n546), .ZN(n671) );
  INV_X1 U450 ( .A(KEYINPUT101), .ZN(n398) );
  XNOR2_X1 U451 ( .A(n619), .B(n364), .ZN(n620) );
  AND2_X1 U452 ( .A1(n407), .A2(n350), .ZN(n406) );
  NAND2_X1 U453 ( .A1(n646), .A2(n349), .ZN(n405) );
  AND2_X1 U454 ( .A1(n713), .A2(n400), .ZN(n715) );
  AND2_X1 U455 ( .A1(n712), .A2(n733), .ZN(n400) );
  NOR2_X1 U456 ( .A1(n674), .A2(n354), .ZN(n347) );
  AND2_X1 U457 ( .A1(n358), .A2(n376), .ZN(n348) );
  AND2_X1 U458 ( .A1(n647), .A2(G217), .ZN(n349) );
  AND2_X1 U459 ( .A1(n409), .A2(n410), .ZN(n350) );
  NOR2_X1 U460 ( .A1(n449), .A2(n562), .ZN(n351) );
  NOR2_X1 U461 ( .A1(n583), .A2(n689), .ZN(n352) );
  AND2_X1 U462 ( .A1(G214), .A2(n501), .ZN(n353) );
  OR2_X1 U463 ( .A1(n742), .A2(n592), .ZN(n354) );
  AND2_X1 U464 ( .A1(n688), .A2(n425), .ZN(n355) );
  XNOR2_X1 U465 ( .A(KEYINPUT77), .B(n558), .ZN(n356) );
  OR2_X1 U466 ( .A1(n719), .A2(n732), .ZN(n357) );
  AND2_X1 U467 ( .A1(n652), .A2(n557), .ZN(n358) );
  AND2_X1 U468 ( .A1(n424), .A2(n548), .ZN(n359) );
  AND2_X1 U469 ( .A1(n543), .A2(KEYINPUT65), .ZN(n360) );
  AND2_X1 U470 ( .A1(n622), .A2(n745), .ZN(n361) );
  AND2_X1 U471 ( .A1(n358), .A2(n540), .ZN(n362) );
  XOR2_X1 U472 ( .A(n487), .B(KEYINPUT22), .Z(n363) );
  XNOR2_X1 U473 ( .A(KEYINPUT15), .B(G902), .ZN(n623) );
  XNOR2_X1 U474 ( .A(KEYINPUT62), .B(n618), .ZN(n364) );
  AND2_X1 U475 ( .A1(n439), .A2(G472), .ZN(n365) );
  AND2_X1 U476 ( .A1(n439), .A2(G469), .ZN(n366) );
  AND2_X1 U477 ( .A1(n439), .A2(G210), .ZN(n367) );
  AND2_X1 U478 ( .A1(n439), .A2(G475), .ZN(n368) );
  NOR2_X1 U479 ( .A1(n733), .A2(G952), .ZN(n650) );
  INV_X1 U480 ( .A(n650), .ZN(n410) );
  NAND2_X1 U481 ( .A1(n377), .A2(n375), .ZN(n404) );
  NAND2_X1 U482 ( .A1(n379), .A2(n348), .ZN(n375) );
  NAND2_X1 U483 ( .A1(n378), .A2(n362), .ZN(n377) );
  NAND2_X1 U484 ( .A1(n379), .A2(n741), .ZN(n378) );
  XNOR2_X2 U485 ( .A(n533), .B(KEYINPUT80), .ZN(n379) );
  INV_X1 U486 ( .A(n719), .ZN(n382) );
  NAND2_X1 U487 ( .A1(n719), .A2(KEYINPUT2), .ZN(n385) );
  NAND2_X1 U488 ( .A1(n388), .A2(n386), .ZN(n399) );
  NAND2_X1 U489 ( .A1(n387), .A2(n390), .ZN(n386) );
  AND2_X1 U490 ( .A1(n415), .A2(n393), .ZN(n387) );
  NAND2_X1 U491 ( .A1(n389), .A2(n360), .ZN(n388) );
  NAND2_X1 U492 ( .A1(n391), .A2(n390), .ZN(n389) );
  INV_X1 U493 ( .A(n392), .ZN(n391) );
  NAND2_X1 U494 ( .A1(n415), .A2(n359), .ZN(n392) );
  NAND2_X1 U495 ( .A1(n394), .A2(n366), .ZN(n627) );
  NAND2_X1 U496 ( .A1(n394), .A2(n367), .ZN(n640) );
  NAND2_X1 U497 ( .A1(n394), .A2(n368), .ZN(n632) );
  NAND2_X1 U498 ( .A1(n394), .A2(n365), .ZN(n619) );
  NAND2_X1 U499 ( .A1(n394), .A2(n439), .ZN(n412) );
  XNOR2_X2 U500 ( .A(n404), .B(KEYINPUT45), .ZN(n719) );
  AND2_X1 U501 ( .A1(n406), .A2(n405), .ZN(G66) );
  NAND2_X1 U502 ( .A1(n412), .A2(n408), .ZN(n407) );
  INV_X1 U503 ( .A(n647), .ZN(n408) );
  OR2_X1 U504 ( .A1(n647), .A2(G217), .ZN(n409) );
  INV_X1 U505 ( .A(n412), .ZN(n646) );
  XNOR2_X1 U506 ( .A(n716), .B(n438), .ZN(n635) );
  XNOR2_X2 U507 ( .A(n411), .B(n444), .ZN(n566) );
  NAND2_X1 U508 ( .A1(n573), .A2(n678), .ZN(n411) );
  NAND2_X1 U509 ( .A1(n527), .A2(n355), .ZN(n415) );
  NAND2_X1 U510 ( .A1(n416), .A2(n361), .ZN(n732) );
  XNOR2_X2 U511 ( .A(G113), .B(KEYINPUT3), .ZN(n422) );
  AND2_X1 U512 ( .A1(n345), .A2(n688), .ZN(n542) );
  INV_X1 U513 ( .A(n527), .ZN(n423) );
  NOR2_X2 U514 ( .A1(n641), .A2(n650), .ZN(n642) );
  NOR2_X2 U515 ( .A1(n628), .A2(n650), .ZN(n629) );
  NOR2_X2 U516 ( .A1(n633), .A2(n650), .ZN(n634) );
  XNOR2_X1 U517 ( .A(n466), .B(n353), .ZN(n470) );
  XNOR2_X1 U518 ( .A(n478), .B(G475), .ZN(n479) );
  BUF_X1 U519 ( .A(n635), .Z(n638) );
  XNOR2_X1 U520 ( .A(n621), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U521 ( .A(G101), .B(KEYINPUT69), .ZN(n426) );
  XNOR2_X2 U522 ( .A(G116), .B(G107), .ZN(n454) );
  XNOR2_X2 U523 ( .A(G122), .B(G104), .ZN(n471) );
  XNOR2_X1 U524 ( .A(n454), .B(n471), .ZN(n430) );
  XNOR2_X1 U525 ( .A(KEYINPUT73), .B(KEYINPUT16), .ZN(n428) );
  INV_X1 U526 ( .A(G110), .ZN(n644) );
  XNOR2_X1 U527 ( .A(n428), .B(n644), .ZN(n429) );
  XNOR2_X1 U528 ( .A(n430), .B(n429), .ZN(n431) );
  NAND2_X1 U529 ( .A1(n733), .A2(G224), .ZN(n432) );
  XNOR2_X1 U530 ( .A(n432), .B(KEYINPUT83), .ZN(n435) );
  XNOR2_X2 U531 ( .A(G146), .B(G125), .ZN(n469) );
  XNOR2_X1 U532 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n433) );
  XNOR2_X1 U533 ( .A(n469), .B(n433), .ZN(n434) );
  XNOR2_X1 U534 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U535 ( .A(n437), .B(n489), .ZN(n438) );
  INV_X1 U536 ( .A(n623), .ZN(n439) );
  OR2_X2 U537 ( .A1(n635), .A2(n439), .ZN(n442) );
  INV_X1 U538 ( .A(G902), .ZN(n521) );
  NAND2_X1 U539 ( .A1(n521), .A2(n440), .ZN(n443) );
  AND2_X1 U540 ( .A1(n443), .A2(G210), .ZN(n441) );
  XNOR2_X2 U541 ( .A(n442), .B(n441), .ZN(n573) );
  XNOR2_X1 U542 ( .A(n445), .B(KEYINPUT14), .ZN(n446) );
  XNOR2_X1 U543 ( .A(KEYINPUT74), .B(n446), .ZN(n448) );
  NAND2_X1 U544 ( .A1(n448), .A2(G902), .ZN(n447) );
  XOR2_X1 U545 ( .A(KEYINPUT84), .B(n447), .Z(n559) );
  NOR2_X1 U546 ( .A1(G898), .A2(n733), .ZN(n717) );
  AND2_X1 U547 ( .A1(n559), .A2(n717), .ZN(n449) );
  NAND2_X1 U548 ( .A1(G952), .A2(n448), .ZN(n706) );
  NOR2_X1 U549 ( .A1(n706), .A2(G953), .ZN(n562) );
  XOR2_X1 U550 ( .A(KEYINPUT94), .B(KEYINPUT9), .Z(n451) );
  XNOR2_X1 U551 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U552 ( .A(n453), .B(n452), .ZN(n457) );
  XNOR2_X1 U553 ( .A(n454), .B(n455), .ZN(n456) );
  XNOR2_X1 U554 ( .A(n457), .B(n456), .ZN(n461) );
  NAND2_X1 U555 ( .A1(G234), .A2(n733), .ZN(n458) );
  XNOR2_X1 U556 ( .A(n459), .B(n458), .ZN(n511) );
  AND2_X1 U557 ( .A1(n511), .A2(G217), .ZN(n460) );
  XNOR2_X1 U558 ( .A(n461), .B(n460), .ZN(n648) );
  NOR2_X1 U559 ( .A1(G902), .A2(n648), .ZN(n462) );
  XNOR2_X1 U560 ( .A(n462), .B(KEYINPUT96), .ZN(n463) );
  XNOR2_X1 U561 ( .A(n463), .B(G478), .ZN(n551) );
  XNOR2_X1 U562 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U563 ( .A(n467), .B(KEYINPUT10), .ZN(n468) );
  XNOR2_X1 U564 ( .A(n469), .B(n468), .ZN(n731) );
  XNOR2_X1 U565 ( .A(n470), .B(n731), .ZN(n477) );
  XNOR2_X1 U566 ( .A(G113), .B(G143), .ZN(n472) );
  XOR2_X1 U567 ( .A(n472), .B(G131), .Z(n473) );
  XNOR2_X1 U568 ( .A(n471), .B(n473), .ZN(n475) );
  XOR2_X1 U569 ( .A(KEYINPUT11), .B(KEYINPUT90), .Z(n474) );
  XNOR2_X1 U570 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U571 ( .A(n477), .B(n476), .ZN(n630) );
  NOR2_X1 U572 ( .A1(G902), .A2(n630), .ZN(n480) );
  XNOR2_X1 U573 ( .A(KEYINPUT93), .B(KEYINPUT13), .ZN(n478) );
  NAND2_X1 U574 ( .A1(n551), .A2(n553), .ZN(n681) );
  NAND2_X1 U575 ( .A1(n623), .A2(G234), .ZN(n482) );
  XNOR2_X1 U576 ( .A(KEYINPUT20), .B(KEYINPUT86), .ZN(n481) );
  XNOR2_X1 U577 ( .A(n482), .B(n481), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n522), .A2(G221), .ZN(n483) );
  XOR2_X1 U579 ( .A(KEYINPUT21), .B(n483), .Z(n692) );
  INV_X1 U580 ( .A(n692), .ZN(n484) );
  XNOR2_X1 U581 ( .A(n485), .B(KEYINPUT99), .ZN(n486) );
  INV_X1 U582 ( .A(KEYINPUT72), .ZN(n487) );
  INV_X1 U583 ( .A(n513), .ZN(n490) );
  NAND2_X1 U584 ( .A1(G227), .A2(n733), .ZN(n491) );
  XNOR2_X1 U585 ( .A(n492), .B(n491), .ZN(n496) );
  XOR2_X1 U586 ( .A(KEYINPUT75), .B(G104), .Z(n494) );
  XNOR2_X1 U587 ( .A(G146), .B(G107), .ZN(n493) );
  XNOR2_X1 U588 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U589 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U590 ( .A(KEYINPUT68), .B(G469), .Z(n498) );
  XNOR2_X1 U591 ( .A(n499), .B(n500), .ZN(n507) );
  XOR2_X1 U592 ( .A(G146), .B(KEYINPUT5), .Z(n503) );
  NAND2_X1 U593 ( .A1(n501), .A2(G210), .ZN(n502) );
  XNOR2_X1 U594 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U595 ( .A(n507), .B(n506), .ZN(n618) );
  NAND2_X1 U596 ( .A1(n618), .A2(n521), .ZN(n510) );
  INV_X1 U597 ( .A(KEYINPUT71), .ZN(n508) );
  XNOR2_X1 U598 ( .A(n508), .B(G472), .ZN(n509) );
  INV_X1 U599 ( .A(n401), .ZN(n548) );
  NAND2_X1 U600 ( .A1(G221), .A2(n511), .ZN(n512) );
  XOR2_X1 U601 ( .A(n512), .B(n731), .Z(n520) );
  XNOR2_X1 U602 ( .A(n514), .B(n513), .ZN(n518) );
  XNOR2_X1 U603 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U604 ( .A(n518), .B(n517), .Z(n519) );
  XNOR2_X1 U605 ( .A(n520), .B(n519), .ZN(n647) );
  NAND2_X1 U606 ( .A1(n647), .A2(n521), .ZN(n526) );
  NAND2_X1 U607 ( .A1(G217), .A2(n522), .ZN(n524) );
  XNOR2_X1 U608 ( .A(KEYINPUT87), .B(KEYINPUT25), .ZN(n523) );
  XNOR2_X1 U609 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U610 ( .A(n526), .B(n525), .ZN(n691) );
  INV_X1 U611 ( .A(n691), .ZN(n543) );
  NAND2_X1 U612 ( .A1(n356), .A2(n543), .ZN(n528) );
  NOR2_X1 U613 ( .A1(n528), .A2(n688), .ZN(n529) );
  NAND2_X1 U614 ( .A1(n345), .A2(n529), .ZN(n532) );
  INV_X1 U615 ( .A(KEYINPUT76), .ZN(n530) );
  XNOR2_X1 U616 ( .A(n530), .B(KEYINPUT32), .ZN(n531) );
  XNOR2_X1 U617 ( .A(n532), .B(n531), .ZN(n743) );
  NOR2_X2 U618 ( .A1(n643), .A2(n743), .ZN(n533) );
  NAND2_X1 U619 ( .A1(n691), .A2(n692), .ZN(n689) );
  BUF_X1 U620 ( .A(n534), .Z(n535) );
  XNOR2_X1 U621 ( .A(n536), .B(KEYINPUT34), .ZN(n537) );
  NOR2_X1 U622 ( .A1(n551), .A2(n553), .ZN(n575) );
  INV_X1 U623 ( .A(KEYINPUT35), .ZN(n538) );
  INV_X1 U624 ( .A(KEYINPUT44), .ZN(n539) );
  AND2_X1 U625 ( .A1(n539), .A2(KEYINPUT70), .ZN(n540) );
  XNOR2_X1 U626 ( .A(KEYINPUT70), .B(KEYINPUT44), .ZN(n541) );
  NOR2_X1 U627 ( .A1(n558), .A2(n543), .ZN(n544) );
  NAND2_X1 U628 ( .A1(n542), .A2(n544), .ZN(n652) );
  NAND2_X1 U629 ( .A1(n401), .A2(n545), .ZN(n698) );
  OR2_X1 U630 ( .A1(n535), .A2(n698), .ZN(n547) );
  XOR2_X1 U631 ( .A(KEYINPUT89), .B(KEYINPUT31), .Z(n546) );
  INV_X1 U632 ( .A(n671), .ZN(n550) );
  NAND2_X1 U633 ( .A1(n352), .A2(n548), .ZN(n549) );
  OR2_X1 U634 ( .A1(n535), .A2(n549), .ZN(n653) );
  NAND2_X1 U635 ( .A1(n550), .A2(n653), .ZN(n556) );
  INV_X1 U636 ( .A(n551), .ZN(n554) );
  OR2_X1 U637 ( .A1(n554), .A2(n553), .ZN(n552) );
  INV_X1 U638 ( .A(n667), .ZN(n604) );
  NAND2_X1 U639 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U640 ( .A(n555), .B(KEYINPUT98), .ZN(n656) );
  NAND2_X1 U641 ( .A1(n604), .A2(n656), .ZN(n593) );
  NAND2_X1 U642 ( .A1(n556), .A2(n593), .ZN(n557) );
  NAND2_X1 U643 ( .A1(n667), .A2(n558), .ZN(n564) );
  NAND2_X1 U644 ( .A1(G953), .A2(n559), .ZN(n560) );
  NOR2_X1 U645 ( .A1(G900), .A2(n560), .ZN(n561) );
  NOR2_X1 U646 ( .A1(n562), .A2(n561), .ZN(n571) );
  NOR2_X1 U647 ( .A1(n571), .A2(n691), .ZN(n563) );
  NAND2_X1 U648 ( .A1(n563), .A2(n692), .ZN(n578) );
  NOR2_X1 U649 ( .A1(n564), .A2(n578), .ZN(n565) );
  XNOR2_X1 U650 ( .A(n565), .B(KEYINPUT102), .ZN(n610) );
  BUF_X1 U651 ( .A(n566), .Z(n567) );
  NAND2_X1 U652 ( .A1(n610), .A2(n567), .ZN(n569) );
  XNOR2_X1 U653 ( .A(KEYINPUT36), .B(KEYINPUT81), .ZN(n568) );
  XOR2_X1 U654 ( .A(n569), .B(n568), .Z(n570) );
  NAND2_X1 U655 ( .A1(n352), .A2(n572), .ZN(n602) );
  INV_X1 U656 ( .A(n614), .ZN(n574) );
  NOR2_X1 U657 ( .A1(n602), .A2(n574), .ZN(n576) );
  NAND2_X1 U658 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U659 ( .A(KEYINPUT103), .B(n577), .ZN(n742) );
  INV_X1 U660 ( .A(n578), .ZN(n579) );
  NAND2_X1 U661 ( .A1(n579), .A2(n695), .ZN(n582) );
  XNOR2_X1 U662 ( .A(KEYINPUT28), .B(KEYINPUT105), .ZN(n580) );
  XNOR2_X1 U663 ( .A(n580), .B(KEYINPUT104), .ZN(n581) );
  XNOR2_X1 U664 ( .A(n582), .B(n581), .ZN(n585) );
  INV_X1 U665 ( .A(n583), .ZN(n584) );
  NAND2_X1 U666 ( .A1(n585), .A2(n584), .ZN(n599) );
  OR2_X1 U667 ( .A1(n599), .A2(n586), .ZN(n594) );
  INV_X1 U668 ( .A(n594), .ZN(n665) );
  NAND2_X1 U669 ( .A1(n665), .A2(KEYINPUT79), .ZN(n591) );
  INV_X1 U670 ( .A(KEYINPUT79), .ZN(n587) );
  NAND2_X1 U671 ( .A1(n594), .A2(n587), .ZN(n588) );
  NAND2_X1 U672 ( .A1(n588), .A2(n593), .ZN(n589) );
  NAND2_X1 U673 ( .A1(n589), .A2(KEYINPUT47), .ZN(n590) );
  NAND2_X1 U674 ( .A1(n591), .A2(n590), .ZN(n592) );
  INV_X1 U675 ( .A(n593), .ZN(n683) );
  NOR2_X1 U676 ( .A1(n683), .A2(n594), .ZN(n595) );
  NOR2_X1 U677 ( .A1(KEYINPUT79), .A2(n595), .ZN(n596) );
  NOR2_X1 U678 ( .A1(KEYINPUT47), .A2(n596), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n614), .B(KEYINPUT38), .ZN(n601) );
  INV_X1 U680 ( .A(n601), .ZN(n679) );
  NAND2_X1 U681 ( .A1(n679), .A2(n678), .ZN(n682) );
  NOR2_X1 U682 ( .A1(n682), .A2(n681), .ZN(n598) );
  XNOR2_X1 U683 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n597) );
  XNOR2_X1 U684 ( .A(n598), .B(n597), .ZN(n707) );
  NOR2_X1 U685 ( .A1(n599), .A2(n707), .ZN(n600) );
  XNOR2_X1 U686 ( .A(n600), .B(KEYINPUT42), .ZN(n747) );
  NOR2_X1 U687 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U688 ( .A(n603), .B(KEYINPUT39), .ZN(n616) );
  NOR2_X1 U689 ( .A1(n604), .A2(n616), .ZN(n605) );
  XNOR2_X1 U690 ( .A(n605), .B(KEYINPUT40), .ZN(n746) );
  NOR2_X1 U691 ( .A1(n747), .A2(n746), .ZN(n606) );
  XOR2_X1 U692 ( .A(KEYINPUT46), .B(n606), .Z(n607) );
  NOR2_X1 U693 ( .A1(n608), .A2(n607), .ZN(n609) );
  INV_X1 U694 ( .A(n688), .ZN(n612) );
  NAND2_X1 U695 ( .A1(n678), .A2(n610), .ZN(n611) );
  NOR2_X1 U696 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U697 ( .A(n613), .B(KEYINPUT43), .ZN(n615) );
  OR2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n622) );
  NOR2_X1 U699 ( .A1(n616), .A2(n656), .ZN(n617) );
  XNOR2_X1 U700 ( .A(n617), .B(KEYINPUT107), .ZN(n745) );
  NAND2_X1 U701 ( .A1(n620), .A2(n410), .ZN(n621) );
  XNOR2_X1 U702 ( .A(n622), .B(G140), .ZN(G42) );
  XOR2_X1 U703 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n624) );
  XNOR2_X1 U704 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U705 ( .A(n629), .B(KEYINPUT120), .ZN(G54) );
  XNOR2_X1 U706 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n634), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U708 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n636), .B(KEYINPUT55), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n642), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U712 ( .A(n644), .B(KEYINPUT110), .ZN(n645) );
  XNOR2_X1 U713 ( .A(n643), .B(n645), .ZN(G12) );
  NAND2_X1 U714 ( .A1(n646), .A2(G478), .ZN(n649) );
  XNOR2_X1 U715 ( .A(n649), .B(n648), .ZN(n651) );
  NOR2_X1 U716 ( .A1(n651), .A2(n650), .ZN(G63) );
  XNOR2_X1 U717 ( .A(G101), .B(n652), .ZN(G3) );
  INV_X1 U718 ( .A(n653), .ZN(n657) );
  NAND2_X1 U719 ( .A1(n657), .A2(n667), .ZN(n654) );
  XNOR2_X1 U720 ( .A(n654), .B(KEYINPUT108), .ZN(n655) );
  XNOR2_X1 U721 ( .A(G104), .B(n655), .ZN(G6) );
  XOR2_X1 U722 ( .A(KEYINPUT26), .B(KEYINPUT109), .Z(n659) );
  INV_X1 U723 ( .A(n656), .ZN(n670) );
  NAND2_X1 U724 ( .A1(n657), .A2(n670), .ZN(n658) );
  XNOR2_X1 U725 ( .A(n659), .B(n658), .ZN(n661) );
  XOR2_X1 U726 ( .A(G107), .B(KEYINPUT27), .Z(n660) );
  XNOR2_X1 U727 ( .A(n661), .B(n660), .ZN(G9) );
  XOR2_X1 U728 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n663) );
  NAND2_X1 U729 ( .A1(n665), .A2(n670), .ZN(n662) );
  XNOR2_X1 U730 ( .A(n663), .B(n662), .ZN(n664) );
  XOR2_X1 U731 ( .A(G128), .B(n664), .Z(G30) );
  NAND2_X1 U732 ( .A1(n667), .A2(n665), .ZN(n666) );
  XNOR2_X1 U733 ( .A(n666), .B(G146), .ZN(G48) );
  NAND2_X1 U734 ( .A1(n671), .A2(n667), .ZN(n668) );
  XNOR2_X1 U735 ( .A(n668), .B(KEYINPUT112), .ZN(n669) );
  XNOR2_X1 U736 ( .A(G113), .B(n669), .ZN(G15) );
  XOR2_X1 U737 ( .A(G116), .B(KEYINPUT113), .Z(n673) );
  NAND2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n673), .B(n672), .ZN(G18) );
  XNOR2_X1 U740 ( .A(n674), .B(KEYINPUT114), .ZN(n675) );
  XNOR2_X1 U741 ( .A(n675), .B(KEYINPUT37), .ZN(n676) );
  XNOR2_X1 U742 ( .A(G125), .B(n676), .ZN(G27) );
  NAND2_X1 U743 ( .A1(n357), .A2(KEYINPUT78), .ZN(n677) );
  XNOR2_X1 U744 ( .A(n677), .B(KEYINPUT2), .ZN(n713) );
  NOR2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n685) );
  NOR2_X1 U747 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U749 ( .A(n686), .B(KEYINPUT116), .ZN(n687) );
  NOR2_X1 U750 ( .A1(n708), .A2(n687), .ZN(n703) );
  NAND2_X1 U751 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U752 ( .A(n690), .B(KEYINPUT50), .ZN(n697) );
  NOR2_X1 U753 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U754 ( .A(KEYINPUT49), .B(n693), .Z(n694) );
  NOR2_X1 U755 ( .A1(n401), .A2(n694), .ZN(n696) );
  NAND2_X1 U756 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U757 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U758 ( .A(KEYINPUT51), .B(n700), .ZN(n701) );
  NOR2_X1 U759 ( .A1(n707), .A2(n701), .ZN(n702) );
  NOR2_X1 U760 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U761 ( .A(n704), .B(KEYINPUT52), .ZN(n705) );
  NOR2_X1 U762 ( .A1(n706), .A2(n705), .ZN(n711) );
  NOR2_X1 U763 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U764 ( .A(KEYINPUT117), .B(n709), .Z(n710) );
  NOR2_X1 U765 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U766 ( .A(KEYINPUT53), .B(KEYINPUT118), .ZN(n714) );
  XNOR2_X1 U767 ( .A(n715), .B(n714), .ZN(G75) );
  XOR2_X1 U768 ( .A(KEYINPUT124), .B(n346), .Z(n718) );
  NOR2_X1 U769 ( .A1(n718), .A2(n717), .ZN(n729) );
  NOR2_X1 U770 ( .A1(n719), .A2(G953), .ZN(n726) );
  XOR2_X1 U771 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n721) );
  NAND2_X1 U772 ( .A1(G224), .A2(G953), .ZN(n720) );
  XNOR2_X1 U773 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U774 ( .A(KEYINPUT121), .B(n722), .ZN(n723) );
  NAND2_X1 U775 ( .A1(n723), .A2(G898), .ZN(n724) );
  XNOR2_X1 U776 ( .A(n724), .B(KEYINPUT123), .ZN(n725) );
  NOR2_X1 U777 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U778 ( .A(n727), .B(KEYINPUT125), .ZN(n728) );
  XNOR2_X1 U779 ( .A(n729), .B(n728), .ZN(G69) );
  XOR2_X1 U780 ( .A(n731), .B(n730), .Z(n735) );
  XNOR2_X1 U781 ( .A(n735), .B(n732), .ZN(n734) );
  NAND2_X1 U782 ( .A1(n734), .A2(n733), .ZN(n740) );
  XNOR2_X1 U783 ( .A(G227), .B(n735), .ZN(n736) );
  NAND2_X1 U784 ( .A1(n736), .A2(G900), .ZN(n737) );
  XNOR2_X1 U785 ( .A(KEYINPUT126), .B(n737), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n738), .A2(G953), .ZN(n739) );
  NAND2_X1 U787 ( .A1(n740), .A2(n739), .ZN(G72) );
  XNOR2_X1 U788 ( .A(G122), .B(n741), .ZN(G24) );
  XOR2_X1 U789 ( .A(G143), .B(n742), .Z(G45) );
  XOR2_X1 U790 ( .A(G119), .B(n743), .Z(G21) );
  XOR2_X1 U791 ( .A(G134), .B(KEYINPUT115), .Z(n744) );
  XNOR2_X1 U792 ( .A(n745), .B(n744), .ZN(G36) );
  XOR2_X1 U793 ( .A(G131), .B(n746), .Z(G33) );
  XOR2_X1 U794 ( .A(G137), .B(n747), .Z(G39) );
endmodule

