//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(KEYINPUT16), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n187), .B(KEYINPUT79), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n193), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT68), .B(G119), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n196), .B1(new_n198), .B2(G128), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G128), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n198), .A2(G128), .B1(new_n200), .B2(G119), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n199), .B1(new_n201), .B2(new_n196), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G110), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT24), .B(G110), .Z(new_n204));
  NOR2_X1   g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n195), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(G110), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n201), .A2(new_n204), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n191), .A2(new_n192), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n193), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT22), .B(G137), .ZN(new_n212));
  INV_X1    g026(.A(G953), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n213), .A2(G221), .A3(G234), .ZN(new_n214));
  XOR2_X1   g028(.A(new_n212), .B(new_n214), .Z(new_n215));
  XNOR2_X1  g029(.A(new_n211), .B(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G902), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G217), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(G234), .B2(new_n217), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(G902), .ZN(new_n224));
  XOR2_X1   g038(.A(new_n224), .B(KEYINPUT80), .Z(new_n225));
  NAND2_X1  g039(.A1(new_n216), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G469), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT3), .B1(new_n229), .B2(G107), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n231));
  INV_X1    g045(.A(G107), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(G104), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n230), .B(new_n233), .C1(G104), .C2(new_n232), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n234), .A2(G101), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n229), .A2(G107), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n232), .A2(G104), .ZN(new_n237));
  OAI21_X1  g051(.A(G101), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT1), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(G143), .B2(new_n192), .ZN(new_n241));
  INV_X1    g055(.A(G128), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G143), .B(G146), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n243), .A2(KEYINPUT83), .A3(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT83), .B1(new_n243), .B2(new_n244), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n240), .A3(G128), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n239), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n192), .A2(G143), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n253), .B1(new_n200), .B2(new_n241), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n247), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n249), .B1(new_n255), .B2(new_n239), .ZN(new_n256));
  INV_X1    g070(.A(G137), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT11), .A3(G134), .ZN(new_n258));
  INV_X1    g072(.A(G134), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G137), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G131), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT64), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n257), .A2(G134), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI211_X1 g080(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n257), .C2(G134), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n261), .B(new_n262), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT65), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n259), .A2(G137), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT64), .B1(new_n270), .B2(KEYINPUT11), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n264), .A2(new_n263), .A3(new_n265), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n262), .B1(new_n273), .B2(new_n261), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n261), .B1(new_n266), .B2(new_n267), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G131), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT65), .A3(new_n268), .ZN(new_n278));
  AND4_X1   g092(.A1(KEYINPUT12), .A2(new_n256), .A3(new_n275), .A4(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n269), .A2(new_n274), .ZN(new_n281));
  AOI211_X1 g095(.A(KEYINPUT65), .B(new_n262), .C1(new_n273), .C2(new_n261), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n275), .A2(new_n278), .A3(KEYINPUT70), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT12), .B1(new_n285), .B2(new_n256), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n284), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n239), .A2(KEYINPUT10), .A3(new_n255), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n234), .A2(G101), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n235), .A2(KEYINPUT4), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n244), .A2(KEYINPUT0), .A3(G128), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT0), .B(G128), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n292), .B1(new_n244), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n290), .A2(KEYINPUT4), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n291), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n289), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT10), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n249), .A2(KEYINPUT84), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT84), .B1(new_n249), .B2(new_n299), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n288), .B(new_n298), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(G110), .B(G140), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n213), .A2(G227), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n303), .B(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n287), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n285), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n308), .B1(new_n312), .B2(new_n302), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n228), .B(new_n217), .C1(new_n310), .C2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n228), .A2(new_n217), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n302), .B1(new_n279), .B2(new_n286), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n307), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n312), .B1(new_n309), .B2(KEYINPUT85), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT85), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n302), .B2(new_n308), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n318), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n314), .B(new_n316), .C1(new_n322), .C2(new_n228), .ZN(new_n323));
  INV_X1    g137(.A(G221), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT9), .B(G234), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n324), .B1(new_n326), .B2(new_n217), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(G214), .B1(G237), .B2(G902), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n294), .A2(G125), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(G125), .B2(new_n255), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n213), .A2(G224), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT7), .ZN(new_n335));
  XOR2_X1   g149(.A(new_n333), .B(new_n335), .Z(new_n336));
  INV_X1    g150(.A(G116), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G119), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT69), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n197), .A2(new_n337), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT2), .B(G113), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n339), .A2(new_n340), .ZN(new_n344));
  INV_X1    g158(.A(new_n342), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n291), .A3(new_n296), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT5), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n340), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(G113), .B(new_n350), .C1(new_n341), .C2(new_n349), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n346), .A3(new_n239), .ZN(new_n352));
  XNOR2_X1  g166(.A(G110), .B(G122), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n336), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n351), .A2(new_n346), .ZN(new_n356));
  INV_X1    g170(.A(new_n239), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n352), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n353), .B(KEYINPUT8), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(G902), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n333), .B(new_n334), .Z(new_n363));
  NAND2_X1  g177(.A1(new_n348), .A2(new_n352), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n353), .A2(KEYINPUT86), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n354), .A2(KEYINPUT6), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n364), .A2(KEYINPUT6), .A3(new_n365), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(G210), .B1(G237), .B2(G902), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n362), .A2(new_n368), .A3(new_n370), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n331), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(G234), .A2(G237), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(G952), .A3(new_n213), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT21), .B(G898), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(G902), .A3(G953), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(KEYINPUT96), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n374), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G478), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(KEYINPUT15), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n200), .A2(G143), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n251), .A2(G128), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT94), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n259), .ZN(new_n391));
  INV_X1    g205(.A(new_n387), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT13), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(KEYINPUT93), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n386), .B1(KEYINPUT13), .B2(new_n392), .ZN(new_n395));
  OAI21_X1  g209(.A(G134), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G122), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G116), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(KEYINPUT91), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n337), .A2(G122), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(KEYINPUT92), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(G107), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n391), .A2(new_n396), .A3(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n388), .B(KEYINPUT94), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G134), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n391), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT95), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n232), .B1(new_n399), .B2(KEYINPUT14), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n409), .B(new_n402), .Z(new_n410));
  AND3_X1   g224(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n408), .B1(new_n407), .B2(new_n410), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n404), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n325), .A2(new_n221), .A3(G953), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n404), .B(new_n414), .C1(new_n411), .C2(new_n412), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n385), .B1(new_n418), .B2(new_n217), .ZN(new_n419));
  AOI211_X1 g233(.A(G902), .B(new_n384), .C1(new_n416), .C2(new_n417), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n422));
  XNOR2_X1  g236(.A(G113), .B(G122), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(new_n229), .ZN(new_n424));
  INV_X1    g238(.A(G237), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n213), .A3(G214), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n251), .A2(KEYINPUT87), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n251), .A2(KEYINPUT87), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n426), .B2(new_n427), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT18), .ZN(new_n431));
  OR3_X1    g245(.A1(new_n430), .A2(new_n431), .A3(new_n262), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n194), .A2(new_n192), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n192), .B2(new_n187), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n430), .B1(new_n431), .B2(new_n262), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n430), .A2(new_n262), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n430), .A2(new_n262), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n209), .A2(new_n193), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n437), .B2(new_n438), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n436), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n193), .B1(new_n437), .B2(new_n439), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT19), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n194), .A2(new_n445), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n446), .A2(KEYINPUT89), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(KEYINPUT89), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n187), .A2(new_n445), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT88), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n444), .B1(new_n451), .B2(G146), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n434), .A2(new_n435), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n424), .B1(new_n453), .B2(new_n432), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n424), .A2(new_n443), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(G475), .A2(G902), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n422), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n422), .A3(new_n456), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n424), .A2(KEYINPUT90), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n443), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n217), .B1(new_n443), .B2(new_n460), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n458), .A2(new_n459), .B1(G475), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n421), .A2(new_n464), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n329), .A2(new_n382), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT76), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n283), .A2(new_n295), .A3(new_n284), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT71), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n283), .A2(KEYINPUT71), .A3(new_n284), .A4(new_n295), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n262), .B1(new_n264), .B2(new_n260), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(new_n254), .B2(new_n247), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n268), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n347), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n470), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n425), .A2(new_n213), .A3(G210), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n478), .B(KEYINPUT27), .Z(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT26), .B(G101), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n479), .B(new_n480), .Z(new_n481));
  NAND2_X1  g295(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT30), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n475), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n470), .A2(new_n471), .A3(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n344), .B(new_n342), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT67), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n473), .A2(new_n488), .A3(new_n268), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n488), .B1(new_n473), .B2(new_n268), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n275), .A2(new_n278), .A3(new_n295), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n487), .B1(new_n493), .B2(new_n484), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n486), .A2(KEYINPUT72), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(KEYINPUT72), .B1(new_n486), .B2(new_n494), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n483), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT73), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g313(.A(KEYINPUT73), .B(new_n483), .C1(new_n495), .C2(new_n496), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(KEYINPUT31), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n486), .A2(new_n494), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT72), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n486), .A2(KEYINPUT72), .A3(new_n494), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n482), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT31), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT28), .B1(new_n468), .B2(new_n476), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT75), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT74), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n493), .B2(new_n347), .ZN(new_n511));
  AOI211_X1 g325(.A(KEYINPUT74), .B(new_n487), .C1(new_n491), .C2(new_n492), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n513), .A2(new_n477), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n481), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n506), .A2(new_n507), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n501), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(G472), .A2(G902), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n467), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n520), .ZN(new_n522));
  AOI211_X1 g336(.A(KEYINPUT76), .B(new_n522), .C1(new_n501), .C2(new_n518), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n521), .A2(new_n523), .A3(KEYINPUT32), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n481), .A2(KEYINPUT29), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n470), .A2(new_n471), .A3(new_n474), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n347), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n477), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT77), .B1(new_n528), .B2(KEYINPUT28), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT77), .ZN(new_n530));
  AOI211_X1 g344(.A(new_n530), .B(new_n515), .C1(new_n527), .C2(new_n477), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n509), .B(new_n525), .C1(new_n529), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT78), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n470), .A2(new_n471), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n534), .A2(new_n476), .B1(new_n526), .B2(new_n347), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n530), .B1(new_n535), .B2(new_n515), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n528), .A2(KEYINPUT77), .A3(KEYINPUT28), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT78), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n538), .A2(new_n539), .A3(new_n509), .A4(new_n525), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT75), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n508), .B(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n515), .B1(new_n513), .B2(new_n477), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT29), .B1(new_n544), .B2(new_n481), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n477), .B1(new_n495), .B2(new_n496), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n517), .ZN(new_n547));
  AOI21_X1  g361(.A(G902), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n533), .A2(new_n540), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G472), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n522), .B1(new_n501), .B2(new_n518), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT32), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n227), .B(new_n466), .C1(new_n524), .C2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT97), .B(G101), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(G3));
  INV_X1    g370(.A(G472), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n519), .B2(new_n217), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n521), .A2(new_n558), .A3(new_n523), .ZN(new_n559));
  INV_X1    g373(.A(new_n227), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(new_n329), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n464), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n217), .A2(G478), .ZN(new_n564));
  NOR2_X1   g378(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n418), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT98), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT33), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n416), .A2(new_n569), .A3(new_n570), .A4(new_n417), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n564), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(G478), .B1(new_n418), .B2(new_n217), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n563), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n562), .A2(new_n381), .A3(new_n374), .A4(new_n575), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT34), .B(G104), .Z(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(G6));
  NOR2_X1   g392(.A1(new_n563), .A2(new_n421), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n381), .B(KEYINPUT99), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n374), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n562), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G107), .Z(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(G9));
  INV_X1    g398(.A(new_n215), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(KEYINPUT36), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n211), .B(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n587), .A2(new_n225), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n220), .B2(new_n222), .ZN(new_n589));
  NOR4_X1   g403(.A1(new_n329), .A2(new_n465), .A3(new_n382), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n519), .A2(new_n520), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT76), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n519), .A2(new_n217), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G472), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n551), .A2(new_n467), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n590), .A2(new_n592), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT37), .B(G110), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G12));
  INV_X1    g412(.A(new_n329), .ZN(new_n599));
  INV_X1    g413(.A(new_n589), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n374), .A3(new_n600), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n379), .A2(G900), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n376), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n464), .B(new_n603), .C1(new_n419), .C2(new_n420), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT100), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n524), .B2(new_n553), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G128), .ZN(G30));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n499), .A2(new_n500), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n535), .A2(new_n481), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n217), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(G472), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n552), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n609), .B1(new_n524), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT32), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n592), .A2(new_n616), .A3(new_n595), .ZN(new_n617));
  INV_X1    g431(.A(new_n614), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n618), .A3(KEYINPUT101), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n603), .B(KEYINPUT39), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT40), .B1(new_n329), .B2(new_n622), .ZN(new_n623));
  OR3_X1    g437(.A1(new_n329), .A2(KEYINPUT40), .A3(new_n622), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n563), .B1(new_n419), .B2(new_n420), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n625), .A2(new_n331), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n372), .A2(new_n373), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT38), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n626), .A2(new_n629), .A3(new_n600), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n620), .A2(new_n623), .A3(new_n624), .A4(new_n630), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n631), .A2(KEYINPUT102), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(KEYINPUT102), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT103), .B(G143), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G45));
  NAND2_X1  g450(.A1(new_n575), .A2(new_n603), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n601), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n638), .B1(new_n524), .B2(new_n553), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G146), .ZN(G48));
  NOR2_X1   g454(.A1(new_n310), .A2(new_n313), .ZN(new_n641));
  OAI21_X1  g455(.A(G469), .B1(new_n641), .B2(G902), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n328), .A3(new_n314), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n574), .A2(new_n643), .A3(new_n382), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n227), .B(new_n644), .C1(new_n524), .C2(new_n553), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT41), .B(G113), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G15));
  NAND4_X1  g461(.A1(new_n374), .A2(new_n642), .A3(new_n328), .A4(new_n314), .ZN(new_n648));
  INV_X1    g462(.A(new_n580), .ZN(new_n649));
  NOR4_X1   g463(.A1(new_n648), .A2(new_n421), .A3(new_n563), .A4(new_n649), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n227), .B(new_n650), .C1(new_n524), .C2(new_n553), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G116), .ZN(G18));
  AOI22_X1  g466(.A1(new_n549), .A2(G472), .B1(new_n551), .B2(KEYINPUT32), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n617), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n381), .ZN(new_n655));
  NOR4_X1   g469(.A1(new_n648), .A2(new_n465), .A3(new_n655), .A4(new_n589), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G119), .ZN(G21));
  NOR3_X1   g472(.A1(new_n648), .A2(new_n625), .A3(new_n649), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n501), .B1(KEYINPUT31), .B2(new_n497), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n481), .B1(new_n538), .B2(new_n509), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n520), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n594), .A2(new_n659), .A3(new_n662), .A4(new_n227), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G122), .ZN(G24));
  NOR2_X1   g478(.A1(new_n637), .A2(new_n648), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n665), .A2(new_n594), .A3(new_n600), .A4(new_n662), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT104), .B(G125), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G27));
  INV_X1    g482(.A(new_n637), .ZN(new_n669));
  INV_X1    g483(.A(new_n627), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n330), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n329), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n654), .A2(new_n227), .A3(new_n669), .A4(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n591), .A2(new_n616), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n560), .B1(new_n653), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n669), .A2(new_n672), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n674), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n673), .A2(new_n674), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n262), .ZN(G33));
  AOI21_X1  g494(.A(new_n560), .B1(new_n617), .B2(new_n653), .ZN(new_n681));
  INV_X1    g495(.A(new_n605), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n672), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G134), .ZN(G36));
  INV_X1    g498(.A(new_n671), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n464), .B1(new_n572), .B2(new_n573), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT43), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n686), .A2(KEYINPUT107), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT107), .B1(new_n686), .B2(new_n690), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OR3_X1    g508(.A1(new_n694), .A2(new_n559), .A3(new_n589), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n685), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT108), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n699), .B(new_n685), .C1(new_n695), .C2(new_n696), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n695), .A2(new_n696), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n322), .A2(new_n702), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n318), .B(KEYINPUT45), .C1(new_n319), .C2(new_n321), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(G469), .A3(new_n704), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n705), .A2(KEYINPUT105), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(KEYINPUT105), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n315), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n314), .B1(new_n708), .B2(KEYINPUT46), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n710));
  AOI211_X1 g524(.A(new_n710), .B(new_n315), .C1(new_n706), .C2(new_n707), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n328), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n622), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n698), .A2(new_n700), .A3(new_n701), .A4(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT109), .B(G137), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G39));
  NOR4_X1   g530(.A1(new_n654), .A2(new_n227), .A3(new_n637), .A4(new_n671), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT47), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n712), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g535(.A(KEYINPUT47), .B(new_n328), .C1(new_n709), .C2(new_n711), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n717), .A2(new_n718), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n719), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G140), .ZN(G42));
  INV_X1    g540(.A(new_n620), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n671), .A2(new_n643), .ZN(new_n728));
  INV_X1    g542(.A(new_n376), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n728), .A2(new_n227), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n727), .A2(new_n575), .A3(new_n730), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n594), .A2(new_n662), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n227), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n729), .B1(new_n692), .B2(new_n693), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n733), .A2(new_n734), .A3(new_n648), .ZN(new_n735));
  INV_X1    g549(.A(G952), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n735), .A2(new_n736), .A3(G953), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n729), .B(new_n728), .C1(new_n692), .C2(new_n693), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AND2_X1   g553(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n676), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n676), .ZN(new_n742));
  NOR2_X1   g556(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n731), .A2(new_n737), .A3(new_n741), .A4(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT118), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n748));
  INV_X1    g562(.A(new_n734), .ZN(new_n749));
  INV_X1    g563(.A(new_n629), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n750), .A2(new_n330), .A3(new_n643), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n749), .A2(new_n227), .A3(new_n732), .A4(new_n751), .ZN(new_n752));
  AOI211_X1 g566(.A(new_n747), .B(new_n748), .C1(new_n752), .C2(KEYINPUT117), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n747), .B1(new_n752), .B2(KEYINPUT117), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n747), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT50), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n753), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n733), .A2(new_n734), .A3(new_n671), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n642), .A2(new_n314), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n328), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n759), .B1(new_n723), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n732), .A2(new_n600), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(new_n738), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n563), .A2(new_n572), .A3(new_n573), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n615), .A2(new_n619), .A3(new_n730), .A4(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n762), .A2(KEYINPUT51), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n746), .B1(new_n758), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n755), .A2(new_n757), .ZN(new_n770));
  INV_X1    g584(.A(new_n753), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n762), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n762), .A2(new_n773), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n772), .B(new_n767), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n769), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n779));
  INV_X1    g593(.A(new_n419), .ZN(new_n780));
  INV_X1    g594(.A(new_n420), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n781), .A3(new_n464), .A4(new_n603), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT113), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n783), .A2(new_n600), .A3(new_n672), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n654), .A2(new_n779), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n779), .B1(new_n654), .B2(new_n784), .ZN(new_n786));
  OAI221_X1 g600(.A(new_n683), .B1(new_n763), .B2(new_n677), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n596), .A2(new_n663), .ZN(new_n788));
  INV_X1    g602(.A(new_n656), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n617), .B2(new_n653), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n681), .B1(new_n644), .B2(new_n650), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n579), .B1(new_n574), .B2(KEYINPUT112), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(KEYINPUT112), .B2(new_n574), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n559), .A2(new_n561), .A3(new_n581), .A4(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n791), .A2(new_n792), .A3(new_n554), .A4(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n787), .A2(new_n679), .A3(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n607), .A2(new_n639), .A3(new_n666), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n626), .A2(new_n670), .ZN(new_n799));
  INV_X1    g613(.A(new_n603), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n600), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n599), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n524), .A2(new_n609), .A3(new_n614), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT101), .B1(new_n617), .B2(new_n618), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n798), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n802), .B1(new_n615), .B2(new_n619), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n607), .A2(new_n639), .A3(new_n666), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT52), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n808), .A2(new_n811), .A3(KEYINPUT115), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT115), .B1(new_n808), .B2(new_n811), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n797), .B(KEYINPUT53), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n657), .A2(new_n554), .A3(new_n596), .A4(new_n663), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n645), .A2(new_n651), .A3(new_n795), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n673), .A2(new_n674), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n678), .A2(new_n676), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n786), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n654), .A2(new_n779), .A3(new_n784), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n763), .A2(new_n677), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n654), .A2(new_n227), .A3(new_n672), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n826), .B1(new_n827), .B2(new_n682), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n819), .A2(new_n822), .A3(new_n825), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n808), .A2(new_n811), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n816), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n814), .A2(new_n815), .A3(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n829), .A2(new_n830), .A3(new_n816), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n797), .B1(new_n812), .B2(new_n813), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n833), .B1(new_n834), .B2(new_n816), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n778), .B(new_n832), .C1(new_n815), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT120), .ZN(new_n837));
  INV_X1    g651(.A(new_n835), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT54), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n840), .A3(new_n832), .A4(new_n778), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n736), .A2(new_n213), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n837), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n760), .A2(KEYINPUT49), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n760), .A2(KEYINPUT49), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n629), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n687), .A2(new_n227), .A3(new_n328), .A4(new_n330), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT111), .ZN(new_n848));
  AOI211_X1 g662(.A(new_n844), .B(new_n846), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n727), .B(new_n849), .C1(new_n848), .C2(new_n847), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n843), .A2(new_n850), .ZN(G75));
  AOI21_X1  g665(.A(new_n217), .B1(new_n814), .B2(new_n831), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(G210), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT56), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n366), .ZN(new_n856));
  INV_X1    g670(.A(new_n367), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(new_n363), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT55), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n855), .A2(new_n860), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n213), .A2(G952), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(G51));
  XOR2_X1   g678(.A(new_n641), .B(KEYINPUT121), .Z(new_n865));
  NAND2_X1  g679(.A1(new_n814), .A2(new_n831), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT54), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n832), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n315), .B(KEYINPUT57), .Z(new_n870));
  OAI21_X1  g684(.A(new_n865), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n852), .A2(new_n706), .A3(new_n707), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n863), .B1(new_n871), .B2(new_n872), .ZN(G54));
  AND2_X1   g687(.A1(KEYINPUT58), .A2(G475), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n852), .A2(new_n455), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n455), .B1(new_n852), .B2(new_n874), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n875), .A2(new_n876), .A3(new_n863), .ZN(G60));
  OAI21_X1  g691(.A(new_n832), .B1(new_n835), .B2(new_n815), .ZN(new_n878));
  NAND2_X1  g692(.A1(G478), .A2(G902), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT59), .Z(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n568), .A2(new_n571), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n884), .A2(new_n880), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n863), .B1(new_n868), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n814), .A2(new_n815), .A3(new_n831), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n815), .B1(new_n814), .B2(new_n831), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n863), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n883), .B1(new_n878), .B2(new_n881), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT122), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n889), .A2(new_n896), .ZN(G63));
  NAND2_X1  g711(.A1(G217), .A2(G902), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT60), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n814), .B2(new_n831), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n587), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n901), .B(new_n893), .C1(new_n216), .C2(new_n900), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n902), .B(new_n903), .ZN(G66));
  INV_X1    g718(.A(G224), .ZN(new_n905));
  OAI21_X1  g719(.A(G953), .B1(new_n377), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n819), .B2(G953), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n856), .B(new_n857), .C1(G898), .C2(new_n213), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(G69));
  NAND2_X1  g723(.A1(new_n493), .A2(new_n484), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n486), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT123), .Z(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(new_n451), .Z(new_n913));
  NAND3_X1  g727(.A1(new_n713), .A2(new_n676), .A3(new_n799), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n914), .A2(new_n683), .A3(new_n798), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n714), .A2(new_n915), .A3(new_n822), .A4(new_n725), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n213), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n213), .A2(G900), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n913), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n632), .A2(new_n633), .A3(new_n798), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(KEYINPUT62), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n794), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n794), .A2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n329), .A2(new_n671), .A3(new_n622), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n924), .A2(new_n681), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT125), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n714), .A2(new_n725), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n921), .A2(KEYINPUT62), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n922), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n213), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n920), .B1(new_n932), .B2(new_n913), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n213), .B1(G227), .B2(G900), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT126), .Z(new_n935));
  XNOR2_X1  g749(.A(new_n933), .B(new_n935), .ZN(G72));
  XNOR2_X1  g750(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n937));
  NAND2_X1  g751(.A1(G472), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n931), .B2(new_n796), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n481), .A3(new_n546), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n499), .A2(new_n547), .A3(new_n500), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n838), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n939), .B1(new_n916), .B2(new_n796), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n546), .A2(new_n481), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n863), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n941), .A2(new_n943), .A3(new_n947), .ZN(G57));
endmodule


