//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT0), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n215), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n211), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n212), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n219), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G226), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT66), .B(G232), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G58), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(G1), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G13), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(new_n209), .ZN(new_n248));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n208), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT67), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n246), .A2(G20), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(G50), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n248), .A2(new_n202), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n209), .A2(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n250), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n254), .A2(KEYINPUT9), .A3(new_n255), .A4(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT9), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT67), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n251), .B(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n253), .A2(G50), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n261), .A2(new_n255), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n263), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G223), .A3(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G77), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G222), .ZN(new_n275));
  OAI221_X1 g0075(.A(new_n271), .B1(new_n272), .B2(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n208), .B1(G33), .B2(G41), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  INV_X1    g0079(.A(G45), .ZN(new_n280));
  AOI21_X1  g0080(.A(G1), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G274), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n277), .A2(new_n281), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(G226), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n278), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G200), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n278), .A2(G190), .A3(new_n285), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n262), .A2(new_n269), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT68), .B1(new_n289), .B2(KEYINPUT10), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n262), .A2(new_n269), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n287), .A2(new_n288), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT68), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT10), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n291), .A2(new_n292), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n289), .A2(KEYINPUT10), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n286), .A2(G169), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n286), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(new_n267), .B2(new_n268), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT18), .ZN(new_n304));
  INV_X1    g0104(.A(new_n258), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n253), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT75), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n307), .A2(new_n252), .B1(new_n248), .B2(new_n258), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G58), .ZN(new_n310));
  INV_X1    g0110(.A(G68), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(G20), .B1(new_n312), .B2(new_n201), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n256), .A2(G159), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT3), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G33), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n321), .A2(new_n322), .A3(new_n209), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT71), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n319), .A2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT71), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n209), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT7), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n323), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(KEYINPUT16), .B(new_n316), .C1(new_n331), .C2(new_n311), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n332), .A2(new_n250), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT16), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT73), .B1(new_n319), .B2(G33), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT73), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(new_n317), .A3(KEYINPUT3), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n337), .A3(new_n320), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n330), .A2(G20), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n341));
  NOR2_X1   g0141(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n270), .B2(G20), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT74), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n346), .A3(G68), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n316), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n311), .B1(new_n340), .B2(new_n344), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(new_n346), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n334), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n309), .B1(new_n333), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n283), .B1(new_n284), .B2(G232), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n318), .A2(new_n320), .A3(G226), .A4(G1698), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT76), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT76), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n270), .A2(new_n356), .A3(G226), .A4(G1698), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT77), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n318), .A2(new_n320), .A3(G223), .A4(new_n273), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G87), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n358), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n277), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n362), .B1(new_n357), .B2(new_n355), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(new_n359), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n300), .B(new_n353), .C1(new_n365), .C2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n353), .ZN(new_n369));
  INV_X1    g0169(.A(new_n277), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n366), .B2(new_n359), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n358), .A2(new_n363), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT77), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n368), .B1(new_n374), .B2(G169), .ZN(new_n375));
  OAI211_X1 g0175(.A(KEYINPUT78), .B(new_n304), .C1(new_n352), .C2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n304), .B1(new_n352), .B2(new_n375), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n332), .A2(new_n250), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n315), .B1(new_n349), .B2(new_n346), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n321), .A2(new_n209), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(new_n343), .B1(new_n338), .B2(new_n339), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT74), .B1(new_n382), .B2(new_n311), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT16), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n308), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n353), .B1(new_n365), .B2(new_n367), .ZN(new_n386));
  INV_X1    g0186(.A(G169), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n385), .A2(KEYINPUT18), .A3(new_n368), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT78), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n377), .B1(new_n378), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT17), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n371), .A2(new_n373), .ZN(new_n393));
  AOI21_X1  g0193(.A(G200), .B1(new_n393), .B2(new_n353), .ZN(new_n394));
  AOI211_X1 g0194(.A(G190), .B(new_n369), .C1(new_n371), .C2(new_n373), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n392), .B1(new_n396), .B2(new_n385), .ZN(new_n397));
  INV_X1    g0197(.A(G190), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n398), .B(new_n353), .C1(new_n365), .C2(new_n367), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n374), .B2(G200), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n352), .A2(KEYINPUT17), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT14), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(KEYINPUT70), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n270), .A2(G232), .A3(G1698), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  INV_X1    g0206(.A(G226), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n405), .B(new_n406), .C1(new_n274), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n277), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT13), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n283), .B1(new_n284), .B2(G238), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n410), .B1(new_n409), .B2(new_n411), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n404), .B1(new_n415), .B2(new_n387), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n409), .A2(new_n411), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT13), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n412), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(G169), .C1(KEYINPUT70), .C2(new_n403), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n415), .A2(G179), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n416), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n247), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(G20), .A3(new_n311), .ZN(new_n424));
  XOR2_X1   g0224(.A(new_n424), .B(KEYINPUT12), .Z(new_n425));
  AOI22_X1  g0225(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n311), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n272), .B2(new_n259), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n427), .A2(new_n250), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n425), .B1(KEYINPUT11), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n251), .A2(G68), .A3(new_n253), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT69), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n428), .A2(KEYINPUT11), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n422), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n270), .A2(G238), .A3(G1698), .ZN(new_n435));
  INV_X1    g0235(.A(G107), .ZN(new_n436));
  INV_X1    g0236(.A(G232), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n435), .B1(new_n436), .B2(new_n270), .C1(new_n274), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n277), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n283), .B1(new_n284), .B2(G244), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G179), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(G169), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n305), .A2(new_n256), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT15), .B(G87), .ZN(new_n447));
  OAI221_X1 g0247(.A(new_n446), .B1(new_n209), .B2(new_n272), .C1(new_n259), .C2(new_n447), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n448), .A2(new_n250), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n251), .A2(G77), .A3(new_n253), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n423), .A2(G20), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(G77), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n445), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n442), .A2(G200), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n441), .A2(G190), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G200), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n419), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n418), .A2(new_n398), .A3(new_n412), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n433), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n434), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  NOR4_X1   g0265(.A1(new_n303), .A2(new_n391), .A3(new_n402), .A4(new_n465), .ZN(new_n466));
  XOR2_X1   g0266(.A(KEYINPUT88), .B(KEYINPUT21), .Z(new_n467));
  NAND2_X1  g0267(.A1(new_n246), .A2(G45), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT5), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n279), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(new_n277), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G270), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(G274), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT83), .ZN(new_n477));
  OAI21_X1  g0277(.A(G303), .B1(new_n325), .B2(new_n326), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n318), .A2(new_n320), .A3(G264), .A4(G1698), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n318), .A2(new_n320), .A3(G257), .A4(new_n273), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n481), .A2(KEYINPUT82), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT82), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n478), .A2(new_n479), .A3(new_n480), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n277), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n477), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n481), .A2(KEYINPUT82), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n487), .A2(KEYINPUT83), .A3(new_n277), .A4(new_n484), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n476), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n250), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n246), .A2(G33), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n451), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT84), .ZN(new_n493));
  INV_X1    g0293(.A(G116), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G20), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n247), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n423), .A2(KEYINPUT84), .A3(G20), .A4(new_n494), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n492), .A2(G116), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G283), .ZN(new_n499));
  INV_X1    g0299(.A(G97), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n499), .B(new_n209), .C1(G33), .C2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(new_n250), .A3(new_n495), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT20), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT85), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n502), .A2(new_n503), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n504), .A2(KEYINPUT85), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n498), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G169), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n467), .B1(new_n489), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n486), .A2(new_n488), .ZN(new_n513));
  INV_X1    g0313(.A(new_n476), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n508), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n505), .A3(new_n506), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n387), .B1(new_n517), .B2(new_n498), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n515), .A2(KEYINPUT21), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n474), .A2(G179), .A3(new_n475), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(new_n486), .B2(new_n488), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n521), .A2(KEYINPUT86), .A3(new_n509), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT86), .B1(new_n521), .B2(new_n509), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT87), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT87), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n526), .B(new_n519), .C1(new_n522), .C2(new_n523), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n512), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n489), .A2(new_n398), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(G200), .B2(new_n489), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(new_n517), .A3(new_n498), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n492), .A2(G97), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n248), .A2(new_n500), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(KEYINPUT6), .A2(G97), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT79), .B1(new_n535), .B2(G107), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT79), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n537), .A2(new_n436), .A3(KEYINPUT6), .A4(G97), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g0339(.A(G97), .B(G107), .Z(new_n540));
  OAI21_X1  g0340(.A(new_n539), .B1(new_n540), .B2(KEYINPUT6), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G20), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n256), .A2(G77), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n543), .C1(new_n436), .C2(new_n382), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n534), .B1(new_n544), .B2(new_n250), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n270), .A2(G244), .A3(new_n273), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT80), .ZN(new_n547));
  OR2_X1    g0347(.A1(new_n547), .A2(KEYINPUT4), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n270), .A2(G244), .A3(new_n548), .A4(new_n273), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n270), .A2(G250), .A3(G1698), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n499), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n277), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n473), .A2(G257), .B1(G274), .B2(new_n472), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G169), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n554), .A2(G179), .A3(new_n555), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n545), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT19), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n209), .B1(new_n406), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(G87), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(new_n500), .A3(new_n436), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n209), .A2(G33), .A3(G97), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n562), .A2(new_n564), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n270), .A2(new_n209), .A3(G68), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n490), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n447), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n569), .A2(new_n451), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n251), .A2(new_n491), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n571), .B1(new_n447), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n468), .A2(G250), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n246), .A2(G45), .A3(G274), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n277), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n270), .A2(G244), .A3(G1698), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G116), .ZN(new_n578));
  INV_X1    g0378(.A(G238), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n577), .B(new_n578), .C1(new_n274), .C2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n576), .B1(new_n580), .B2(new_n277), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n581), .A2(new_n387), .ZN(new_n582));
  AOI211_X1 g0382(.A(new_n300), .B(new_n576), .C1(new_n580), .C2(new_n277), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n573), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(G190), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n572), .A2(new_n563), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n586), .A2(new_n568), .A3(new_n570), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n585), .B(new_n587), .C1(new_n460), .C2(new_n581), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n554), .A2(new_n398), .A3(new_n555), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n473), .A2(G257), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n475), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n546), .A2(new_n549), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n593), .A2(new_n499), .A3(new_n551), .A4(new_n552), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n592), .B1(new_n594), .B2(new_n277), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n590), .B1(new_n595), .B2(G200), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(KEYINPUT81), .A3(new_n545), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT81), .B1(new_n596), .B2(new_n545), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n560), .B(new_n589), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n572), .A2(new_n436), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n423), .A2(G20), .A3(new_n436), .ZN(new_n602));
  XNOR2_X1  g0402(.A(new_n602), .B(KEYINPUT25), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n318), .A2(new_n320), .A3(new_n209), .A4(G87), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT22), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT22), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n270), .A2(new_n607), .A3(new_n209), .A4(G87), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n578), .A2(G20), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT23), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n209), .B2(G107), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n436), .A2(KEYINPUT23), .A3(G20), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n609), .A2(KEYINPUT24), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n250), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT24), .B1(new_n609), .B2(new_n614), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n604), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT89), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n270), .A2(G250), .A3(new_n273), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n270), .A2(G257), .A3(G1698), .ZN(new_n622));
  NAND2_X1  g0422(.A1(G33), .A2(G294), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n277), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n473), .A2(G264), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n300), .A2(new_n625), .A3(new_n475), .A4(new_n626), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n624), .A2(new_n277), .B1(G264), .B2(new_n473), .ZN(new_n628));
  AOI21_X1  g0428(.A(G169), .B1(new_n628), .B2(new_n475), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n604), .B(KEYINPUT89), .C1(new_n616), .C2(new_n617), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n620), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT90), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n628), .A2(new_n475), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n460), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(G190), .B2(new_n635), .ZN(new_n637));
  INV_X1    g0437(.A(new_n618), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n620), .A2(new_n630), .A3(KEYINPUT90), .A4(new_n631), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n634), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n600), .A2(new_n641), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n466), .A2(new_n528), .A3(new_n531), .A4(new_n642), .ZN(G372));
  NAND2_X1  g0443(.A1(new_n557), .A2(new_n558), .ZN(new_n644));
  INV_X1    g0444(.A(new_n545), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(new_n584), .A4(new_n588), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n584), .B1(new_n646), .B2(KEYINPUT26), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n589), .B2(new_n559), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n511), .B(new_n519), .C1(new_n522), .C2(new_n523), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n630), .A2(new_n618), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n554), .A2(new_n398), .A3(new_n555), .ZN(new_n655));
  AOI21_X1  g0455(.A(G200), .B1(new_n554), .B2(new_n555), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n545), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT81), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n597), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n660), .A2(new_n560), .A3(new_n589), .A4(new_n639), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n650), .B1(new_n654), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n466), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n302), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n378), .A2(new_n389), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n453), .B1(new_n443), .B2(new_n444), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n464), .A2(new_n667), .B1(new_n422), .B2(new_n433), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n666), .B1(new_n668), .B2(new_n402), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n664), .B1(new_n669), .B2(new_n298), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n663), .A2(new_n670), .ZN(G369));
  OR3_X1    g0471(.A1(new_n247), .A2(KEYINPUT27), .A3(G20), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT27), .B1(new_n247), .B2(G20), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G343), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT91), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n528), .A2(new_n531), .B1(new_n509), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G330), .ZN(new_n678));
  INV_X1    g0478(.A(new_n676), .ZN(new_n679));
  AOI211_X1 g0479(.A(new_n679), .B(new_n651), .C1(new_n517), .C2(new_n498), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n620), .A2(new_n631), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n679), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n641), .A2(new_n683), .B1(new_n632), .B2(new_n679), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n528), .A2(new_n676), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n641), .A2(new_n683), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n686), .A2(new_n687), .B1(new_n653), .B2(new_n679), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n213), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR4_X1   g0492(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G1), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n207), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(new_n692), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT28), .ZN(new_n697));
  INV_X1    g0497(.A(new_n520), .ZN(new_n698));
  INV_X1    g0498(.A(new_n485), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT83), .B1(new_n699), .B2(new_n487), .ZN(new_n700));
  INV_X1    g0500(.A(new_n488), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n509), .B(new_n698), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT86), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n521), .A2(KEYINPUT86), .A3(new_n509), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(new_n511), .A3(new_n519), .A4(new_n652), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n559), .B1(new_n659), .B2(new_n597), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n707), .A2(new_n708), .A3(new_n589), .A4(new_n639), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n676), .B1(new_n709), .B2(new_n650), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n634), .A2(new_n640), .ZN(new_n714));
  INV_X1    g0514(.A(new_n527), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n526), .B1(new_n706), .B2(new_n519), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n714), .B(new_n511), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n708), .A2(new_n588), .A3(new_n639), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n676), .B1(new_n720), .B2(new_n650), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n713), .B1(new_n722), .B2(new_n712), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n528), .A2(new_n642), .A3(new_n531), .A4(new_n679), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n581), .A2(new_n628), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT92), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT92), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n581), .A2(new_n628), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT93), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n726), .A2(new_n595), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n521), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n731), .A2(new_n732), .B1(KEYINPUT93), .B2(new_n729), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n728), .A2(new_n595), .A3(new_n730), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n729), .A2(KEYINPUT93), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(new_n521), .A3(new_n726), .A4(new_n735), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n595), .A2(G179), .A3(new_n581), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n515), .A3(new_n635), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n733), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT31), .B1(new_n739), .B2(new_n676), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n678), .B1(new_n724), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n723), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n697), .B1(new_n746), .B2(G1), .ZN(G364));
  INV_X1    g0547(.A(G13), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G45), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n692), .A2(G1), .A3(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n677), .A2(new_n680), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n678), .B1(new_n677), .B2(new_n680), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n208), .B1(G20), .B2(new_n387), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n327), .A2(new_n328), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n690), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n241), .A2(new_n280), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n207), .A2(G45), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n690), .A2(new_n321), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n769), .A2(G355), .B1(new_n494), .B2(new_n690), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n762), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n209), .A2(new_n398), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n460), .A2(G179), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G303), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g0576(.A(KEYINPUT33), .B(G317), .Z(new_n777));
  NOR2_X1   g0577(.A1(new_n300), .A2(new_n460), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n209), .A2(G190), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n300), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n777), .A2(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n772), .A2(new_n778), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n776), .B(new_n784), .C1(G326), .C2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G179), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G190), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G294), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n772), .A2(new_n781), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n270), .B1(new_n793), .B2(G322), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n779), .A2(new_n773), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n779), .A2(new_n788), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G283), .A2(new_n796), .B1(new_n798), .B2(G329), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n787), .A2(new_n791), .A3(new_n794), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT94), .B(G159), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT95), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT32), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n792), .A2(new_n310), .B1(new_n795), .B2(new_n436), .ZN(new_n805));
  INV_X1    g0605(.A(new_n782), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(G77), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n790), .A2(G97), .ZN(new_n808));
  INV_X1    g0608(.A(new_n780), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n321), .B1(new_n809), .B2(G68), .ZN(new_n810));
  INV_X1    g0610(.A(new_n774), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G50), .A2(new_n786), .B1(new_n811), .B2(G87), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n807), .A2(new_n808), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n800), .B1(new_n804), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n771), .B1(new_n814), .B2(new_n760), .ZN(new_n815));
  INV_X1    g0615(.A(new_n759), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n753), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n756), .B1(new_n752), .B2(new_n817), .ZN(G396));
  INV_X1    g0618(.A(KEYINPUT97), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n455), .B2(new_n679), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n667), .A2(KEYINPUT97), .A3(new_n676), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n455), .B(new_n458), .C1(new_n453), .C2(new_n679), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n710), .B(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n751), .B1(new_n825), .B2(new_n744), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n744), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n826), .B1(new_n828), .B2(KEYINPUT98), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(KEYINPUT98), .B2(new_n828), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n774), .A2(new_n436), .B1(new_n797), .B2(new_n783), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n270), .B(new_n831), .C1(G87), .C2(new_n796), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G294), .A2(new_n793), .B1(new_n806), .B2(G116), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n786), .A2(G303), .B1(new_n809), .B2(G283), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n832), .A2(new_n808), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n801), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n786), .A2(G137), .B1(new_n806), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G150), .ZN(new_n838));
  XNOR2_X1  g0638(.A(KEYINPUT96), .B(G143), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(new_n838), .B2(new_n780), .C1(new_n792), .C2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n796), .A2(G68), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G50), .A2(new_n811), .B1(new_n798), .B2(G132), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n763), .B1(G58), .B2(new_n790), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n842), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n840), .A2(new_n841), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n835), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n760), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n760), .A2(new_n757), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n751), .B1(new_n272), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n849), .B(new_n851), .C1(new_n824), .C2(new_n758), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n830), .A2(new_n852), .ZN(G384));
  OAI211_X1 g0653(.A(G116), .B(new_n210), .C1(new_n541), .C2(KEYINPUT35), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT99), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n541), .A2(KEYINPUT35), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT36), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  NOR3_X1   g0662(.A1(new_n695), .A2(new_n272), .A3(new_n312), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n311), .A2(G50), .ZN(new_n864));
  OAI211_X1 g0664(.A(G1), .B(new_n748), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n861), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT100), .Z(new_n867));
  NAND2_X1  g0667(.A1(new_n433), .A2(new_n676), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n434), .B2(new_n464), .ZN(new_n869));
  INV_X1    g0669(.A(new_n868), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n870), .B(new_n463), .C1(new_n422), .C2(new_n433), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n824), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n724), .B2(new_n742), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n385), .A2(new_n368), .A3(new_n388), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n351), .A2(new_n250), .A3(new_n332), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n400), .A2(new_n875), .A3(new_n308), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n385), .A2(new_n674), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n874), .A2(new_n876), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n674), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n375), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n316), .B1(new_n331), .B2(new_n311), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n882), .A2(new_n334), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n308), .B1(new_n883), .B2(new_n379), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n881), .A2(new_n884), .B1(new_n352), .B2(new_n400), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n879), .B1(new_n885), .B2(new_n877), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n390), .A2(new_n378), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n402), .B1(new_n887), .B2(new_n376), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(new_n674), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT102), .ZN(new_n893));
  OAI211_X1 g0693(.A(KEYINPUT38), .B(new_n886), .C1(new_n888), .C2(new_n889), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n893), .B1(new_n892), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n873), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n894), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n874), .A2(new_n876), .A3(new_n878), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT103), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n901), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(new_n879), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n878), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n665), .B2(new_n402), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n873), .B(KEYINPUT40), .C1(new_n900), .C2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n899), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n724), .A2(new_n742), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n466), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n911), .B(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n914), .A2(new_n678), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n667), .A2(new_n679), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT101), .Z(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n710), .B2(new_n824), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n869), .A2(new_n871), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n895), .B2(new_n896), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n434), .A2(new_n676), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n905), .A2(new_n879), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT103), .B1(new_n901), .B2(KEYINPUT37), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n908), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n891), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT39), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n927), .A2(new_n928), .A3(new_n894), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n928), .B1(new_n892), .B2(new_n894), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n923), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n666), .A2(new_n674), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n922), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n466), .B(new_n713), .C1(new_n722), .C2(new_n712), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n670), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n934), .B(new_n936), .Z(new_n937));
  OAI22_X1  g0737(.A1(new_n915), .A2(new_n937), .B1(new_n246), .B2(new_n749), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n915), .A2(new_n937), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n867), .B1(new_n938), .B2(new_n939), .ZN(G367));
  OAI21_X1  g0740(.A(new_n708), .B1(new_n545), .B2(new_n679), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n559), .A2(new_n676), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n686), .A2(new_n684), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n560), .B1(new_n941), .B2(new_n714), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n944), .A2(KEYINPUT42), .B1(new_n679), .B2(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT104), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n944), .A2(KEYINPUT42), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n946), .B2(KEYINPUT104), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n679), .A2(new_n587), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n584), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n589), .B2(new_n951), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT43), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n950), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n947), .A2(new_n949), .A3(new_n954), .A4(new_n953), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n685), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n943), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n959), .B(new_n961), .Z(new_n962));
  XOR2_X1   g0762(.A(new_n691), .B(KEYINPUT41), .Z(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n688), .A2(new_n943), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n964), .B1(new_n688), .B2(new_n943), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n688), .A2(new_n943), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n688), .A2(KEYINPUT45), .A3(new_n943), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n968), .A2(new_n685), .A3(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n971), .A2(new_n972), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n960), .B1(new_n975), .B2(new_n967), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n686), .A2(new_n687), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n684), .B2(new_n686), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT106), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n978), .B1(new_n754), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n681), .A2(KEYINPUT106), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n978), .A2(KEYINPUT106), .A3(new_n681), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n745), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n974), .A2(new_n976), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT107), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n974), .A2(new_n976), .A3(new_n984), .A4(KEYINPUT107), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n963), .B1(new_n989), .B2(new_n746), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n750), .A2(G1), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n962), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n953), .A2(new_n759), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n765), .A2(new_n237), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n762), .B1(new_n690), .B2(new_n569), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n751), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(G317), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n795), .A2(new_n500), .B1(new_n797), .B2(new_n997), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n998), .B(new_n764), .C1(G107), .C2(new_n790), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n811), .A2(G116), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT46), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G294), .A2(new_n809), .B1(new_n806), .B2(G283), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G311), .A2(new_n786), .B1(new_n793), .B2(G303), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(G137), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n795), .A2(new_n272), .B1(new_n797), .B2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n321), .B(new_n1006), .C1(G58), .C2(new_n811), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n809), .A2(new_n836), .B1(new_n806), .B2(G50), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n839), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n786), .A2(new_n1009), .B1(new_n793), .B2(G150), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n790), .A2(G68), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(KEYINPUT47), .B1(new_n1004), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1004), .A2(KEYINPUT47), .A3(new_n1012), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n760), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n993), .B(new_n996), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n992), .A2(new_n1016), .ZN(G387));
  NAND2_X1  g0817(.A1(new_n982), .A2(new_n983), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n991), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT108), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n769), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1021), .A2(new_n693), .B1(G107), .B2(new_n213), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n233), .A2(G45), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n765), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT109), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n280), .B1(new_n311), .B2(new_n272), .C1(new_n693), .C2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n1025), .B2(new_n693), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n258), .A2(G50), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT50), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1024), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1022), .B1(new_n1023), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n752), .B1(new_n1031), .B2(new_n762), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n763), .B1(new_n569), .B2(new_n790), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n792), .A2(new_n202), .B1(new_n797), .B2(new_n838), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G77), .B2(new_n811), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n786), .A2(G159), .B1(new_n796), .B2(G97), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n305), .A2(new_n809), .B1(new_n806), .B2(G68), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G116), .A2(new_n796), .B1(new_n798), .B2(G326), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n790), .ZN(new_n1040));
  INV_X1    g0840(.A(G283), .ZN(new_n1041));
  INV_X1    g0841(.A(G294), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1040), .A2(new_n1041), .B1(new_n774), .B2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n786), .A2(G322), .B1(new_n806), .B2(G303), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n783), .B2(new_n780), .C1(new_n997), .C2(new_n792), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT110), .Z(new_n1046));
  AOI21_X1  g0846(.A(new_n1043), .B1(new_n1046), .B2(KEYINPUT48), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(KEYINPUT48), .B2(new_n1046), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT49), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n763), .B(new_n1039), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1038), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1032), .B1(new_n1052), .B2(new_n760), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n684), .B2(new_n816), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1020), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n984), .A2(new_n692), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n746), .B2(new_n1018), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(G393));
  INV_X1    g0858(.A(new_n984), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n685), .B1(new_n968), .B2(new_n973), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n975), .A2(new_n967), .A3(new_n960), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n691), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n987), .B2(new_n988), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n974), .A2(new_n976), .A3(new_n991), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n761), .B1(new_n500), .B2(new_n213), .C1(new_n1024), .C2(new_n244), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n752), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT111), .Z(new_n1068));
  OAI22_X1  g0868(.A1(new_n785), .A2(new_n997), .B1(new_n792), .B2(new_n783), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT52), .Z(new_n1070));
  OAI21_X1  g0870(.A(new_n321), .B1(new_n795), .B2(new_n436), .ZN(new_n1071));
  INV_X1    g0871(.A(G322), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n782), .A2(new_n1042), .B1(new_n797), .B2(new_n1072), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(G283), .C2(new_n811), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT113), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n1040), .A2(new_n494), .B1(new_n780), .B2(new_n775), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1070), .B(new_n1077), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G87), .A2(new_n796), .B1(new_n798), .B2(new_n1009), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n764), .B(new_n1079), .C1(new_n311), .C2(new_n774), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT112), .Z(new_n1081));
  AOI22_X1  g0881(.A1(G150), .A2(new_n786), .B1(new_n793), .B2(G159), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT51), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1040), .A2(new_n272), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n780), .A2(new_n202), .B1(new_n782), .B2(new_n258), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1078), .B1(new_n1081), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT114), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n760), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1087), .A2(KEYINPUT114), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1068), .B1(new_n943), .B2(new_n816), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1065), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(KEYINPUT115), .B1(new_n1064), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT115), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1092), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n989), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1094), .B(new_n1095), .C1(new_n1096), .C2(new_n1063), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1093), .A2(new_n1097), .ZN(G390));
  INV_X1    g0898(.A(new_n872), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n912), .A2(new_n1099), .A3(G330), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n662), .A2(new_n679), .A3(new_n824), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n917), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n920), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n923), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n929), .A2(new_n930), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n718), .B1(new_n528), .B2(new_n714), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n650), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n679), .B(new_n824), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n920), .B1(new_n1108), .B2(new_n917), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n923), .B(KEYINPUT116), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n900), .B2(new_n909), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1100), .B1(new_n1105), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(KEYINPUT117), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n889), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n391), .B2(new_n402), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT38), .B1(new_n1117), .B2(new_n886), .ZN(new_n1118));
  OAI21_X1  g0918(.A(KEYINPUT39), .B1(new_n1118), .B2(new_n900), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n927), .A2(new_n928), .A3(new_n894), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n919), .A2(new_n920), .B1(new_n434), .B2(new_n676), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1110), .B1(new_n927), .B2(new_n894), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n918), .B1(new_n721), .B2(new_n824), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n920), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT117), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n1127), .A3(new_n1100), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT118), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n743), .A2(new_n1099), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1122), .A2(new_n1125), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1122), .A2(new_n1125), .A3(new_n1130), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(KEYINPUT118), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1115), .A2(new_n1128), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n991), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n751), .B1(new_n258), .B2(new_n850), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n760), .ZN(new_n1137));
  INV_X1    g0937(.A(G128), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n785), .A2(new_n1138), .B1(new_n782), .B2(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G132), .A2(new_n793), .B1(new_n798), .B2(G125), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n1005), .B2(new_n780), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(G159), .C2(new_n790), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n811), .A2(G150), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT53), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n270), .B1(new_n795), .B2(new_n202), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1146), .A2(KEYINPUT120), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1146), .A2(KEYINPUT120), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n436), .A2(new_n780), .B1(new_n792), .B2(new_n494), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n782), .A2(new_n500), .B1(new_n797), .B2(new_n1042), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n843), .B1(new_n1041), .B2(new_n785), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n321), .B1(new_n774), .B2(new_n563), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n1153), .A2(new_n1084), .A3(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1143), .A2(new_n1149), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1136), .B1(new_n1137), .B2(new_n1156), .C1(new_n1157), .C2(new_n758), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1135), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1134), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n466), .A2(G330), .A3(new_n912), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n935), .A2(new_n670), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n912), .A2(G330), .A3(new_n824), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n920), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1165), .A2(KEYINPUT119), .A3(new_n1124), .A4(new_n1130), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1103), .B1(new_n743), .B2(new_n824), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1102), .B1(new_n1167), .B2(new_n1100), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1167), .A2(new_n1100), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT119), .B1(new_n1170), .B2(new_n1124), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1163), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n692), .B1(new_n1160), .B2(new_n1172), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT119), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1165), .A2(new_n1130), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1124), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1162), .B1(new_n1174), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1133), .A2(new_n1131), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1128), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1127), .B1(new_n1126), .B2(new_n1100), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1179), .B(new_n1180), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1159), .B1(new_n1173), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(G378));
  INV_X1    g0985(.A(new_n910), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n678), .B(new_n1186), .C1(new_n897), .C2(new_n898), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n674), .B1(new_n267), .B2(new_n268), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n303), .B(new_n1188), .Z(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n932), .B1(new_n1157), .B2(new_n923), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n1192), .B2(new_n922), .ZN(new_n1193));
  AND4_X1   g0993(.A1(new_n922), .A2(new_n931), .A3(new_n1191), .A4(new_n933), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1187), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1191), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n934), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n899), .A2(G330), .A3(new_n910), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1192), .A2(new_n922), .A3(new_n1191), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  AOI221_X4 g1000(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1200), .C1(new_n1183), .C2(new_n1163), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT57), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1183), .A2(new_n1163), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1195), .A2(new_n1200), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n691), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n751), .B1(new_n202), .B2(new_n850), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n774), .A2(new_n272), .B1(new_n795), .B2(new_n310), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n763), .A2(new_n279), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(G283), .C2(new_n798), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT122), .Z(new_n1211));
  OAI22_X1  g1011(.A1(new_n780), .A2(new_n500), .B1(new_n782), .B2(new_n447), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT123), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G116), .A2(new_n786), .B1(new_n793), .B2(G107), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n1011), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n317), .B(new_n279), .C1(new_n795), .C2(new_n801), .ZN(new_n1218));
  INV_X1    g1018(.A(G125), .ZN(new_n1219));
  INV_X1    g1019(.A(G132), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n785), .A2(new_n1219), .B1(new_n780), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1139), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1222), .A2(new_n811), .B1(new_n793), .B2(G128), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1005), .B2(new_n782), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1221), .B(new_n1224), .C1(G150), .C2(new_n790), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1218), .B(new_n1227), .C1(G124), .C2(new_n798), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(KEYINPUT59), .B2(new_n1226), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1209), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT121), .ZN(new_n1232));
  AND4_X1   g1032(.A1(new_n1217), .A2(new_n1229), .A3(new_n1230), .A4(new_n1232), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1207), .B1(new_n1137), .B2(new_n1233), .C1(new_n1196), .C2(new_n758), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1204), .B2(new_n991), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1206), .A2(new_n1236), .ZN(G375));
  NAND2_X1  g1037(.A1(new_n920), .A2(new_n757), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n494), .A2(new_n780), .B1(new_n792), .B2(new_n1041), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n270), .B(new_n1239), .C1(G77), .C2(new_n796), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n569), .A2(new_n790), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G97), .A2(new_n811), .B1(new_n798), .B2(G303), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n786), .A2(G294), .B1(new_n806), .B2(G107), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n763), .B1(G50), .B2(new_n790), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n785), .A2(new_n1220), .B1(new_n792), .B2(new_n1005), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G159), .B2(new_n811), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G58), .A2(new_n796), .B1(new_n806), .B2(G150), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n809), .A2(new_n1222), .B1(new_n798), .B2(G128), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1245), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1137), .B1(new_n1244), .B2(new_n1250), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n751), .B(new_n1251), .C1(new_n311), .C2(new_n850), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1238), .A2(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n991), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1253), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1174), .A2(new_n1162), .A3(new_n1178), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n963), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1172), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1257), .A2(new_n1260), .ZN(G381));
  NAND3_X1  g1061(.A1(new_n1206), .A2(new_n1184), .A3(new_n1236), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n992), .A2(new_n1093), .A3(new_n1016), .A4(new_n1097), .ZN(new_n1263));
  INV_X1    g1063(.A(G396), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1055), .A2(new_n1264), .A3(new_n1057), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1265), .A2(G384), .ZN(new_n1266));
  OR4_X1    g1066(.A1(G381), .A2(new_n1262), .A3(new_n1263), .A4(new_n1266), .ZN(G407));
  INV_X1    g1067(.A(G213), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1268), .A2(G343), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1262), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(G407), .A2(new_n1271), .A3(G213), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(KEYINPUT124), .ZN(G409));
  NAND3_X1  g1073(.A1(new_n1206), .A2(G378), .A3(new_n1236), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1203), .A2(new_n1259), .A3(new_n1204), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1236), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1184), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1269), .B1(new_n1274), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1258), .A2(KEYINPUT60), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1254), .A2(new_n1280), .A3(new_n1162), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1172), .A2(new_n691), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1285), .A2(new_n1286), .A3(G384), .A4(new_n1257), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1283), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n830), .B(new_n852), .C1(new_n1288), .C2(new_n1256), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1288), .A2(new_n1256), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1286), .B1(new_n1291), .B2(G384), .ZN(new_n1292));
  INV_X1    g1092(.A(G2897), .ZN(new_n1293));
  OAI22_X1  g1093(.A1(new_n1290), .A2(new_n1292), .B1(new_n1293), .B2(new_n1270), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1285), .A2(G384), .A3(new_n1257), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(KEYINPUT125), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1270), .A2(new_n1293), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1296), .A2(new_n1287), .A3(new_n1289), .A4(new_n1297), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1294), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT63), .B1(new_n1278), .B2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1162), .B1(new_n1134), .B2(new_n1179), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1195), .A2(new_n1200), .ZN(new_n1303));
  OAI21_X1  g1103(.A(KEYINPUT57), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1203), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n692), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1236), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1306), .A2(new_n1184), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1277), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1270), .B(new_n1301), .C1(new_n1308), .C2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1300), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(G393), .A2(G396), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1265), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT126), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1313), .A2(KEYINPUT126), .A3(new_n1265), .ZN(new_n1317));
  AND4_X1   g1117(.A1(new_n992), .A2(new_n1093), .A3(new_n1016), .A4(new_n1097), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n992), .A2(new_n1016), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1316), .B(new_n1317), .C1(new_n1318), .C2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G387), .A2(G390), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1321), .A2(new_n1315), .A3(new_n1263), .A4(new_n1314), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1278), .A2(KEYINPUT63), .A3(new_n1301), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1311), .A2(new_n1312), .A3(new_n1324), .A4(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1310), .A2(new_n1327), .A3(KEYINPUT62), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT62), .B1(new_n1310), .B2(new_n1327), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1312), .B1(new_n1278), .B2(new_n1299), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1328), .A2(new_n1329), .A3(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1326), .B1(new_n1331), .B2(new_n1324), .ZN(G405));
  NAND2_X1  g1132(.A1(G375), .A2(G378), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1262), .ZN(new_n1334));
  AND2_X1   g1134(.A1(new_n1323), .A2(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1323), .A2(new_n1334), .ZN(new_n1336));
  OAI22_X1  g1136(.A1(new_n1335), .A2(new_n1336), .B1(new_n1292), .B2(new_n1290), .ZN(new_n1337));
  OR2_X1    g1137(.A1(new_n1323), .A2(new_n1334), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1323), .A2(new_n1334), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1338), .A2(new_n1301), .A3(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1337), .A2(new_n1340), .ZN(G402));
endmodule


