//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT72), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT0), .A2(G128), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G146), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n192), .A2(KEYINPUT64), .A3(G143), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n191), .B(new_n193), .C1(new_n196), .C2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n193), .A2(new_n199), .ZN(new_n200));
  OR2_X1    g014(.A1(KEYINPUT0), .A2(G128), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n190), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G137), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(G134), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI211_X1 g026(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n204), .C2(G134), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n208), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G131), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n208), .B(new_n216), .C1(new_n212), .C2(new_n213), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n203), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n193), .B(new_n220), .C1(new_n196), .C2(new_n197), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n222), .B1(G143), .B2(new_n192), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n200), .B1(new_n223), .B2(new_n219), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n210), .A2(new_n207), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n225), .A2(new_n217), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n218), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G113), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT2), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT2), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G113), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G116), .B(G119), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT28), .B1(new_n229), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT28), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n195), .A2(G146), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT64), .B1(new_n192), .B2(G143), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n194), .A2(new_n195), .A3(G146), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n201), .A2(new_n190), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n243), .A2(new_n191), .B1(new_n244), .B2(new_n200), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n205), .A2(new_n207), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n211), .B1(new_n206), .B2(G137), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT65), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n210), .A2(new_n209), .A3(new_n211), .ZN(new_n249));
  AOI211_X1 g063(.A(G131), .B(new_n246), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n249), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n216), .B1(new_n251), .B2(new_n208), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n245), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n225), .A2(new_n217), .A3(new_n227), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n237), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n239), .B1(new_n255), .B2(KEYINPUT71), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n236), .B1(new_n218), .B2(new_n228), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n253), .A2(new_n237), .A3(new_n254), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n238), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(KEYINPUT66), .A2(G953), .ZN(new_n264));
  NOR2_X1   g078(.A1(KEYINPUT66), .A2(G953), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G237), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(G210), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(G101), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n268), .A2(new_n269), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n263), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n272), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(new_n262), .A3(new_n270), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n276), .B(KEYINPUT70), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n189), .B1(new_n261), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n238), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT28), .B1(new_n257), .B2(new_n258), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n277), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(KEYINPUT72), .A3(new_n283), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n218), .A2(new_n228), .A3(KEYINPUT30), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT30), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n253), .B2(new_n254), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n236), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n259), .A2(new_n276), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT68), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n259), .A2(new_n292), .A3(new_n276), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n288), .A2(new_n290), .A3(new_n291), .A4(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT69), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n288), .A2(new_n290), .A3(new_n293), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT31), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n278), .A2(new_n284), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n295), .A3(KEYINPUT31), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n188), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n282), .A2(new_n283), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n304));
  INV_X1    g118(.A(new_n259), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT30), .B1(new_n218), .B2(new_n228), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n253), .A2(new_n286), .A3(new_n254), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n305), .B1(new_n308), .B2(new_n236), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n304), .B1(new_n309), .B2(new_n276), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n302), .B1(new_n303), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT28), .B1(new_n305), .B2(new_n255), .ZN(new_n312));
  INV_X1    g126(.A(new_n276), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(new_n304), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n279), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n312), .A2(new_n279), .A3(KEYINPUT76), .A4(new_n314), .ZN(new_n318));
  AOI21_X1  g132(.A(G902), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OR2_X1    g133(.A1(new_n309), .A2(new_n276), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n261), .A2(new_n277), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT75), .A4(new_n304), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n311), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n301), .A2(KEYINPUT32), .B1(G472), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n284), .A2(new_n278), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n296), .A2(new_n298), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n300), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n187), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT73), .B(KEYINPUT32), .Z(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n325), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  AOI211_X1 g146(.A(KEYINPUT74), .B(new_n330), .C1(new_n328), .C2(new_n187), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n324), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G217), .ZN(new_n335));
  INV_X1    g149(.A(G902), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n335), .B1(G234), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G110), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT24), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT24), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G110), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n219), .A2(G119), .ZN(new_n342));
  INV_X1    g156(.A(G119), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(G128), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n339), .B(new_n341), .C1(new_n342), .C2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n343), .B2(G128), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n219), .A2(KEYINPUT23), .A3(G119), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(G128), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n338), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(KEYINPUT78), .ZN(new_n352));
  INV_X1    g166(.A(G140), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G125), .ZN(new_n354));
  INV_X1    g168(.A(G125), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G140), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n356), .A3(KEYINPUT16), .ZN(new_n357));
  OR3_X1    g171(.A1(new_n355), .A2(KEYINPUT16), .A3(G140), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(G146), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT79), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n357), .A2(new_n358), .A3(new_n361), .A4(G146), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n354), .A2(new_n356), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n192), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n360), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n352), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n347), .A2(new_n349), .A3(new_n348), .ZN(new_n367));
  XNOR2_X1  g181(.A(G119), .B(G128), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n339), .A2(new_n341), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n367), .A2(G110), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n357), .A2(G146), .A3(new_n358), .ZN(new_n371));
  AOI21_X1  g185(.A(G146), .B1(new_n357), .B2(new_n358), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT77), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n370), .B(new_n375), .C1(new_n371), .C2(new_n372), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n266), .A2(G221), .A3(G234), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT22), .B(G137), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n378), .B(new_n379), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n366), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n380), .B1(new_n366), .B2(new_n377), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT25), .B1(new_n383), .B2(new_n336), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n366), .A2(new_n377), .ZN(new_n385));
  INV_X1    g199(.A(new_n380), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n366), .A2(new_n377), .A3(new_n380), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n387), .A2(KEYINPUT25), .A3(new_n336), .A4(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n337), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n337), .A2(G902), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n383), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n337), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n387), .A2(new_n336), .A3(new_n388), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT25), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n396), .B1(new_n399), .B2(new_n389), .ZN(new_n400));
  INV_X1    g214(.A(new_n394), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT80), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(G210), .B1(G237), .B2(G902), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n355), .B1(new_n198), .B2(new_n202), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n221), .A2(new_n224), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n407), .B1(new_n355), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G224), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT7), .B1(new_n410), .B2(G953), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n234), .A2(new_n235), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n343), .A2(G116), .ZN(new_n414));
  INV_X1    g228(.A(G116), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G119), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n414), .A2(new_n416), .A3(KEYINPUT5), .ZN(new_n417));
  OAI21_X1  g231(.A(G113), .B1(new_n414), .B2(KEYINPUT5), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n413), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G104), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT3), .B1(new_n420), .B2(G107), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT3), .ZN(new_n422));
  INV_X1    g236(.A(G107), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(G104), .ZN(new_n424));
  INV_X1    g238(.A(G101), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n420), .A2(G107), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n421), .A2(new_n424), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n420), .A2(G107), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n423), .A2(G104), .ZN(new_n429));
  OAI21_X1  g243(.A(G101), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n419), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n414), .A2(new_n416), .A3(KEYINPUT5), .ZN(new_n433));
  OR3_X1    g247(.A1(new_n415), .A2(KEYINPUT5), .A3(G119), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(G113), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n435), .A2(new_n413), .A3(new_n427), .A4(new_n430), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G122), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n338), .A2(G122), .ZN(new_n441));
  INV_X1    g255(.A(G122), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(G110), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT85), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n440), .A2(new_n444), .A3(KEYINPUT8), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT8), .B1(new_n440), .B2(new_n444), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n409), .A2(new_n412), .B1(new_n437), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT87), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n221), .A2(new_n355), .A3(new_n224), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n245), .B2(new_n355), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT86), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n411), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n451), .B2(new_n411), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n448), .B(new_n449), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n421), .A2(new_n424), .A3(new_n426), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G101), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(KEYINPUT4), .A3(new_n427), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT4), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n460), .A3(G101), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n236), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n440), .A2(new_n444), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n436), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n456), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n455), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n453), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n449), .B1(new_n467), .B2(new_n448), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n462), .A2(new_n436), .ZN(new_n470));
  INV_X1    g284(.A(new_n463), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(KEYINPUT6), .A3(new_n464), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n474), .A3(new_n471), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n410), .A2(G953), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n451), .B(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n336), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n406), .B1(new_n469), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n478), .A2(new_n336), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n454), .A2(new_n455), .ZN(new_n482));
  INV_X1    g296(.A(new_n448), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT87), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(new_n464), .A3(new_n456), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n485), .A3(new_n405), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n427), .A2(new_n430), .ZN(new_n488));
  INV_X1    g302(.A(new_n221), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n223), .A2(new_n219), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n243), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n488), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n215), .A2(new_n217), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n459), .A2(new_n245), .A3(new_n461), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n225), .A2(new_n488), .A3(KEYINPUT10), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n495), .A2(new_n497), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n225), .A2(new_n488), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n193), .B1(new_n196), .B2(new_n197), .ZN(new_n502));
  OAI21_X1  g316(.A(G128), .B1(new_n240), .B2(new_n222), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n431), .B1(new_n504), .B2(new_n221), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n496), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT12), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT12), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n508), .B(new_n496), .C1(new_n501), .C2(new_n505), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n500), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT83), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n266), .A2(G227), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT81), .ZN(new_n513));
  XNOR2_X1  g327(.A(G110), .B(G140), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT83), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n500), .A2(new_n507), .A3(new_n517), .A4(new_n509), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n511), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n499), .B1(new_n505), .B2(new_n493), .ZN(new_n520));
  INV_X1    g334(.A(new_n498), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n496), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n500), .A3(new_n515), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n519), .A2(G469), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n500), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n516), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n500), .A2(new_n507), .A3(new_n515), .A4(new_n509), .ZN(new_n527));
  AOI21_X1  g341(.A(G902), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G469), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n336), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n524), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT9), .B(G234), .ZN(new_n534));
  OAI21_X1  g348(.A(G221), .B1(new_n534), .B2(G902), .ZN(new_n535));
  INV_X1    g349(.A(new_n266), .ZN(new_n536));
  NAND2_X1  g350(.A1(G234), .A2(G237), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(G902), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT21), .B(G898), .ZN(new_n540));
  INV_X1    g354(.A(G952), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(G953), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n539), .A2(new_n540), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(G214), .B1(G237), .B2(G902), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n545), .B(KEYINPUT84), .Z(new_n546));
  AND2_X1   g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n487), .A2(new_n533), .A3(new_n535), .A4(new_n547), .ZN(new_n548));
  XOR2_X1   g362(.A(G113), .B(G122), .Z(new_n549));
  XOR2_X1   g363(.A(KEYINPUT88), .B(G104), .Z(new_n550));
  XOR2_X1   g364(.A(new_n549), .B(new_n550), .Z(new_n551));
  AND3_X1   g365(.A1(new_n354), .A2(new_n356), .A3(KEYINPUT19), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT19), .B1(new_n354), .B2(new_n356), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n192), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n360), .A2(new_n362), .A3(new_n554), .ZN(new_n555));
  OR2_X1    g369(.A1(KEYINPUT66), .A2(G953), .ZN(new_n556));
  NAND2_X1  g370(.A1(KEYINPUT66), .A2(G953), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n556), .A2(G214), .A3(new_n267), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n195), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n266), .A2(G143), .A3(G214), .A4(new_n267), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n216), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n560), .A3(new_n216), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n555), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n559), .A2(new_n560), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT18), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(new_n216), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n363), .B(new_n192), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n559), .B(new_n560), .C1(new_n566), .C2(new_n216), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n551), .B1(new_n564), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n573));
  INV_X1    g387(.A(new_n551), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n559), .A2(new_n560), .A3(new_n216), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n575), .A2(new_n561), .A3(KEYINPUT17), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n565), .A2(KEYINPUT17), .A3(G131), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n371), .A2(new_n372), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n573), .B(new_n574), .C1(new_n576), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(G475), .A2(G902), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT20), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT20), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n581), .A2(new_n585), .A3(new_n582), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n573), .B1(new_n576), .B2(new_n579), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n588), .A2(new_n551), .ZN(new_n589));
  INV_X1    g403(.A(new_n580), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n336), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G475), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n534), .A2(new_n335), .A3(G953), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT94), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT89), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n442), .B2(G116), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n415), .A2(KEYINPUT89), .A3(G122), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n442), .A2(G116), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n423), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n219), .A2(G143), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n195), .A2(KEYINPUT90), .A3(G128), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT90), .B1(new_n195), .B2(G128), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n206), .B(new_n603), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT90), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n219), .B2(G143), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n195), .A2(KEYINPUT90), .A3(G128), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n206), .B1(new_n611), .B2(new_n603), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n602), .B1(new_n607), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT14), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n598), .A2(new_n614), .A3(new_n599), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT93), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n615), .A2(new_n616), .B1(G116), .B2(new_n442), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n598), .A2(new_n599), .A3(KEYINPUT93), .A4(new_n614), .ZN(new_n618));
  AOI211_X1 g432(.A(KEYINPUT92), .B(new_n614), .C1(new_n598), .C2(new_n599), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT92), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n600), .B2(KEYINPUT14), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n613), .B1(new_n622), .B2(G107), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n606), .A2(KEYINPUT91), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT91), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n611), .A2(new_n625), .A3(new_n206), .A4(new_n603), .ZN(new_n626));
  INV_X1    g440(.A(new_n602), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n423), .B1(new_n600), .B2(new_n601), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n624), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT13), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n611), .A2(new_n630), .B1(new_n219), .B2(G143), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n609), .A2(KEYINPUT13), .A3(new_n610), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n206), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n596), .B1(new_n623), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n621), .A2(new_n619), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n615), .A2(new_n616), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n618), .A3(new_n601), .ZN(new_n638));
  OAI21_X1  g452(.A(G107), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n613), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n631), .A2(new_n632), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(G134), .ZN(new_n643));
  INV_X1    g457(.A(new_n628), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n602), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n643), .A2(new_n645), .A3(new_n626), .A4(new_n624), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n641), .A2(new_n646), .A3(new_n595), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n635), .A2(new_n647), .A3(KEYINPUT95), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT95), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n641), .A2(new_n646), .A3(new_n649), .A4(new_n595), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n648), .A2(new_n336), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(G478), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(KEYINPUT15), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n653), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n648), .A2(new_n336), .A3(new_n650), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT96), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n654), .A2(KEYINPUT96), .A3(new_n656), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n593), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n548), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n334), .A2(new_n404), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT97), .B(G101), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G3));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n651), .A2(new_n652), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n595), .B1(new_n641), .B2(new_n646), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT98), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n668), .B1(new_n669), .B2(new_n647), .ZN(new_n670));
  AOI211_X1 g484(.A(KEYINPUT98), .B(new_n595), .C1(new_n641), .C2(new_n646), .ZN(new_n671));
  OAI21_X1  g485(.A(KEYINPUT33), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n648), .A2(new_n650), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT33), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n652), .A2(G902), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n667), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n666), .B1(new_n678), .B2(new_n593), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n647), .A2(new_n669), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n635), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n668), .A2(new_n669), .A3(new_n647), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n674), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(KEYINPUT33), .B1(new_n648), .B2(new_n650), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n677), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n651), .A2(new_n652), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n587), .A2(new_n592), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(KEYINPUT99), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n679), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n545), .ZN(new_n691));
  AOI211_X1 g505(.A(new_n691), .B(new_n543), .C1(new_n480), .C2(new_n486), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n690), .A2(KEYINPUT100), .A3(new_n692), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n535), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n531), .B1(new_n528), .B2(new_n529), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n698), .B1(new_n699), .B2(new_n524), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n395), .A3(new_n402), .ZN(new_n701));
  INV_X1    g515(.A(G472), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n328), .B2(new_n336), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n701), .A2(new_n703), .A3(new_n301), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n697), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT34), .B(G104), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G6));
  NAND2_X1  g521(.A1(new_n659), .A2(new_n660), .ZN(new_n708));
  MUX2_X1   g522(.A(new_n584), .B(new_n587), .S(KEYINPUT101), .Z(new_n709));
  AND4_X1   g523(.A1(new_n592), .A2(new_n692), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n704), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT35), .B(G107), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G9));
  NOR2_X1   g527(.A1(new_n386), .A2(KEYINPUT36), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n385), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n366), .A3(new_n377), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n393), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT102), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n716), .A2(new_n720), .A3(new_n393), .A4(new_n717), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n400), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n548), .A2(new_n661), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n703), .A2(new_n301), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT37), .B(G110), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G12));
  NAND2_X1  g542(.A1(new_n542), .A2(new_n537), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n729), .B(KEYINPUT103), .Z(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(G900), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n731), .B1(new_n539), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n591), .B2(G475), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n708), .A2(new_n709), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n723), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n691), .B1(new_n480), .B2(new_n486), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n737), .A3(new_n700), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n334), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G128), .ZN(G30));
  NAND2_X1  g555(.A1(new_n533), .A2(new_n535), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n733), .B(KEYINPUT39), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT40), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(KEYINPUT40), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n487), .B(KEYINPUT38), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n708), .A2(new_n688), .ZN(new_n749));
  NOR4_X1   g563(.A1(new_n748), .A2(new_n691), .A3(new_n736), .A4(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n305), .A2(new_n255), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n297), .B1(new_n277), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n702), .B1(new_n752), .B2(new_n336), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n301), .B2(KEYINPUT32), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n332), .B2(new_n333), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n750), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G143), .ZN(G45));
  INV_X1    g571(.A(new_n733), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n687), .A2(new_n688), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n738), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n334), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G146), .ZN(G48));
  OR2_X1    g576(.A1(new_n528), .A2(new_n529), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n763), .A2(new_n535), .A3(new_n530), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n404), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT100), .B1(new_n690), .B2(new_n692), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n469), .A2(new_n406), .A3(new_n479), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n405), .B1(new_n481), .B2(new_n485), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n545), .B(new_n544), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  AOI211_X1 g584(.A(new_n694), .B(new_n770), .C1(new_n679), .C2(new_n689), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n334), .B(new_n766), .C1(new_n767), .C2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT41), .B(G113), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G15));
  NAND3_X1  g588(.A1(new_n334), .A2(new_n710), .A3(new_n766), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G116), .ZN(G18));
  NAND3_X1  g590(.A1(new_n764), .A2(new_n737), .A3(new_n736), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n777), .A2(new_n661), .A3(new_n543), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n334), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G119), .ZN(G21));
  INV_X1    g594(.A(KEYINPUT104), .ZN(new_n781));
  AOI21_X1  g595(.A(G902), .B1(new_n299), .B2(new_n300), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n781), .B1(new_n782), .B2(new_n702), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n703), .A2(KEYINPUT104), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AND4_X1   g599(.A1(new_n688), .A2(new_n692), .A3(new_n708), .A4(new_n764), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n391), .A2(new_n394), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n312), .A2(new_n279), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n298), .B1(new_n789), .B2(new_n277), .ZN(new_n790));
  INV_X1    g604(.A(new_n294), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n187), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n785), .A2(new_n786), .A3(new_n788), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G122), .ZN(G24));
  NOR2_X1   g608(.A1(new_n777), .A2(new_n759), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n785), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G125), .ZN(G27));
  NAND3_X1  g611(.A1(new_n480), .A2(new_n486), .A3(new_n545), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n523), .A2(KEYINPUT105), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n523), .A2(KEYINPUT105), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n519), .A2(G469), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n698), .B1(new_n699), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n759), .ZN(new_n805));
  INV_X1    g619(.A(new_n324), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n301), .A2(KEYINPUT32), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n805), .B(new_n788), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT74), .B1(new_n301), .B2(new_n330), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n329), .A2(new_n325), .A3(new_n331), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n403), .B1(new_n811), .B2(new_n324), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n804), .A2(KEYINPUT42), .A3(new_n759), .ZN(new_n813));
  AOI22_X1  g627(.A1(KEYINPUT42), .A2(new_n808), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G131), .ZN(G33));
  NOR2_X1   g629(.A1(new_n735), .A2(new_n804), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n334), .A2(new_n404), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT106), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n334), .A2(KEYINPUT106), .A3(new_n404), .A4(new_n816), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G134), .ZN(G36));
  NAND4_X1  g636(.A1(new_n519), .A2(KEYINPUT45), .A3(new_n800), .A4(new_n801), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(G469), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT45), .B1(new_n519), .B2(new_n523), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT46), .B1(new_n826), .B2(new_n532), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n529), .B2(new_n528), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n826), .A2(KEYINPUT46), .A3(new_n532), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n698), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n743), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n678), .A2(new_n688), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT43), .Z(new_n834));
  NOR3_X1   g648(.A1(new_n834), .A2(new_n725), .A3(new_n723), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n798), .B1(new_n835), .B2(KEYINPUT44), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n832), .B(new_n836), .C1(KEYINPUT44), .C2(new_n835), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(G137), .ZN(G39));
  XOR2_X1   g652(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n839));
  NOR2_X1   g653(.A1(new_n830), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n840), .B1(new_n830), .B2(new_n841), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n334), .A2(new_n404), .A3(new_n759), .A4(new_n798), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(G140), .ZN(G42));
  NAND2_X1  g659(.A1(new_n799), .A2(new_n764), .ZN(new_n846));
  OR3_X1    g660(.A1(new_n834), .A2(new_n730), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n788), .B1(new_n806), .B2(new_n807), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT113), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT48), .ZN(new_n852));
  XNOR2_X1  g666(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n834), .A2(new_n730), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n785), .A2(new_n792), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n855), .A2(new_n788), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n737), .A3(new_n764), .ZN(new_n858));
  INV_X1    g672(.A(new_n690), .ZN(new_n859));
  OR4_X1    g673(.A1(new_n403), .A2(new_n755), .A3(new_n729), .A4(new_n846), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n858), .B(new_n542), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n852), .A2(new_n854), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n763), .A2(new_n530), .ZN(new_n863));
  NOR4_X1   g677(.A1(new_n747), .A2(new_n698), .A3(new_n545), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT50), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n856), .A2(new_n736), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n847), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n860), .A2(new_n688), .A3(new_n687), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n698), .B1(new_n863), .B2(KEYINPUT111), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(KEYINPUT111), .B2(new_n863), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n799), .B(new_n857), .C1(new_n842), .C2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n870), .A2(KEYINPUT51), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n862), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT112), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n873), .A2(new_n877), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n870), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n875), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n772), .A2(new_n775), .A3(new_n779), .A4(new_n793), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n547), .B1(new_n768), .B2(new_n769), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n687), .A2(new_n688), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n593), .A2(new_n657), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n704), .A2(new_n886), .B1(new_n724), .B2(new_n725), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n785), .A2(new_n805), .A3(new_n736), .A4(new_n792), .ZN(new_n888));
  INV_X1    g702(.A(new_n657), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n709), .A2(new_n736), .A3(new_n889), .A4(new_n734), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n890), .A2(new_n742), .A3(new_n798), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n334), .A2(new_n891), .ZN(new_n892));
  AND4_X1   g706(.A1(new_n663), .A2(new_n887), .A3(new_n888), .A4(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n882), .A2(new_n814), .A3(new_n821), .A4(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n332), .A2(new_n333), .ZN(new_n895));
  OAI22_X1  g709(.A1(new_n895), .A2(new_n806), .B1(new_n739), .B2(new_n760), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n400), .A2(new_n722), .A3(new_n733), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT108), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n803), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n708), .A2(new_n688), .A3(new_n737), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n898), .B1(new_n803), .B2(new_n897), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n755), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n896), .A2(new_n903), .A3(KEYINPUT52), .A4(new_n796), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n894), .B1(new_n905), .B2(KEYINPUT109), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n896), .A2(new_n796), .A3(new_n903), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT52), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT109), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n910), .A3(new_n904), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT53), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n821), .A2(new_n814), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n909), .A2(new_n904), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(new_n917), .A3(new_n882), .A4(new_n893), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n914), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT54), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n909), .A2(new_n904), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n913), .B1(new_n894), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT110), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n765), .B1(new_n811), .B2(new_n324), .ZN(new_n926));
  AOI22_X1  g740(.A1(new_n697), .A2(new_n926), .B1(new_n334), .B2(new_n778), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n775), .A2(new_n793), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n700), .A2(new_n395), .A3(new_n402), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n328), .A2(new_n336), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(G472), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n886), .A2(new_n329), .A3(new_n929), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n726), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n812), .B2(new_n662), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n888), .A2(new_n892), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n927), .A2(new_n928), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n915), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n905), .A2(KEYINPUT109), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n937), .A2(KEYINPUT53), .A3(new_n911), .A4(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(KEYINPUT110), .B(new_n913), .C1(new_n894), .C2(new_n921), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n924), .A2(new_n925), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n881), .A2(new_n920), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(G952), .B2(G953), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n788), .A2(new_n535), .A3(new_n546), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n863), .A2(KEYINPUT49), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n863), .A2(KEYINPUT49), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n944), .A2(new_n833), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  OR3_X1    g761(.A1(new_n755), .A2(new_n947), .A3(new_n747), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n943), .A2(new_n948), .ZN(G75));
  AND2_X1   g763(.A1(new_n473), .A2(new_n475), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(new_n477), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT55), .ZN(new_n952));
  XOR2_X1   g766(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n924), .A2(new_n939), .A3(new_n940), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(G902), .ZN(new_n956));
  INV_X1    g770(.A(G210), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n266), .A2(G952), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT56), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n956), .B2(new_n957), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n963), .A2(new_n952), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n964), .A2(KEYINPUT115), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(KEYINPUT115), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n961), .B1(new_n965), .B2(new_n966), .ZN(G51));
  NAND2_X1  g781(.A1(new_n939), .A2(new_n940), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT110), .B1(new_n918), .B2(new_n913), .ZN(new_n969));
  OAI21_X1  g783(.A(KEYINPUT54), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT118), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n971), .A3(new_n941), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n955), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n973));
  XNOR2_X1  g787(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(new_n531), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n526), .A2(new_n527), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n826), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n955), .A2(G902), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n981), .A2(KEYINPUT119), .A3(new_n960), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT119), .ZN(new_n983));
  INV_X1    g797(.A(new_n980), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n976), .B2(new_n977), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n983), .B1(new_n985), .B2(new_n959), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n982), .A2(new_n986), .ZN(G54));
  INV_X1    g801(.A(new_n956), .ZN(new_n988));
  NAND2_X1  g802(.A1(KEYINPUT58), .A2(G475), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT120), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n988), .A2(new_n581), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n581), .B1(new_n988), .B2(new_n990), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n991), .A2(new_n992), .A3(new_n959), .ZN(G60));
  NAND2_X1  g807(.A1(G478), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT59), .Z(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n920), .B2(new_n941), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n676), .B(KEYINPUT121), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n960), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n995), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n972), .A2(new_n973), .A3(new_n999), .A4(new_n997), .ZN(new_n1000));
  OR2_X1    g814(.A1(new_n1000), .A2(KEYINPUT122), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(KEYINPUT122), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(G63));
  NAND2_X1  g817(.A1(G217), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT60), .Z(new_n1005));
  NAND4_X1  g819(.A1(new_n955), .A2(new_n717), .A3(new_n716), .A4(new_n1005), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n955), .A2(new_n1005), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n960), .B(new_n1006), .C1(new_n1007), .C2(new_n383), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g823(.A(G953), .B1(new_n540), .B2(new_n410), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT123), .Z(new_n1011));
  AND2_X1   g825(.A1(new_n882), .A2(new_n934), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1011), .B1(new_n1012), .B2(new_n536), .ZN(new_n1013));
  INV_X1    g827(.A(G898), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n950), .B1(new_n1014), .B2(new_n536), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1013), .B(new_n1015), .Z(G69));
  NOR2_X1   g830(.A1(new_n552), .A2(new_n553), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n308), .B(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1018), .B1(G900), .B2(new_n536), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n844), .A2(new_n837), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n896), .A2(new_n796), .ZN(new_n1021));
  NOR4_X1   g835(.A1(new_n831), .A2(new_n743), .A3(new_n848), .A4(new_n900), .ZN(new_n1022));
  NOR3_X1   g836(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  OR2_X1    g837(.A1(new_n915), .A2(KEYINPUT124), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n915), .A2(KEYINPUT124), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1019), .B1(new_n1026), .B2(new_n536), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n896), .A2(new_n796), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n756), .A2(new_n1028), .ZN(new_n1029));
  AND2_X1   g843(.A1(new_n1029), .A2(KEYINPUT62), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1029), .A2(KEYINPUT62), .ZN(new_n1031));
  OR2_X1    g845(.A1(new_n744), .A2(new_n798), .ZN(new_n1032));
  INV_X1    g846(.A(new_n812), .ZN(new_n1033));
  AOI211_X1 g847(.A(new_n1032), .B(new_n1033), .C1(new_n884), .C2(new_n885), .ZN(new_n1034));
  NOR4_X1   g848(.A1(new_n1030), .A2(new_n1020), .A3(new_n1031), .A4(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1018), .B1(new_n1035), .B2(new_n536), .ZN(new_n1036));
  INV_X1    g850(.A(KEYINPUT126), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1027), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1037), .B1(new_n1027), .B2(new_n1036), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT125), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n1018), .A2(new_n1041), .ZN(new_n1042));
  AOI211_X1 g856(.A(new_n266), .B(new_n1042), .C1(G227), .C2(G900), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1043), .ZN(new_n1044));
  NOR3_X1   g858(.A1(new_n1039), .A2(new_n1040), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1027), .A2(new_n1036), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(KEYINPUT126), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1043), .B1(new_n1047), .B2(new_n1038), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n1045), .A2(new_n1048), .ZN(G72));
  NOR2_X1   g863(.A1(new_n309), .A2(new_n313), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1035), .A2(new_n1012), .ZN(new_n1052));
  NAND2_X1  g866(.A1(G472), .A2(G902), .ZN(new_n1053));
  XOR2_X1   g867(.A(new_n1053), .B(KEYINPUT63), .Z(new_n1054));
  AOI21_X1  g868(.A(new_n1051), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g869(.A(new_n1055), .B(KEYINPUT127), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n320), .A2(new_n297), .ZN(new_n1057));
  NAND3_X1  g871(.A1(new_n919), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  NAND4_X1  g872(.A1(new_n1023), .A2(new_n1012), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1059));
  AND2_X1   g873(.A1(new_n1059), .A2(new_n1054), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n309), .A2(new_n313), .ZN(new_n1061));
  OAI211_X1 g875(.A(new_n960), .B(new_n1058), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g876(.A1(new_n1056), .A2(new_n1062), .ZN(G57));
endmodule


