

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782;

  AND2_X1 U378 ( .A1(n607), .A2(n720), .ZN(n617) );
  AND2_X2 U379 ( .A1(n380), .A2(n608), .ZN(n693) );
  NOR2_X2 U380 ( .A1(n746), .A2(n620), .ZN(n402) );
  NOR2_X1 U381 ( .A1(n669), .A2(G902), .ZN(n442) );
  AND2_X1 U382 ( .A1(n621), .A2(n486), .ZN(n553) );
  XNOR2_X1 U383 ( .A(n597), .B(KEYINPUT0), .ZN(n603) );
  XNOR2_X1 U384 ( .A(n442), .B(n423), .ZN(n609) );
  NOR2_X2 U385 ( .A1(G953), .A2(G237), .ZN(n509) );
  NAND2_X1 U386 ( .A1(n644), .A2(n374), .ZN(n365) );
  NAND2_X1 U387 ( .A1(n364), .A2(n366), .ZN(n374) );
  XNOR2_X1 U388 ( .A(n387), .B(KEYINPUT40), .ZN(n668) );
  XNOR2_X1 U389 ( .A(n421), .B(n619), .ZN(n703) );
  XNOR2_X1 U390 ( .A(n382), .B(n381), .ZN(n782) );
  OR2_X1 U391 ( .A1(n732), .A2(n541), .ZN(n542) );
  NAND2_X1 U392 ( .A1(n553), .A2(n552), .ZN(n386) );
  NAND2_X1 U393 ( .A1(n395), .A2(n393), .ZN(n746) );
  AND2_X1 U394 ( .A1(n398), .A2(n396), .ZN(n395) );
  NOR2_X1 U395 ( .A1(n603), .A2(n602), .ZN(n605) );
  INV_X1 U396 ( .A(n556), .ZN(n727) );
  OR2_X1 U397 ( .A1(n646), .A2(G902), .ZN(n478) );
  INV_X2 U398 ( .A(G107), .ZN(n413) );
  INV_X2 U399 ( .A(G119), .ZN(n416) );
  INV_X2 U400 ( .A(G122), .ZN(n415) );
  XNOR2_X1 U401 ( .A(n415), .B(G104), .ZN(n355) );
  XNOR2_X1 U402 ( .A(n415), .B(G104), .ZN(n503) );
  XNOR2_X1 U403 ( .A(n556), .B(KEYINPUT6), .ZN(n626) );
  BUF_X1 U404 ( .A(n640), .Z(n356) );
  BUF_X1 U405 ( .A(n639), .Z(n640) );
  BUF_X1 U406 ( .A(n522), .Z(n357) );
  XNOR2_X1 U407 ( .A(n605), .B(n604), .ZN(n613) );
  BUF_X1 U408 ( .A(n603), .Z(n620) );
  OR2_X2 U409 ( .A1(n643), .A2(n770), .ZN(n644) );
  NOR2_X1 U410 ( .A1(n613), .A2(n598), .ZN(n625) );
  NAND2_X1 U411 ( .A1(n375), .A2(n373), .ZN(n372) );
  NOR2_X1 U412 ( .A1(n384), .A2(n410), .ZN(n383) );
  NOR2_X2 U413 ( .A1(n782), .A2(n693), .ZN(n616) );
  INV_X1 U414 ( .A(KEYINPUT95), .ZN(n417) );
  NOR2_X1 U415 ( .A1(n361), .A2(n376), .ZN(n375) );
  INV_X1 U416 ( .A(n377), .ZN(n376) );
  INV_X1 U417 ( .A(KEYINPUT92), .ZN(n373) );
  OR2_X1 U418 ( .A1(n626), .A2(n399), .ZN(n398) );
  XNOR2_X1 U419 ( .A(n378), .B(n500), .ZN(n558) );
  INV_X1 U420 ( .A(KEYINPUT16), .ZN(n488) );
  XOR2_X1 U421 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n471) );
  AND2_X1 U422 ( .A1(n727), .A2(n735), .ZN(n480) );
  AND2_X1 U423 ( .A1(n408), .A2(KEYINPUT47), .ZN(n407) );
  AND2_X1 U424 ( .A1(n386), .A2(n568), .ZN(n569) );
  AND2_X1 U425 ( .A1(n383), .A2(n575), .ZN(n576) );
  AND2_X1 U426 ( .A1(n630), .A2(n390), .ZN(n389) );
  INV_X1 U427 ( .A(KEYINPUT10), .ZN(n424) );
  XNOR2_X1 U428 ( .A(G902), .B(KEYINPUT15), .ZN(n635) );
  NOR2_X1 U429 ( .A1(G902), .A2(G237), .ZN(n479) );
  XNOR2_X1 U430 ( .A(G137), .B(KEYINPUT102), .ZN(n466) );
  XNOR2_X1 U431 ( .A(G116), .B(G119), .ZN(n467) );
  XNOR2_X1 U432 ( .A(KEYINPUT5), .B(KEYINPUT82), .ZN(n464) );
  XNOR2_X1 U433 ( .A(G113), .B(G131), .ZN(n504) );
  XNOR2_X1 U434 ( .A(G143), .B(G140), .ZN(n505) );
  XOR2_X1 U435 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n506) );
  XNOR2_X1 U436 ( .A(n427), .B(n426), .ZN(n513) );
  XNOR2_X1 U437 ( .A(G146), .B(G125), .ZN(n427) );
  XNOR2_X1 U438 ( .A(n425), .B(n424), .ZN(n426) );
  INV_X1 U439 ( .A(KEYINPUT71), .ZN(n425) );
  XOR2_X1 U440 ( .A(KEYINPUT78), .B(KEYINPUT17), .Z(n492) );
  XNOR2_X1 U441 ( .A(n535), .B(KEYINPUT73), .ZN(n536) );
  INV_X1 U442 ( .A(G902), .ZN(n514) );
  INV_X1 U443 ( .A(KEYINPUT64), .ZN(n430) );
  XNOR2_X1 U444 ( .A(G134), .B(G122), .ZN(n519) );
  INV_X1 U445 ( .A(n419), .ZN(n367) );
  NAND2_X1 U446 ( .A1(n358), .A2(KEYINPUT92), .ZN(n371) );
  NAND2_X1 U447 ( .A1(n370), .A2(n369), .ZN(n368) );
  NAND2_X1 U448 ( .A1(n358), .A2(n373), .ZN(n369) );
  NAND2_X1 U449 ( .A1(n375), .A2(KEYINPUT92), .ZN(n370) );
  XNOR2_X1 U450 ( .A(G104), .B(G101), .ZN(n450) );
  XNOR2_X1 U451 ( .A(G110), .B(G107), .ZN(n449) );
  XNOR2_X1 U452 ( .A(G137), .B(G140), .ZN(n454) );
  NAND2_X1 U453 ( .A1(G234), .A2(G237), .ZN(n483) );
  NAND2_X1 U454 ( .A1(n394), .A2(n626), .ZN(n393) );
  NAND2_X1 U455 ( .A1(n558), .A2(n735), .ZN(n563) );
  XNOR2_X1 U456 ( .A(n563), .B(KEYINPUT19), .ZN(n596) );
  XNOR2_X1 U457 ( .A(n463), .B(n462), .ZN(n621) );
  XNOR2_X1 U458 ( .A(n414), .B(n412), .ZN(n490) );
  XNOR2_X1 U459 ( .A(n518), .B(n488), .ZN(n412) );
  XNOR2_X1 U460 ( .A(n487), .B(n503), .ZN(n414) );
  XNOR2_X1 U461 ( .A(n403), .B(n768), .ZN(n669) );
  INV_X1 U462 ( .A(G953), .ZN(n756) );
  INV_X1 U463 ( .A(G134), .ZN(n530) );
  INV_X1 U464 ( .A(KEYINPUT32), .ZN(n381) );
  NAND2_X1 U465 ( .A1(n622), .A2(n422), .ZN(n421) );
  INV_X1 U466 ( .A(n729), .ZN(n422) );
  AND2_X1 U467 ( .A1(n377), .A2(n638), .ZN(n358) );
  OR2_X1 U468 ( .A1(n551), .A2(n544), .ZN(n700) );
  AND2_X1 U469 ( .A1(n617), .A2(n399), .ZN(n359) );
  NAND2_X1 U470 ( .A1(n571), .A2(KEYINPUT89), .ZN(n360) );
  AND2_X1 U471 ( .A1(n637), .A2(n638), .ZN(n361) );
  NAND2_X1 U472 ( .A1(n372), .A2(n371), .ZN(n362) );
  XNOR2_X1 U473 ( .A(n764), .B(n379), .ZN(n661) );
  XNOR2_X1 U474 ( .A(n490), .B(n489), .ZN(n764) );
  NAND2_X1 U475 ( .A1(n363), .A2(n418), .ZN(n388) );
  XNOR2_X1 U476 ( .A(n616), .B(n615), .ZN(n363) );
  NAND2_X1 U477 ( .A1(n367), .A2(n362), .ZN(n364) );
  XNOR2_X2 U478 ( .A(n365), .B(n645), .ZN(n677) );
  XNOR2_X1 U479 ( .A(n391), .B(n417), .ZN(n390) );
  NAND2_X1 U480 ( .A1(n419), .A2(n368), .ZN(n366) );
  OR2_X1 U481 ( .A1(n637), .A2(n638), .ZN(n377) );
  NAND2_X1 U482 ( .A1(n661), .A2(n635), .ZN(n378) );
  XNOR2_X1 U483 ( .A(n497), .B(n498), .ZN(n379) );
  XNOR2_X1 U484 ( .A(n625), .B(n606), .ZN(n380) );
  OR2_X1 U485 ( .A1(n614), .A2(n613), .ZN(n382) );
  NAND2_X1 U486 ( .A1(n360), .A2(n385), .ZN(n384) );
  NAND2_X1 U487 ( .A1(n570), .A2(n572), .ZN(n385) );
  NOR2_X1 U488 ( .A1(n386), .A2(n568), .ZN(n555) );
  XNOR2_X1 U489 ( .A(n386), .B(n697), .ZN(G45) );
  NAND2_X1 U490 ( .A1(n529), .A2(n406), .ZN(n387) );
  XNOR2_X1 U491 ( .A(n502), .B(KEYINPUT39), .ZN(n529) );
  NAND2_X1 U492 ( .A1(n389), .A2(n388), .ZN(n632) );
  NAND2_X1 U493 ( .A1(n781), .A2(KEYINPUT44), .ZN(n391) );
  XNOR2_X1 U494 ( .A(n392), .B(n474), .ZN(n646) );
  XNOR2_X1 U495 ( .A(n392), .B(n457), .ZN(n680) );
  XNOR2_X2 U496 ( .A(n769), .B(G146), .ZN(n392) );
  NAND2_X1 U497 ( .A1(n598), .A2(n617), .ZN(n397) );
  XNOR2_X2 U498 ( .A(n560), .B(KEYINPUT1), .ZN(n598) );
  AND2_X1 U499 ( .A1(n598), .A2(n359), .ZN(n394) );
  NAND2_X1 U500 ( .A1(n397), .A2(n599), .ZN(n396) );
  INV_X1 U501 ( .A(n599), .ZN(n399) );
  INV_X1 U502 ( .A(n626), .ZN(n611) );
  XNOR2_X2 U503 ( .A(n496), .B(n448), .ZN(n769) );
  XNOR2_X2 U504 ( .A(n522), .B(KEYINPUT4), .ZN(n496) );
  XNOR2_X2 U505 ( .A(n400), .B(KEYINPUT35), .ZN(n781) );
  NAND2_X1 U506 ( .A1(n401), .A2(n601), .ZN(n400) );
  XNOR2_X1 U507 ( .A(n402), .B(KEYINPUT34), .ZN(n401) );
  XNOR2_X1 U508 ( .A(n405), .B(n404), .ZN(n403) );
  XNOR2_X1 U509 ( .A(n435), .B(n436), .ZN(n404) );
  NAND2_X1 U510 ( .A1(n517), .A2(G221), .ZN(n405) );
  AND2_X1 U511 ( .A1(n406), .A2(n536), .ZN(n557) );
  INV_X1 U512 ( .A(n700), .ZN(n406) );
  NAND2_X1 U513 ( .A1(n409), .A2(n407), .ZN(n411) );
  NAND2_X1 U514 ( .A1(n566), .A2(KEYINPUT89), .ZN(n408) );
  NAND2_X1 U515 ( .A1(n571), .A2(n566), .ZN(n409) );
  NAND2_X1 U516 ( .A1(n567), .A2(n411), .ZN(n410) );
  XNOR2_X2 U517 ( .A(n413), .B(G116), .ZN(n518) );
  XNOR2_X2 U518 ( .A(n416), .B(G110), .ZN(n487) );
  NAND2_X1 U519 ( .A1(n616), .A2(n781), .ZN(n418) );
  NAND2_X1 U520 ( .A1(n633), .A2(n634), .ZN(n419) );
  NAND2_X1 U521 ( .A1(n420), .A2(n741), .ZN(n628) );
  NAND2_X1 U522 ( .A1(n689), .A2(n703), .ZN(n420) );
  XNOR2_X1 U523 ( .A(n632), .B(n631), .ZN(n639) );
  XOR2_X1 U524 ( .A(n441), .B(n440), .Z(n423) );
  XNOR2_X1 U525 ( .A(n465), .B(n464), .ZN(n469) );
  XNOR2_X1 U526 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(n473) );
  BUF_X1 U528 ( .A(n642), .Z(n770) );
  INV_X1 U529 ( .A(n513), .ZN(n429) );
  INV_X1 U530 ( .A(n454), .ZN(n428) );
  XNOR2_X1 U531 ( .A(n429), .B(n428), .ZN(n768) );
  XNOR2_X2 U532 ( .A(n430), .B(G953), .ZN(n771) );
  NAND2_X1 U533 ( .A1(n771), .A2(G234), .ZN(n434) );
  XNOR2_X1 U534 ( .A(KEYINPUT70), .B(KEYINPUT90), .ZN(n432) );
  XNOR2_X1 U535 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n431) );
  XNOR2_X1 U536 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U537 ( .A(n434), .B(n433), .ZN(n517) );
  XNOR2_X1 U538 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n436) );
  XNOR2_X1 U539 ( .A(G128), .B(n487), .ZN(n435) );
  NAND2_X1 U540 ( .A1(n635), .A2(G234), .ZN(n437) );
  XNOR2_X1 U541 ( .A(n437), .B(KEYINPUT20), .ZN(n443) );
  NAND2_X1 U542 ( .A1(n443), .A2(G217), .ZN(n441) );
  XNOR2_X1 U543 ( .A(KEYINPUT85), .B(KEYINPUT99), .ZN(n439) );
  XNOR2_X1 U544 ( .A(KEYINPUT25), .B(KEYINPUT84), .ZN(n438) );
  XNOR2_X1 U545 ( .A(n439), .B(n438), .ZN(n440) );
  INV_X1 U546 ( .A(n609), .ZN(n607) );
  INV_X1 U547 ( .A(n443), .ZN(n445) );
  INV_X1 U548 ( .A(G221), .ZN(n444) );
  OR2_X1 U549 ( .A1(n445), .A2(n444), .ZN(n447) );
  INV_X1 U550 ( .A(KEYINPUT21), .ZN(n446) );
  XNOR2_X1 U551 ( .A(n447), .B(n446), .ZN(n720) );
  XNOR2_X2 U552 ( .A(G143), .B(G128), .ZN(n522) );
  XNOR2_X1 U553 ( .A(n530), .B(G131), .ZN(n448) );
  NAND2_X1 U554 ( .A1(n771), .A2(G227), .ZN(n452) );
  XNOR2_X1 U555 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U556 ( .A(n452), .B(n451), .ZN(n456) );
  XNOR2_X1 U557 ( .A(KEYINPUT78), .B(KEYINPUT98), .ZN(n453) );
  XNOR2_X1 U558 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U559 ( .A(n456), .B(n455), .ZN(n457) );
  OR2_X2 U560 ( .A1(n680), .A2(G902), .ZN(n461) );
  XNOR2_X1 U561 ( .A(KEYINPUT75), .B(G469), .ZN(n459) );
  INV_X1 U562 ( .A(KEYINPUT74), .ZN(n458) );
  XNOR2_X1 U563 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X2 U564 ( .A(n461), .B(n460), .ZN(n560) );
  NAND2_X1 U565 ( .A1(n617), .A2(n560), .ZN(n463) );
  INV_X1 U566 ( .A(KEYINPUT100), .ZN(n462) );
  AND2_X1 U567 ( .A1(n509), .A2(G210), .ZN(n465) );
  XNOR2_X1 U568 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U569 ( .A(G113), .B(G101), .ZN(n470) );
  XNOR2_X1 U570 ( .A(n470), .B(KEYINPUT3), .ZN(n472) );
  XNOR2_X1 U571 ( .A(n472), .B(n471), .ZN(n489) );
  XNOR2_X1 U572 ( .A(n473), .B(n489), .ZN(n474) );
  XNOR2_X1 U573 ( .A(G472), .B(KEYINPUT103), .ZN(n476) );
  INV_X1 U574 ( .A(KEYINPUT79), .ZN(n475) );
  XNOR2_X1 U575 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X2 U576 ( .A(n478), .B(n477), .ZN(n556) );
  XNOR2_X1 U577 ( .A(n479), .B(KEYINPUT81), .ZN(n499) );
  NAND2_X1 U578 ( .A1(n499), .A2(G214), .ZN(n735) );
  XNOR2_X1 U579 ( .A(n480), .B(KEYINPUT30), .ZN(n485) );
  NAND2_X1 U580 ( .A1(G952), .A2(n756), .ZN(n591) );
  INV_X1 U581 ( .A(n771), .ZN(n651) );
  NOR2_X1 U582 ( .A1(n514), .A2(G900), .ZN(n481) );
  NAND2_X1 U583 ( .A1(n651), .A2(n481), .ZN(n482) );
  NAND2_X1 U584 ( .A1(n591), .A2(n482), .ZN(n484) );
  XNOR2_X1 U585 ( .A(n483), .B(KEYINPUT14), .ZN(n750) );
  AND2_X1 U586 ( .A1(n484), .A2(n750), .ZN(n533) );
  AND2_X1 U587 ( .A1(n485), .A2(n533), .ZN(n486) );
  NAND2_X1 U588 ( .A1(n771), .A2(G224), .ZN(n491) );
  XNOR2_X1 U589 ( .A(n492), .B(n491), .ZN(n498) );
  XOR2_X1 U590 ( .A(G146), .B(G125), .Z(n494) );
  XOR2_X1 U591 ( .A(KEYINPUT18), .B(KEYINPUT86), .Z(n493) );
  XNOR2_X1 U592 ( .A(n494), .B(n493), .ZN(n495) );
  AND2_X1 U593 ( .A1(n499), .A2(G210), .ZN(n500) );
  BUF_X1 U594 ( .A(n558), .Z(n549) );
  INV_X1 U595 ( .A(KEYINPUT38), .ZN(n501) );
  XNOR2_X1 U596 ( .A(n549), .B(n501), .ZN(n736) );
  NAND2_X1 U597 ( .A1(n553), .A2(n736), .ZN(n502) );
  XNOR2_X1 U598 ( .A(n504), .B(n355), .ZN(n508) );
  XNOR2_X1 U599 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U600 ( .A(n508), .B(n507), .Z(n511) );
  NAND2_X1 U601 ( .A1(G214), .A2(n509), .ZN(n510) );
  XNOR2_X1 U602 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U603 ( .A(n513), .B(n512), .ZN(n655) );
  NAND2_X1 U604 ( .A1(n655), .A2(n514), .ZN(n516) );
  XNOR2_X1 U605 ( .A(KEYINPUT13), .B(G475), .ZN(n515) );
  XNOR2_X1 U606 ( .A(n516), .B(n515), .ZN(n551) );
  INV_X1 U607 ( .A(n551), .ZN(n528) );
  NAND2_X1 U608 ( .A1(n517), .A2(G217), .ZN(n526) );
  XNOR2_X1 U609 ( .A(n519), .B(KEYINPUT105), .ZN(n520) );
  XNOR2_X1 U610 ( .A(n518), .B(n520), .ZN(n524) );
  XNOR2_X1 U611 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n521) );
  XNOR2_X1 U612 ( .A(n357), .B(n521), .ZN(n523) );
  XNOR2_X1 U613 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U614 ( .A(n526), .B(n525), .ZN(n673) );
  OR2_X1 U615 ( .A1(n673), .A2(G902), .ZN(n527) );
  XNOR2_X1 U616 ( .A(n527), .B(G478), .ZN(n544) );
  INV_X1 U617 ( .A(n544), .ZN(n550) );
  OR2_X1 U618 ( .A1(n528), .A2(n550), .ZN(n702) );
  INV_X1 U619 ( .A(n702), .ZN(n694) );
  AND2_X1 U620 ( .A1(n529), .A2(n694), .ZN(n588) );
  XNOR2_X1 U621 ( .A(n588), .B(n530), .ZN(G36) );
  XOR2_X1 U622 ( .A(G137), .B(KEYINPUT126), .Z(n543) );
  AND2_X1 U623 ( .A1(n736), .A2(n735), .ZN(n742) );
  AND2_X1 U624 ( .A1(n551), .A2(n550), .ZN(n738) );
  NAND2_X1 U625 ( .A1(n742), .A2(n738), .ZN(n532) );
  INV_X1 U626 ( .A(KEYINPUT41), .ZN(n531) );
  XNOR2_X1 U627 ( .A(n532), .B(n531), .ZN(n732) );
  AND2_X1 U628 ( .A1(n720), .A2(n533), .ZN(n534) );
  NAND2_X1 U629 ( .A1(n609), .A2(n534), .ZN(n535) );
  NAND2_X1 U630 ( .A1(n536), .A2(n727), .ZN(n539) );
  INV_X1 U631 ( .A(KEYINPUT112), .ZN(n537) );
  XNOR2_X1 U632 ( .A(n537), .B(KEYINPUT28), .ZN(n538) );
  XNOR2_X1 U633 ( .A(n539), .B(n538), .ZN(n540) );
  AND2_X1 U634 ( .A1(n560), .A2(n540), .ZN(n564) );
  INV_X1 U635 ( .A(n564), .ZN(n541) );
  XNOR2_X1 U636 ( .A(n542), .B(KEYINPUT42), .ZN(n545) );
  XOR2_X1 U637 ( .A(n543), .B(n545), .Z(G39) );
  NAND2_X1 U638 ( .A1(n668), .A2(n545), .ZN(n548) );
  XNOR2_X1 U639 ( .A(KEYINPUT65), .B(KEYINPUT94), .ZN(n546) );
  XNOR2_X1 U640 ( .A(n546), .B(KEYINPUT46), .ZN(n547) );
  XNOR2_X1 U641 ( .A(n548), .B(n547), .ZN(n577) );
  INV_X1 U642 ( .A(KEYINPUT88), .ZN(n568) );
  INV_X1 U643 ( .A(n549), .ZN(n584) );
  OR2_X1 U644 ( .A1(n551), .A2(n550), .ZN(n600) );
  NOR2_X1 U645 ( .A1(n584), .A2(n600), .ZN(n552) );
  NAND2_X1 U646 ( .A1(n700), .A2(n702), .ZN(n741) );
  INV_X1 U647 ( .A(n741), .ZN(n565) );
  NOR2_X1 U648 ( .A1(n565), .A2(KEYINPUT88), .ZN(n554) );
  NOR2_X1 U649 ( .A1(n555), .A2(n554), .ZN(n562) );
  NAND2_X1 U650 ( .A1(n557), .A2(n626), .ZN(n581) );
  NOR2_X1 U651 ( .A1(n581), .A2(n563), .ZN(n559) );
  XNOR2_X1 U652 ( .A(KEYINPUT36), .B(n559), .ZN(n561) );
  NAND2_X1 U653 ( .A1(n561), .A2(n598), .ZN(n705) );
  AND2_X1 U654 ( .A1(n562), .A2(n705), .ZN(n567) );
  AND2_X1 U655 ( .A1(n596), .A2(n564), .ZN(n571) );
  NAND2_X1 U656 ( .A1(KEYINPUT88), .A2(n565), .ZN(n566) );
  OR2_X1 U657 ( .A1(KEYINPUT89), .A2(n569), .ZN(n570) );
  INV_X1 U658 ( .A(KEYINPUT47), .ZN(n572) );
  AND2_X1 U659 ( .A1(n741), .A2(n572), .ZN(n573) );
  NAND2_X1 U660 ( .A1(n571), .A2(n573), .ZN(n574) );
  XNOR2_X1 U661 ( .A(n574), .B(KEYINPUT80), .ZN(n575) );
  NAND2_X1 U662 ( .A1(n577), .A2(n576), .ZN(n580) );
  XNOR2_X1 U663 ( .A(KEYINPUT93), .B(KEYINPUT48), .ZN(n578) );
  XNOR2_X1 U664 ( .A(n578), .B(KEYINPUT72), .ZN(n579) );
  XNOR2_X1 U665 ( .A(n580), .B(n579), .ZN(n590) );
  NOR2_X1 U666 ( .A1(n581), .A2(n598), .ZN(n582) );
  NAND2_X1 U667 ( .A1(n582), .A2(n735), .ZN(n583) );
  XNOR2_X1 U668 ( .A(n583), .B(KEYINPUT43), .ZN(n585) );
  AND2_X1 U669 ( .A1(n585), .A2(n584), .ZN(n587) );
  INV_X1 U670 ( .A(KEYINPUT111), .ZN(n586) );
  XNOR2_X1 U671 ( .A(n587), .B(n586), .ZN(n780) );
  NOR2_X1 U672 ( .A1(n780), .A2(n588), .ZN(n589) );
  NAND2_X1 U673 ( .A1(n590), .A2(n589), .ZN(n642) );
  XNOR2_X1 U674 ( .A(n642), .B(KEYINPUT83), .ZN(n634) );
  XOR2_X1 U675 ( .A(KEYINPUT97), .B(G898), .Z(n759) );
  NOR2_X1 U676 ( .A1(n759), .A2(n756), .ZN(n765) );
  NAND2_X1 U677 ( .A1(n765), .A2(G902), .ZN(n592) );
  AND2_X1 U678 ( .A1(n592), .A2(n591), .ZN(n594) );
  INV_X1 U679 ( .A(n750), .ZN(n593) );
  NOR2_X1 U680 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U681 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U682 ( .A(KEYINPUT110), .B(KEYINPUT33), .Z(n599) );
  XNOR2_X1 U683 ( .A(n600), .B(KEYINPUT87), .ZN(n601) );
  NAND2_X1 U684 ( .A1(n738), .A2(n720), .ZN(n602) );
  INV_X1 U685 ( .A(KEYINPUT22), .ZN(n604) );
  INV_X1 U686 ( .A(KEYINPUT109), .ZN(n606) );
  NOR2_X1 U687 ( .A1(n607), .A2(n727), .ZN(n608) );
  XNOR2_X1 U688 ( .A(n609), .B(KEYINPUT106), .ZN(n722) );
  NAND2_X1 U689 ( .A1(n722), .A2(n598), .ZN(n610) );
  XOR2_X1 U690 ( .A(KEYINPUT108), .B(n610), .Z(n612) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n614) );
  INV_X1 U692 ( .A(KEYINPUT44), .ZN(n615) );
  XOR2_X1 U693 ( .A(KEYINPUT104), .B(KEYINPUT31), .Z(n619) );
  INV_X1 U694 ( .A(n617), .ZN(n717) );
  NOR2_X1 U695 ( .A1(n717), .A2(n556), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n618), .A2(n598), .ZN(n729) );
  INV_X1 U697 ( .A(n620), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n623), .B(KEYINPUT101), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n624), .A2(n556), .ZN(n689) );
  NOR2_X1 U701 ( .A1(n626), .A2(n722), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n625), .A2(n627), .ZN(n687) );
  NAND2_X1 U703 ( .A1(n628), .A2(n687), .ZN(n629) );
  XNOR2_X1 U704 ( .A(KEYINPUT107), .B(n629), .ZN(n630) );
  INV_X1 U705 ( .A(KEYINPUT45), .ZN(n631) );
  NOR2_X1 U706 ( .A1(n639), .A2(n635), .ZN(n633) );
  INV_X1 U707 ( .A(n635), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n636), .A2(KEYINPUT2), .ZN(n637) );
  INV_X1 U709 ( .A(KEYINPUT67), .ZN(n638) );
  INV_X1 U710 ( .A(n640), .ZN(n641) );
  NAND2_X1 U711 ( .A1(n641), .A2(KEYINPUT2), .ZN(n643) );
  INV_X1 U712 ( .A(KEYINPUT66), .ZN(n645) );
  NAND2_X1 U713 ( .A1(n677), .A2(G472), .ZN(n649) );
  INV_X1 U714 ( .A(n646), .ZN(n647) );
  XNOR2_X1 U715 ( .A(n647), .B(KEYINPUT62), .ZN(n648) );
  XNOR2_X1 U716 ( .A(n649), .B(n648), .ZN(n652) );
  INV_X1 U717 ( .A(G952), .ZN(n650) );
  NAND2_X1 U718 ( .A1(n651), .A2(n650), .ZN(n671) );
  NAND2_X1 U719 ( .A1(n652), .A2(n671), .ZN(n653) );
  XNOR2_X1 U720 ( .A(n653), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U721 ( .A1(n677), .A2(G475), .ZN(n657) );
  XOR2_X1 U722 ( .A(KEYINPUT96), .B(KEYINPUT59), .Z(n654) );
  XNOR2_X1 U723 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U724 ( .A(n657), .B(n656), .ZN(n658) );
  NAND2_X1 U725 ( .A1(n658), .A2(n671), .ZN(n660) );
  XOR2_X1 U726 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n659) );
  XNOR2_X1 U727 ( .A(n660), .B(n659), .ZN(G60) );
  NAND2_X1 U728 ( .A1(n677), .A2(G210), .ZN(n664) );
  XOR2_X1 U729 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n662) );
  XNOR2_X1 U730 ( .A(n661), .B(n662), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n665), .A2(n671), .ZN(n667) );
  INV_X1 U733 ( .A(KEYINPUT56), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n667), .B(n666), .ZN(G51) );
  XNOR2_X1 U735 ( .A(n668), .B(G131), .ZN(G33) );
  NAND2_X1 U736 ( .A1(n677), .A2(G217), .ZN(n670) );
  XNOR2_X1 U737 ( .A(n670), .B(n669), .ZN(n672) );
  INV_X1 U738 ( .A(n671), .ZN(n684) );
  NOR2_X1 U739 ( .A1(n672), .A2(n684), .ZN(G66) );
  NAND2_X1 U740 ( .A1(n677), .A2(G478), .ZN(n675) );
  XNOR2_X1 U741 ( .A(n673), .B(KEYINPUT122), .ZN(n674) );
  XNOR2_X1 U742 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X1 U743 ( .A1(n676), .A2(n684), .ZN(G63) );
  NAND2_X1 U744 ( .A1(n677), .A2(G469), .ZN(n683) );
  XOR2_X1 U745 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n679) );
  XNOR2_X1 U746 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n679), .B(n678), .ZN(n681) );
  XOR2_X1 U748 ( .A(n681), .B(n680), .Z(n682) );
  XNOR2_X1 U749 ( .A(n683), .B(n682), .ZN(n685) );
  NOR2_X1 U750 ( .A1(n685), .A2(n684), .ZN(G54) );
  XOR2_X1 U751 ( .A(G101), .B(KEYINPUT113), .Z(n686) );
  XNOR2_X1 U752 ( .A(n687), .B(n686), .ZN(G3) );
  NOR2_X1 U753 ( .A1(n689), .A2(n700), .ZN(n688) );
  XOR2_X1 U754 ( .A(G104), .B(n688), .Z(G6) );
  NOR2_X1 U755 ( .A1(n689), .A2(n702), .ZN(n691) );
  XNOR2_X1 U756 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n690) );
  XNOR2_X1 U757 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U758 ( .A(G107), .B(n692), .ZN(G9) );
  XOR2_X1 U759 ( .A(G110), .B(n693), .Z(G12) );
  XOR2_X1 U760 ( .A(G128), .B(KEYINPUT29), .Z(n696) );
  NAND2_X1 U761 ( .A1(n571), .A2(n694), .ZN(n695) );
  XNOR2_X1 U762 ( .A(n696), .B(n695), .ZN(G30) );
  XNOR2_X1 U763 ( .A(G143), .B(KEYINPUT114), .ZN(n697) );
  INV_X1 U764 ( .A(n571), .ZN(n698) );
  NOR2_X1 U765 ( .A1(n698), .A2(n700), .ZN(n699) );
  XOR2_X1 U766 ( .A(G146), .B(n699), .Z(G48) );
  NOR2_X1 U767 ( .A1(n703), .A2(n700), .ZN(n701) );
  XOR2_X1 U768 ( .A(G113), .B(n701), .Z(G15) );
  NOR2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U770 ( .A(G116), .B(n704), .Z(G18) );
  XNOR2_X1 U771 ( .A(KEYINPUT37), .B(KEYINPUT115), .ZN(n706) );
  XNOR2_X1 U772 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U773 ( .A(G125), .B(n707), .ZN(G27) );
  NOR2_X1 U774 ( .A1(n356), .A2(n770), .ZN(n708) );
  NOR2_X1 U775 ( .A1(n708), .A2(KEYINPUT91), .ZN(n709) );
  XNOR2_X1 U776 ( .A(n709), .B(KEYINPUT2), .ZN(n713) );
  INV_X1 U777 ( .A(n770), .ZN(n710) );
  NAND2_X1 U778 ( .A1(n356), .A2(n710), .ZN(n711) );
  NAND2_X1 U779 ( .A1(n711), .A2(KEYINPUT91), .ZN(n712) );
  NAND2_X1 U780 ( .A1(n713), .A2(n712), .ZN(n716) );
  NOR2_X1 U781 ( .A1(n746), .A2(n732), .ZN(n714) );
  XNOR2_X1 U782 ( .A(n714), .B(KEYINPUT119), .ZN(n715) );
  NAND2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n754) );
  INV_X1 U784 ( .A(n598), .ZN(n718) );
  NAND2_X1 U785 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U786 ( .A(KEYINPUT50), .B(n719), .ZN(n726) );
  XOR2_X1 U787 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n724) );
  INV_X1 U788 ( .A(n720), .ZN(n721) );
  NAND2_X1 U789 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U790 ( .A(n724), .B(n723), .ZN(n725) );
  NAND2_X1 U791 ( .A1(n726), .A2(n725), .ZN(n728) );
  OR2_X1 U792 ( .A1(n728), .A2(n727), .ZN(n730) );
  NAND2_X1 U793 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U794 ( .A(n731), .B(KEYINPUT51), .ZN(n733) );
  NOR2_X1 U795 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U796 ( .A(KEYINPUT117), .B(n734), .Z(n748) );
  NOR2_X1 U797 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U798 ( .A(n737), .B(KEYINPUT118), .ZN(n740) );
  INV_X1 U799 ( .A(n738), .ZN(n739) );
  NOR2_X1 U800 ( .A1(n740), .A2(n739), .ZN(n744) );
  AND2_X1 U801 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U802 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U803 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U804 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U805 ( .A(KEYINPUT52), .B(n749), .ZN(n752) );
  NAND2_X1 U806 ( .A1(n750), .A2(G952), .ZN(n751) );
  NOR2_X1 U807 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U808 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U809 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U810 ( .A(KEYINPUT53), .B(n757), .Z(G75) );
  NAND2_X1 U811 ( .A1(G953), .A2(G224), .ZN(n758) );
  XNOR2_X1 U812 ( .A(KEYINPUT61), .B(n758), .ZN(n760) );
  NAND2_X1 U813 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U814 ( .A(n761), .B(KEYINPUT123), .ZN(n763) );
  NOR2_X1 U815 ( .A1(n356), .A2(G953), .ZN(n762) );
  NOR2_X1 U816 ( .A1(n763), .A2(n762), .ZN(n767) );
  NOR2_X1 U817 ( .A1(n764), .A2(n765), .ZN(n766) );
  XOR2_X1 U818 ( .A(n767), .B(n766), .Z(G69) );
  XOR2_X1 U819 ( .A(n769), .B(n768), .Z(n774) );
  XNOR2_X1 U820 ( .A(n770), .B(n774), .ZN(n772) );
  NAND2_X1 U821 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U822 ( .A(n773), .B(KEYINPUT124), .ZN(n778) );
  XNOR2_X1 U823 ( .A(n774), .B(G227), .ZN(n775) );
  NAND2_X1 U824 ( .A1(n775), .A2(G900), .ZN(n776) );
  NAND2_X1 U825 ( .A1(n776), .A2(G953), .ZN(n777) );
  NAND2_X1 U826 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U827 ( .A(KEYINPUT125), .B(n779), .Z(G72) );
  XOR2_X1 U828 ( .A(G140), .B(n780), .Z(G42) );
  XOR2_X1 U829 ( .A(n781), .B(G122), .Z(G24) );
  XOR2_X1 U830 ( .A(G119), .B(n782), .Z(G21) );
endmodule

