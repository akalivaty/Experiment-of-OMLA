

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U552 ( .A1(n522), .A2(G2104), .ZN(n884) );
  NOR2_X1 U553 ( .A1(n561), .A2(n560), .ZN(G164) );
  NOR2_X2 U554 ( .A1(n690), .A2(n950), .ZN(n692) );
  BUF_X1 U555 ( .A(n565), .Z(n536) );
  NOR2_X2 U556 ( .A1(G2104), .A2(n522), .ZN(n887) );
  NOR2_X2 U557 ( .A1(n777), .A2(n778), .ZN(n710) );
  XNOR2_X1 U558 ( .A(n756), .B(n755), .ZN(n757) );
  NOR2_X2 U559 ( .A1(n530), .A2(n529), .ZN(G160) );
  AND2_X1 U560 ( .A1(n823), .A2(n971), .ZN(n518) );
  NOR2_X1 U561 ( .A1(n723), .A2(n844), .ZN(n687) );
  XNOR2_X1 U562 ( .A(KEYINPUT32), .B(KEYINPUT100), .ZN(n735) );
  INV_X1 U563 ( .A(KEYINPUT64), .ZN(n755) );
  XNOR2_X1 U564 ( .A(n736), .B(n735), .ZN(n763) );
  INV_X1 U565 ( .A(KEYINPUT13), .ZN(n545) );
  OR2_X1 U566 ( .A1(n808), .A2(n518), .ZN(n809) );
  NOR2_X1 U567 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U568 ( .A1(G651), .A2(n653), .ZN(n647) );
  INV_X1 U569 ( .A(KEYINPUT75), .ZN(n554) );
  XNOR2_X1 U570 ( .A(n555), .B(n554), .ZN(n950) );
  INV_X1 U571 ( .A(G2105), .ZN(n522) );
  NAND2_X1 U572 ( .A1(G101), .A2(n884), .ZN(n521) );
  XNOR2_X1 U573 ( .A(KEYINPUT23), .B(KEYINPUT69), .ZN(n519) );
  XNOR2_X1 U574 ( .A(n519), .B(KEYINPUT68), .ZN(n520) );
  XNOR2_X1 U575 ( .A(n521), .B(n520), .ZN(n525) );
  NAND2_X1 U576 ( .A1(G125), .A2(n887), .ZN(n523) );
  XOR2_X1 U577 ( .A(KEYINPUT67), .B(n523), .Z(n524) );
  NAND2_X1 U578 ( .A1(n525), .A2(n524), .ZN(n530) );
  NOR2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XOR2_X1 U580 ( .A(KEYINPUT17), .B(n526), .Z(n607) );
  NAND2_X1 U581 ( .A1(G137), .A2(n607), .ZN(n528) );
  AND2_X1 U582 ( .A1(G2104), .A2(G2105), .ZN(n889) );
  NAND2_X1 U583 ( .A1(G113), .A2(n889), .ZN(n527) );
  NAND2_X1 U584 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U585 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .Z(n653) );
  NAND2_X1 U587 ( .A1(G52), .A2(n647), .ZN(n533) );
  NOR2_X1 U588 ( .A1(G543), .A2(n534), .ZN(n531) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n531), .Z(n547) );
  BUF_X1 U590 ( .A(n547), .Z(n651) );
  NAND2_X1 U591 ( .A1(G64), .A2(n651), .ZN(n532) );
  NAND2_X1 U592 ( .A1(n533), .A2(n532), .ZN(n541) );
  INV_X1 U593 ( .A(G651), .ZN(n534) );
  NOR2_X2 U594 ( .A1(n653), .A2(n534), .ZN(n637) );
  NAND2_X1 U595 ( .A1(n637), .A2(G77), .ZN(n538) );
  NOR2_X1 U596 ( .A1(G651), .A2(G543), .ZN(n535) );
  XNOR2_X1 U597 ( .A(n535), .B(KEYINPUT66), .ZN(n565) );
  NAND2_X1 U598 ( .A1(G90), .A2(n536), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n539), .Z(n540) );
  NOR2_X1 U601 ( .A1(n541), .A2(n540), .ZN(G171) );
  NAND2_X1 U602 ( .A1(G81), .A2(n565), .ZN(n542) );
  XNOR2_X1 U603 ( .A(n542), .B(KEYINPUT12), .ZN(n544) );
  NAND2_X1 U604 ( .A1(G68), .A2(n637), .ZN(n543) );
  NAND2_X1 U605 ( .A1(n544), .A2(n543), .ZN(n546) );
  XNOR2_X1 U606 ( .A(n546), .B(n545), .ZN(n550) );
  NAND2_X1 U607 ( .A1(n547), .A2(G56), .ZN(n548) );
  XOR2_X1 U608 ( .A(KEYINPUT14), .B(n548), .Z(n549) );
  XNOR2_X1 U609 ( .A(n551), .B(KEYINPUT74), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G43), .A2(n647), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n555) );
  INV_X1 U612 ( .A(G860), .ZN(n596) );
  OR2_X1 U613 ( .A1(n950), .A2(n596), .ZN(G153) );
  INV_X1 U614 ( .A(G132), .ZN(G219) );
  INV_X1 U615 ( .A(G82), .ZN(G220) );
  INV_X1 U616 ( .A(G57), .ZN(G237) );
  AND2_X1 U617 ( .A1(n607), .A2(G138), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G126), .A2(n887), .ZN(n557) );
  NAND2_X1 U619 ( .A1(G114), .A2(n889), .ZN(n556) );
  AND2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G102), .A2(n884), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U623 ( .A1(G51), .A2(n647), .ZN(n563) );
  NAND2_X1 U624 ( .A1(G63), .A2(n651), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U626 ( .A(KEYINPUT6), .B(n564), .ZN(n572) );
  NAND2_X1 U627 ( .A1(G89), .A2(n565), .ZN(n566) );
  XNOR2_X1 U628 ( .A(n566), .B(KEYINPUT4), .ZN(n568) );
  NAND2_X1 U629 ( .A1(G76), .A2(n637), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U631 ( .A(KEYINPUT5), .B(n569), .Z(n570) );
  XNOR2_X1 U632 ( .A(KEYINPUT78), .B(n570), .ZN(n571) );
  NOR2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n574) );
  XNOR2_X1 U634 ( .A(KEYINPUT79), .B(KEYINPUT7), .ZN(n573) );
  XNOR2_X1 U635 ( .A(n574), .B(n573), .ZN(G168) );
  XOR2_X1 U636 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U637 ( .A1(G94), .A2(G452), .ZN(n575) );
  XOR2_X1 U638 ( .A(KEYINPUT72), .B(n575), .Z(G173) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U640 ( .A(n576), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U641 ( .A(G223), .B(KEYINPUT73), .ZN(n828) );
  NAND2_X1 U642 ( .A1(n828), .A2(G567), .ZN(n577) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(n577), .Z(G234) );
  XOR2_X1 U644 ( .A(KEYINPUT76), .B(G171), .Z(G301) );
  NAND2_X1 U645 ( .A1(G868), .A2(G301), .ZN(n587) );
  NAND2_X1 U646 ( .A1(G54), .A2(n647), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n637), .A2(G79), .ZN(n579) );
  NAND2_X1 U648 ( .A1(G92), .A2(n536), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U650 ( .A1(G66), .A2(n651), .ZN(n580) );
  XNOR2_X1 U651 ( .A(KEYINPUT77), .B(n580), .ZN(n581) );
  NOR2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U653 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U654 ( .A(n585), .B(KEYINPUT15), .ZN(n969) );
  OR2_X1 U655 ( .A1(n969), .A2(G868), .ZN(n586) );
  NAND2_X1 U656 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U657 ( .A1(G53), .A2(n647), .ZN(n589) );
  NAND2_X1 U658 ( .A1(G65), .A2(n651), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U660 ( .A1(n637), .A2(G78), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G91), .A2(n536), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U663 ( .A1(n593), .A2(n592), .ZN(n951) );
  INV_X1 U664 ( .A(n951), .ZN(G299) );
  NOR2_X1 U665 ( .A1(G868), .A2(G299), .ZN(n595) );
  INV_X1 U666 ( .A(G868), .ZN(n665) );
  NOR2_X1 U667 ( .A1(G286), .A2(n665), .ZN(n594) );
  NOR2_X1 U668 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U669 ( .A1(n596), .A2(G559), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n597), .A2(n969), .ZN(n598) );
  XNOR2_X1 U671 ( .A(n598), .B(KEYINPUT80), .ZN(n599) );
  XNOR2_X1 U672 ( .A(KEYINPUT16), .B(n599), .ZN(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n950), .ZN(n600) );
  XOR2_X1 U674 ( .A(KEYINPUT81), .B(n600), .Z(n603) );
  NAND2_X1 U675 ( .A1(G868), .A2(n969), .ZN(n601) );
  NOR2_X1 U676 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n603), .A2(n602), .ZN(G282) );
  XOR2_X1 U678 ( .A(G2100), .B(KEYINPUT82), .Z(n613) );
  NAND2_X1 U679 ( .A1(n887), .A2(G123), .ZN(n604) );
  XNOR2_X1 U680 ( .A(n604), .B(KEYINPUT18), .ZN(n606) );
  NAND2_X1 U681 ( .A1(G111), .A2(n889), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n611) );
  BUF_X1 U683 ( .A(n607), .Z(n883) );
  NAND2_X1 U684 ( .A1(G135), .A2(n883), .ZN(n609) );
  NAND2_X1 U685 ( .A1(G99), .A2(n884), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n928) );
  XNOR2_X1 U688 ( .A(G2096), .B(n928), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(G156) );
  NAND2_X1 U690 ( .A1(n637), .A2(G80), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G93), .A2(n536), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U693 ( .A1(G55), .A2(n647), .ZN(n617) );
  NAND2_X1 U694 ( .A1(G67), .A2(n651), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n618) );
  OR2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n664) );
  NAND2_X1 U697 ( .A1(G559), .A2(n969), .ZN(n620) );
  XOR2_X1 U698 ( .A(n950), .B(n620), .Z(n662) );
  XNOR2_X1 U699 ( .A(KEYINPUT83), .B(n662), .ZN(n621) );
  NOR2_X1 U700 ( .A1(G860), .A2(n621), .ZN(n622) );
  XOR2_X1 U701 ( .A(n664), .B(n622), .Z(G145) );
  NAND2_X1 U702 ( .A1(n637), .A2(G75), .ZN(n624) );
  NAND2_X1 U703 ( .A1(G88), .A2(n536), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G50), .A2(n647), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G62), .A2(n651), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U708 ( .A1(n628), .A2(n627), .ZN(G166) );
  INV_X1 U709 ( .A(G166), .ZN(G303) );
  NAND2_X1 U710 ( .A1(n637), .A2(G72), .ZN(n630) );
  NAND2_X1 U711 ( .A1(G85), .A2(n536), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U713 ( .A(KEYINPUT70), .B(n631), .ZN(n634) );
  NAND2_X1 U714 ( .A1(G47), .A2(n647), .ZN(n632) );
  XNOR2_X1 U715 ( .A(KEYINPUT71), .B(n632), .ZN(n633) );
  NOR2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n651), .A2(G60), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(G290) );
  NAND2_X1 U719 ( .A1(n637), .A2(G73), .ZN(n638) );
  XNOR2_X1 U720 ( .A(KEYINPUT2), .B(n638), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n651), .A2(G61), .ZN(n640) );
  NAND2_X1 U722 ( .A1(G86), .A2(n536), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U724 ( .A(KEYINPUT86), .B(n641), .Z(n642) );
  NAND2_X1 U725 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U726 ( .A(n644), .B(KEYINPUT87), .ZN(n646) );
  NAND2_X1 U727 ( .A1(G48), .A2(n647), .ZN(n645) );
  NAND2_X1 U728 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U729 ( .A1(G49), .A2(n647), .ZN(n649) );
  NAND2_X1 U730 ( .A1(G74), .A2(G651), .ZN(n648) );
  NAND2_X1 U731 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U732 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U733 ( .A(KEYINPUT84), .B(n652), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n653), .A2(G87), .ZN(n654) );
  XOR2_X1 U735 ( .A(KEYINPUT85), .B(n654), .Z(n655) );
  NAND2_X1 U736 ( .A1(n656), .A2(n655), .ZN(G288) );
  XNOR2_X1 U737 ( .A(KEYINPUT19), .B(n664), .ZN(n658) );
  XOR2_X1 U738 ( .A(G303), .B(n951), .Z(n657) );
  XNOR2_X1 U739 ( .A(n658), .B(n657), .ZN(n661) );
  XNOR2_X1 U740 ( .A(G290), .B(G305), .ZN(n659) );
  XNOR2_X1 U741 ( .A(n659), .B(G288), .ZN(n660) );
  XNOR2_X1 U742 ( .A(n661), .B(n660), .ZN(n901) );
  XNOR2_X1 U743 ( .A(n901), .B(n662), .ZN(n663) );
  NAND2_X1 U744 ( .A1(n663), .A2(G868), .ZN(n667) );
  NAND2_X1 U745 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U746 ( .A1(n667), .A2(n666), .ZN(G295) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n669) );
  NAND2_X1 U748 ( .A1(G2084), .A2(G2078), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U752 ( .A1(n672), .A2(G2072), .ZN(G158) );
  NAND2_X1 U753 ( .A1(G108), .A2(G120), .ZN(n673) );
  NOR2_X1 U754 ( .A1(G237), .A2(n673), .ZN(n674) );
  NAND2_X1 U755 ( .A1(G69), .A2(n674), .ZN(n833) );
  NAND2_X1 U756 ( .A1(G567), .A2(n833), .ZN(n675) );
  XNOR2_X1 U757 ( .A(n675), .B(KEYINPUT89), .ZN(n680) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n676) );
  XNOR2_X1 U759 ( .A(KEYINPUT22), .B(n676), .ZN(n677) );
  NAND2_X1 U760 ( .A1(n677), .A2(G96), .ZN(n678) );
  OR2_X1 U761 ( .A1(G218), .A2(n678), .ZN(n834) );
  AND2_X1 U762 ( .A1(G2106), .A2(n834), .ZN(n679) );
  NOR2_X1 U763 ( .A1(n680), .A2(n679), .ZN(G319) );
  NAND2_X1 U764 ( .A1(G483), .A2(G661), .ZN(n682) );
  INV_X1 U765 ( .A(G319), .ZN(n681) );
  NOR2_X1 U766 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U767 ( .A(n683), .B(KEYINPUT90), .ZN(n831) );
  NAND2_X1 U768 ( .A1(G36), .A2(n831), .ZN(G176) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n685) );
  XNOR2_X1 U770 ( .A(n685), .B(KEYINPUT65), .ZN(n777) );
  NAND2_X1 U771 ( .A1(G160), .A2(G40), .ZN(n778) );
  INV_X1 U772 ( .A(n710), .ZN(n723) );
  INV_X1 U773 ( .A(G1996), .ZN(n844) );
  XOR2_X1 U774 ( .A(KEYINPUT26), .B(KEYINPUT98), .Z(n686) );
  XNOR2_X1 U775 ( .A(n687), .B(n686), .ZN(n689) );
  NAND2_X1 U776 ( .A1(n723), .A2(G1341), .ZN(n688) );
  NAND2_X1 U777 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U778 ( .A1(n692), .A2(n969), .ZN(n691) );
  XNOR2_X1 U779 ( .A(n691), .B(KEYINPUT99), .ZN(n698) );
  NAND2_X1 U780 ( .A1(n692), .A2(n969), .ZN(n696) );
  NOR2_X1 U781 ( .A1(n710), .A2(G1348), .ZN(n694) );
  NOR2_X1 U782 ( .A1(G2067), .A2(n723), .ZN(n693) );
  NOR2_X1 U783 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U785 ( .A1(n698), .A2(n697), .ZN(n703) );
  NAND2_X1 U786 ( .A1(n710), .A2(G2072), .ZN(n699) );
  XNOR2_X1 U787 ( .A(n699), .B(KEYINPUT27), .ZN(n701) );
  AND2_X1 U788 ( .A1(G1956), .A2(n723), .ZN(n700) );
  NOR2_X1 U789 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U790 ( .A1(n951), .A2(n704), .ZN(n702) );
  NAND2_X1 U791 ( .A1(n703), .A2(n702), .ZN(n707) );
  NOR2_X1 U792 ( .A1(n951), .A2(n704), .ZN(n705) );
  XOR2_X1 U793 ( .A(n705), .B(KEYINPUT28), .Z(n706) );
  NAND2_X1 U794 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U795 ( .A(n708), .B(KEYINPUT29), .ZN(n739) );
  XNOR2_X1 U796 ( .A(G2078), .B(KEYINPUT25), .ZN(n1004) );
  NAND2_X1 U797 ( .A1(n710), .A2(n1004), .ZN(n709) );
  XOR2_X1 U798 ( .A(KEYINPUT96), .B(n709), .Z(n712) );
  NOR2_X1 U799 ( .A1(n710), .A2(G1961), .ZN(n711) );
  NOR2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U801 ( .A(KEYINPUT97), .B(n713), .ZN(n721) );
  AND2_X1 U802 ( .A1(G171), .A2(n721), .ZN(n738) );
  INV_X1 U803 ( .A(G8), .ZN(n718) );
  NAND2_X1 U804 ( .A1(G8), .A2(n723), .ZN(n774) );
  NOR2_X1 U805 ( .A1(G1971), .A2(n774), .ZN(n715) );
  NOR2_X1 U806 ( .A1(G2090), .A2(n723), .ZN(n714) );
  NOR2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U808 ( .A1(n716), .A2(G303), .ZN(n717) );
  NOR2_X1 U809 ( .A1(n718), .A2(n717), .ZN(n730) );
  OR2_X1 U810 ( .A1(n730), .A2(G286), .ZN(n732) );
  INV_X1 U811 ( .A(n732), .ZN(n719) );
  OR2_X1 U812 ( .A1(n738), .A2(n719), .ZN(n720) );
  NOR2_X1 U813 ( .A1(n739), .A2(n720), .ZN(n734) );
  NOR2_X1 U814 ( .A1(G171), .A2(n721), .ZN(n728) );
  NOR2_X1 U815 ( .A1(n718), .A2(G1966), .ZN(n722) );
  AND2_X1 U816 ( .A1(n723), .A2(n722), .ZN(n743) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n723), .ZN(n737) );
  NOR2_X1 U818 ( .A1(n743), .A2(n737), .ZN(n724) );
  NAND2_X1 U819 ( .A1(G8), .A2(n724), .ZN(n725) );
  XNOR2_X1 U820 ( .A(KEYINPUT30), .B(n725), .ZN(n726) );
  NOR2_X1 U821 ( .A1(G168), .A2(n726), .ZN(n727) );
  NOR2_X1 U822 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U823 ( .A(n729), .B(KEYINPUT31), .ZN(n740) );
  OR2_X1 U824 ( .A1(n740), .A2(n730), .ZN(n731) );
  AND2_X1 U825 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U826 ( .A1(n734), .A2(n733), .ZN(n736) );
  NAND2_X1 U827 ( .A1(n737), .A2(G8), .ZN(n745) );
  NOR2_X1 U828 ( .A1(n739), .A2(n738), .ZN(n741) );
  NOR2_X1 U829 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U831 ( .A1(n745), .A2(n744), .ZN(n764) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n952) );
  INV_X1 U833 ( .A(n774), .ZN(n746) );
  AND2_X1 U834 ( .A1(n952), .A2(n746), .ZN(n748) );
  AND2_X1 U835 ( .A1(n764), .A2(n748), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n763), .A2(n747), .ZN(n754) );
  INV_X1 U837 ( .A(n748), .ZN(n752) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n749) );
  XNOR2_X1 U839 ( .A(KEYINPUT101), .B(n749), .ZN(n750) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n758) );
  INV_X1 U841 ( .A(n758), .ZN(n953) );
  AND2_X1 U842 ( .A1(n750), .A2(n953), .ZN(n751) );
  OR2_X1 U843 ( .A1(n752), .A2(n751), .ZN(n753) );
  AND2_X1 U844 ( .A1(n754), .A2(n753), .ZN(n756) );
  NOR2_X1 U845 ( .A1(KEYINPUT33), .A2(n757), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n758), .A2(KEYINPUT33), .ZN(n759) );
  NOR2_X1 U847 ( .A1(n759), .A2(n774), .ZN(n760) );
  NOR2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n965) );
  NAND2_X1 U850 ( .A1(n762), .A2(n965), .ZN(n770) );
  NAND2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n767) );
  NOR2_X1 U852 ( .A1(G2090), .A2(G303), .ZN(n765) );
  NAND2_X1 U853 ( .A1(G8), .A2(n765), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U855 ( .A1(n768), .A2(n774), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n776) );
  NOR2_X1 U857 ( .A1(G1981), .A2(G305), .ZN(n771) );
  XNOR2_X1 U858 ( .A(n771), .B(KEYINPUT95), .ZN(n772) );
  XNOR2_X1 U859 ( .A(KEYINPUT24), .B(n772), .ZN(n773) );
  NOR2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U861 ( .A1(n776), .A2(n775), .ZN(n810) );
  INV_X1 U862 ( .A(n777), .ZN(n779) );
  NOR2_X1 U863 ( .A1(n779), .A2(n778), .ZN(n823) );
  NAND2_X1 U864 ( .A1(n884), .A2(G104), .ZN(n780) );
  XOR2_X1 U865 ( .A(KEYINPUT91), .B(n780), .Z(n782) );
  NAND2_X1 U866 ( .A1(n883), .A2(G140), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U868 ( .A(KEYINPUT34), .B(n783), .ZN(n789) );
  NAND2_X1 U869 ( .A1(G128), .A2(n887), .ZN(n785) );
  NAND2_X1 U870 ( .A1(G116), .A2(n889), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U872 ( .A(KEYINPUT92), .B(n786), .Z(n787) );
  XNOR2_X1 U873 ( .A(KEYINPUT35), .B(n787), .ZN(n788) );
  NOR2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U875 ( .A(KEYINPUT36), .B(n790), .ZN(n898) );
  XNOR2_X1 U876 ( .A(KEYINPUT37), .B(G2067), .ZN(n820) );
  OR2_X1 U877 ( .A1(n898), .A2(n820), .ZN(n791) );
  XNOR2_X1 U878 ( .A(KEYINPUT93), .B(n791), .ZN(n945) );
  NAND2_X1 U879 ( .A1(n823), .A2(n945), .ZN(n818) );
  NAND2_X1 U880 ( .A1(G131), .A2(n883), .ZN(n793) );
  NAND2_X1 U881 ( .A1(G119), .A2(n887), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n797) );
  NAND2_X1 U883 ( .A1(G95), .A2(n884), .ZN(n795) );
  NAND2_X1 U884 ( .A1(G107), .A2(n889), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n796) );
  OR2_X1 U886 ( .A1(n797), .A2(n796), .ZN(n875) );
  NAND2_X1 U887 ( .A1(G1991), .A2(n875), .ZN(n806) );
  NAND2_X1 U888 ( .A1(G141), .A2(n883), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G129), .A2(n887), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U891 ( .A1(n884), .A2(G105), .ZN(n800) );
  XOR2_X1 U892 ( .A(KEYINPUT38), .B(n800), .Z(n801) );
  NOR2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n804) );
  NAND2_X1 U894 ( .A1(n889), .A2(G117), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n873) );
  NAND2_X1 U896 ( .A1(G1996), .A2(n873), .ZN(n805) );
  NAND2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n933) );
  NAND2_X1 U898 ( .A1(n823), .A2(n933), .ZN(n812) );
  NAND2_X1 U899 ( .A1(n818), .A2(n812), .ZN(n807) );
  XNOR2_X1 U900 ( .A(n807), .B(KEYINPUT94), .ZN(n808) );
  XNOR2_X1 U901 ( .A(G1986), .B(G290), .ZN(n971) );
  OR2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U903 ( .A(n811), .B(KEYINPUT102), .ZN(n825) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n873), .ZN(n925) );
  INV_X1 U905 ( .A(n812), .ZN(n815) );
  NOR2_X1 U906 ( .A1(G1991), .A2(n875), .ZN(n929) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U908 ( .A1(n929), .A2(n813), .ZN(n814) );
  NOR2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U910 ( .A1(n925), .A2(n816), .ZN(n817) );
  XNOR2_X1 U911 ( .A(n817), .B(KEYINPUT39), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U913 ( .A1(n898), .A2(n820), .ZN(n934) );
  NAND2_X1 U914 ( .A1(n821), .A2(n934), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(n827) );
  XOR2_X1 U917 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n826) );
  XNOR2_X1 U918 ( .A(n827), .B(n826), .ZN(G329) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U921 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n830) );
  XOR2_X1 U923 ( .A(KEYINPUT105), .B(n830), .Z(n832) );
  NAND2_X1 U924 ( .A1(n832), .A2(n831), .ZN(G188) );
  XOR2_X1 U925 ( .A(G120), .B(KEYINPUT106), .Z(G236) );
  INV_X1 U927 ( .A(G108), .ZN(G238) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  NOR2_X1 U929 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  XOR2_X1 U931 ( .A(KEYINPUT107), .B(G2084), .Z(n836) );
  XNOR2_X1 U932 ( .A(G2090), .B(G2078), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U934 ( .A(n837), .B(G2096), .Z(n839) );
  XNOR2_X1 U935 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U937 ( .A(G2100), .B(KEYINPUT43), .Z(n841) );
  XNOR2_X1 U938 ( .A(G2678), .B(KEYINPUT42), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U940 ( .A(n843), .B(n842), .Z(G227) );
  XOR2_X1 U941 ( .A(G1976), .B(G1956), .Z(n846) );
  XOR2_X1 U942 ( .A(n844), .B(G1991), .Z(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n856) );
  XOR2_X1 U944 ( .A(G2474), .B(KEYINPUT41), .Z(n848) );
  XNOR2_X1 U945 ( .A(G1986), .B(KEYINPUT109), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U947 ( .A(G1981), .B(G1966), .Z(n850) );
  XNOR2_X1 U948 ( .A(G1971), .B(G1961), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U950 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U951 ( .A(KEYINPUT110), .B(KEYINPUT108), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U954 ( .A1(G112), .A2(n889), .ZN(n863) );
  NAND2_X1 U955 ( .A1(G136), .A2(n883), .ZN(n858) );
  NAND2_X1 U956 ( .A1(G100), .A2(n884), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n861) );
  NAND2_X1 U958 ( .A1(n887), .A2(G124), .ZN(n859) );
  XOR2_X1 U959 ( .A(KEYINPUT44), .B(n859), .Z(n860) );
  NOR2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n862) );
  NAND2_X1 U961 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n864), .B(KEYINPUT111), .ZN(G162) );
  NAND2_X1 U963 ( .A1(G130), .A2(n887), .ZN(n866) );
  NAND2_X1 U964 ( .A1(G118), .A2(n889), .ZN(n865) );
  NAND2_X1 U965 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U966 ( .A(KEYINPUT112), .B(n867), .ZN(n872) );
  NAND2_X1 U967 ( .A1(G142), .A2(n883), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G106), .A2(n884), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U970 ( .A(n870), .B(KEYINPUT45), .Z(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(n879) );
  XNOR2_X1 U973 ( .A(KEYINPUT46), .B(KEYINPUT113), .ZN(n877) );
  XNOR2_X1 U974 ( .A(n875), .B(KEYINPUT48), .ZN(n876) );
  XNOR2_X1 U975 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U976 ( .A(n879), .B(n878), .Z(n881) );
  XNOR2_X1 U977 ( .A(G160), .B(G162), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U979 ( .A(n882), .B(n928), .Z(n897) );
  NAND2_X1 U980 ( .A1(G139), .A2(n883), .ZN(n886) );
  NAND2_X1 U981 ( .A1(G103), .A2(n884), .ZN(n885) );
  NAND2_X1 U982 ( .A1(n886), .A2(n885), .ZN(n895) );
  NAND2_X1 U983 ( .A1(n887), .A2(G127), .ZN(n888) );
  XNOR2_X1 U984 ( .A(n888), .B(KEYINPUT114), .ZN(n891) );
  NAND2_X1 U985 ( .A1(G115), .A2(n889), .ZN(n890) );
  NAND2_X1 U986 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U987 ( .A(KEYINPUT47), .B(n892), .ZN(n893) );
  XNOR2_X1 U988 ( .A(KEYINPUT115), .B(n893), .ZN(n894) );
  NOR2_X1 U989 ( .A1(n895), .A2(n894), .ZN(n936) );
  XNOR2_X1 U990 ( .A(G164), .B(n936), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n899) );
  XOR2_X1 U992 ( .A(n899), .B(n898), .Z(n900) );
  NOR2_X1 U993 ( .A1(G37), .A2(n900), .ZN(G395) );
  XOR2_X1 U994 ( .A(KEYINPUT116), .B(n901), .Z(n903) );
  XNOR2_X1 U995 ( .A(G171), .B(n969), .ZN(n902) );
  XNOR2_X1 U996 ( .A(n903), .B(n902), .ZN(n905) );
  XOR2_X1 U997 ( .A(n950), .B(G286), .Z(n904) );
  XNOR2_X1 U998 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U999 ( .A1(G37), .A2(n906), .ZN(G397) );
  XOR2_X1 U1000 ( .A(G2443), .B(G2427), .Z(n908) );
  XNOR2_X1 U1001 ( .A(G2438), .B(G2454), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1003 ( .A(n909), .B(G2435), .Z(n911) );
  XNOR2_X1 U1004 ( .A(G1348), .B(G1341), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1006 ( .A(G2430), .B(G2446), .Z(n913) );
  XNOR2_X1 U1007 ( .A(KEYINPUT104), .B(G2451), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1009 ( .A(n915), .B(n914), .Z(n916) );
  NAND2_X1 U1010 ( .A1(G14), .A2(n916), .ZN(n923) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n923), .ZN(n920) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n917) );
  XOR2_X1 U1013 ( .A(KEYINPUT117), .B(n917), .Z(n918) );
  XNOR2_X1 U1014 ( .A(n918), .B(KEYINPUT49), .ZN(n919) );
  NOR2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G69), .ZN(G235) );
  INV_X1 U1020 ( .A(n923), .ZN(G401) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1023 ( .A(KEYINPUT51), .B(n926), .Z(n943) );
  XNOR2_X1 U1024 ( .A(G2084), .B(G160), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(n927), .B(KEYINPUT118), .ZN(n931) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n935) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n941) );
  XOR2_X1 U1030 ( .A(G2072), .B(n936), .Z(n938) );
  XOR2_X1 U1031 ( .A(G164), .B(G2078), .Z(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1033 ( .A(KEYINPUT50), .B(n939), .Z(n940) );
  NOR2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1036 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n946), .ZN(n947) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n1019) );
  NAND2_X1 U1039 ( .A1(n947), .A2(n1019), .ZN(n948) );
  NAND2_X1 U1040 ( .A1(n948), .A2(G29), .ZN(n1028) );
  XOR2_X1 U1041 ( .A(G16), .B(KEYINPUT56), .Z(n977) );
  XNOR2_X1 U1042 ( .A(G171), .B(G1961), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(n949), .B(KEYINPUT121), .ZN(n975) );
  XOR2_X1 U1044 ( .A(n950), .B(G1341), .Z(n962) );
  XOR2_X1 U1045 ( .A(n951), .B(G1956), .Z(n959) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(KEYINPUT122), .B(n954), .ZN(n956) );
  XOR2_X1 U1048 ( .A(G1971), .B(G166), .Z(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(KEYINPUT123), .B(n957), .ZN(n958) );
  NOR2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(KEYINPUT124), .B(n960), .ZN(n961) );
  NAND2_X1 U1053 ( .A1(n962), .A2(n961), .ZN(n968) );
  XNOR2_X1 U1054 ( .A(G168), .B(G1966), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(n963), .B(KEYINPUT120), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1057 ( .A(KEYINPUT57), .B(n966), .Z(n967) );
  NOR2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n973) );
  XOR2_X1 U1059 ( .A(G1348), .B(n969), .Z(n970) );
  NOR2_X1 U1060 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1061 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1062 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1063 ( .A1(n977), .A2(n976), .ZN(n1025) );
  XNOR2_X1 U1064 ( .A(G1961), .B(G5), .ZN(n979) );
  XNOR2_X1 U1065 ( .A(G21), .B(G1966), .ZN(n978) );
  NOR2_X1 U1066 ( .A1(n979), .A2(n978), .ZN(n991) );
  XOR2_X1 U1067 ( .A(KEYINPUT126), .B(G4), .Z(n981) );
  XNOR2_X1 U1068 ( .A(G1348), .B(KEYINPUT59), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(n981), .B(n980), .ZN(n984) );
  XOR2_X1 U1070 ( .A(KEYINPUT125), .B(G1956), .Z(n982) );
  XNOR2_X1 U1071 ( .A(G20), .B(n982), .ZN(n983) );
  NOR2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n988) );
  XNOR2_X1 U1073 ( .A(G1341), .B(G19), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(G6), .B(G1981), .ZN(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1077 ( .A(KEYINPUT60), .B(n989), .Z(n990) );
  NAND2_X1 U1078 ( .A1(n991), .A2(n990), .ZN(n998) );
  XNOR2_X1 U1079 ( .A(G1971), .B(G22), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(G23), .B(G1976), .ZN(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n995) );
  XOR2_X1 U1082 ( .A(G1986), .B(G24), .Z(n994) );
  NAND2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(KEYINPUT58), .B(n996), .ZN(n997) );
  NOR2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1086 ( .A(KEYINPUT61), .B(n999), .Z(n1000) );
  NOR2_X1 U1087 ( .A1(G16), .A2(n1000), .ZN(n1022) );
  XNOR2_X1 U1088 ( .A(G2067), .B(G26), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(G1991), .B(G25), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1011) );
  XOR2_X1 U1091 ( .A(G2072), .B(G33), .Z(n1003) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(G28), .ZN(n1009) );
  XOR2_X1 U1093 ( .A(n1004), .B(G27), .Z(n1006) );
  XNOR2_X1 U1094 ( .A(G1996), .B(G32), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(n1007), .B(KEYINPUT119), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(n1012), .B(KEYINPUT53), .ZN(n1015) );
  XOR2_X1 U1100 ( .A(G2084), .B(G34), .Z(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT54), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(G35), .B(G2090), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(n1019), .B(n1018), .ZN(n1020) );
  NOR2_X1 U1106 ( .A1(G29), .A2(n1020), .ZN(n1021) );
  NOR2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1108 ( .A1(G11), .A2(n1023), .ZN(n1024) );
  NOR2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1110 ( .A(KEYINPUT127), .B(n1026), .Z(n1027) );
  NAND2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1029), .ZN(G150) );
  INV_X1 U1113 ( .A(G150), .ZN(G311) );
endmodule

