//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT74), .ZN(new_n189));
  XNOR2_X1  g003(.A(G125), .B(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT16), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  OR3_X1    g006(.A1(new_n192), .A2(KEYINPUT16), .A3(G140), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(G146), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n190), .A2(new_n195), .ZN(new_n196));
  XOR2_X1   g010(.A(G119), .B(G128), .Z(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT24), .B(G110), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n199), .B(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G128), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT23), .A3(G119), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n204), .B(new_n206), .C1(G119), .C2(new_n205), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT75), .B1(new_n207), .B2(G110), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n201), .A2(new_n208), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n207), .A2(KEYINPUT75), .A3(G110), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n194), .B(new_n196), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n191), .A2(new_n193), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n195), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n194), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(G110), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n214), .B(new_n215), .C1(new_n197), .C2(new_n198), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G137), .ZN(new_n218));
  INV_X1    g032(.A(G221), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n219), .A2(new_n187), .A3(G953), .ZN(new_n220));
  XOR2_X1   g034(.A(new_n218), .B(new_n220), .Z(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n211), .A2(new_n216), .A3(new_n221), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G902), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n225), .A2(KEYINPUT25), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT25), .B1(new_n225), .B2(new_n226), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n189), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n189), .A2(G902), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT29), .ZN(new_n233));
  INV_X1    g047(.A(G143), .ZN(new_n234));
  OAI211_X1 g048(.A(KEYINPUT68), .B(KEYINPUT1), .C1(new_n234), .C2(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G128), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n195), .A2(G143), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT68), .B1(new_n237), .B2(KEYINPUT1), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(G146), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n234), .A2(KEYINPUT64), .A3(G146), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n242), .A2(new_n243), .B1(G143), .B2(new_n195), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT69), .B1(new_n239), .B2(new_n244), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n234), .A2(KEYINPUT64), .A3(G146), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT64), .B1(new_n234), .B2(G146), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n237), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n248), .B(new_n249), .C1(new_n238), .C2(new_n236), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n237), .A3(new_n240), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT67), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n251), .A2(new_n237), .A3(new_n240), .A4(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n245), .A2(new_n250), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G137), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT65), .A2(G134), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT65), .A2(G134), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT11), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  OR2_X1    g078(.A1(KEYINPUT65), .A2(G134), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT65), .A2(G134), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(G137), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n258), .A2(KEYINPUT66), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT66), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G137), .ZN(new_n270));
  AND2_X1   g084(.A1(KEYINPUT11), .A2(G134), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n263), .A2(new_n264), .A3(new_n267), .A4(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n261), .ZN(new_n274));
  AOI21_X1  g088(.A(G134), .B1(new_n268), .B2(new_n270), .ZN(new_n275));
  OAI21_X1  g089(.A(G131), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n257), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n203), .A2(G116), .ZN(new_n279));
  INV_X1    g093(.A(G116), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G119), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT2), .B(G113), .ZN(new_n283));
  OR2_X1    g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n283), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n265), .A2(new_n266), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT11), .B1(new_n288), .B2(new_n258), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n267), .A2(new_n272), .ZN(new_n290));
  OAI21_X1  g104(.A(G131), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n273), .ZN(new_n292));
  AND2_X1   g106(.A1(KEYINPUT0), .A2(G128), .ZN(new_n293));
  NOR2_X1   g107(.A1(KEYINPUT0), .A2(G128), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n237), .A2(new_n240), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n248), .A2(new_n295), .B1(new_n297), .B2(new_n293), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n278), .A2(new_n287), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT28), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g116(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n303));
  INV_X1    g117(.A(G237), .ZN(new_n304));
  INV_X1    g118(.A(G953), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(G210), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n303), .B(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT26), .B(G101), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n273), .A2(new_n276), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n248), .B1(new_n238), .B2(new_n236), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n312), .A2(KEYINPUT69), .B1(new_n255), .B2(new_n253), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n311), .B1(new_n313), .B2(new_n250), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n297), .A2(new_n293), .ZN(new_n315));
  INV_X1    g129(.A(new_n295), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n315), .B1(new_n244), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(new_n291), .B2(new_n273), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n286), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n301), .B1(new_n319), .B2(new_n300), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n233), .B1(new_n310), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n309), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n278), .A2(new_n299), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n324), .B1(new_n292), .B2(new_n298), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT70), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n326), .A2(new_n278), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n326), .B2(new_n278), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n325), .B(new_n286), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n300), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n321), .B1(new_n322), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n314), .A2(new_n286), .A3(new_n318), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n287), .B1(new_n278), .B2(new_n299), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n319), .A2(KEYINPUT72), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n301), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n322), .B1(new_n300), .B2(new_n301), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT29), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n226), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(G472), .B1(new_n332), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT73), .ZN(new_n343));
  INV_X1    g157(.A(G472), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT72), .B1(new_n319), .B2(new_n300), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n335), .A2(new_n333), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT28), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n340), .ZN(new_n348));
  AOI21_X1  g162(.A(G902), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT28), .B1(new_n334), .B2(new_n335), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT29), .B1(new_n350), .B2(new_n339), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n326), .A2(new_n278), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT70), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n326), .A2(new_n278), .A3(new_n327), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n257), .A2(new_n277), .B1(new_n292), .B2(new_n298), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n286), .B1(new_n356), .B2(KEYINPUT30), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n334), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n351), .B1(new_n359), .B2(new_n309), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n344), .B1(new_n349), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT73), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n343), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n309), .B1(new_n350), .B2(new_n302), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT31), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n357), .B1(new_n354), .B2(new_n353), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n300), .A2(new_n309), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n368), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n330), .A2(KEYINPUT31), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n365), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(G472), .A2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT32), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n365), .ZN(new_n376));
  AOI211_X1 g190(.A(new_n366), .B(new_n368), .C1(new_n355), .C2(new_n358), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT31), .B1(new_n330), .B2(new_n370), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT32), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(new_n373), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n232), .B1(new_n364), .B2(new_n382), .ZN(new_n383));
  XOR2_X1   g197(.A(KEYINPUT9), .B(G234), .Z(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT77), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n219), .B1(new_n385), .B2(new_n226), .ZN(new_n386));
  XNOR2_X1  g200(.A(G110), .B(G140), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n305), .A2(G227), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n387), .B(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT81), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT12), .B1(new_n292), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n257), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT78), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT78), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G104), .ZN(new_n397));
  AOI21_X1  g211(.A(G107), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G107), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(G104), .ZN(new_n400));
  OAI21_X1  g214(.A(G101), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n402));
  NOR2_X1   g216(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n403));
  OAI211_X1 g217(.A(G104), .B(new_n399), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT3), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n404), .B1(new_n398), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n395), .A2(new_n397), .A3(G107), .ZN(new_n407));
  INV_X1    g221(.A(G101), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n401), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n237), .A2(KEYINPUT1), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G128), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n253), .A2(new_n255), .B1(new_n412), .B2(new_n296), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT80), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n296), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n256), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT78), .B(G104), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT3), .B1(new_n417), .B2(G107), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n418), .A2(new_n408), .A3(new_n404), .A4(new_n407), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT80), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n416), .A2(new_n419), .A3(new_n420), .A4(new_n401), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n393), .A2(new_n410), .B1(new_n414), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n292), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n392), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n414), .A2(new_n421), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n313), .A2(new_n250), .A3(new_n410), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n392), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n292), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT10), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n404), .B(new_n407), .C1(new_n398), .C2(new_n405), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT4), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(G101), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n298), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(G101), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n419), .A3(KEYINPUT4), .ZN(new_n439));
  OAI211_X1 g253(.A(KEYINPUT10), .B(new_n401), .C1(new_n406), .C2(new_n409), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n437), .A2(new_n439), .B1(new_n257), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n432), .A2(new_n442), .A3(new_n423), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n390), .B1(new_n430), .B2(new_n443), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n433), .A2(G101), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT4), .B1(new_n406), .B2(new_n409), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI22_X1  g261(.A1(new_n393), .A2(new_n440), .B1(new_n447), .B2(new_n436), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT10), .B1(new_n414), .B2(new_n421), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n448), .A2(new_n449), .A3(new_n292), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n423), .B1(new_n432), .B2(new_n442), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n450), .A2(new_n451), .A3(new_n389), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT82), .B1(new_n444), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n448), .A2(new_n449), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n389), .B1(new_n454), .B2(new_n423), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n292), .B1(new_n448), .B2(new_n449), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT82), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n450), .B1(new_n429), .B2(new_n424), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n457), .B(new_n458), .C1(new_n459), .C2(new_n390), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n453), .A2(new_n460), .A3(G469), .ZN(new_n461));
  INV_X1    g275(.A(G469), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(new_n226), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n422), .A2(new_n423), .A3(new_n392), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n428), .B1(new_n427), .B2(new_n292), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n443), .B(new_n390), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n389), .B1(new_n450), .B2(new_n451), .ZN(new_n467));
  AOI21_X1  g281(.A(G902), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n463), .B1(new_n468), .B2(new_n462), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n386), .B1(new_n461), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G214), .B1(G237), .B2(G902), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n279), .A2(new_n281), .A3(KEYINPUT5), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n473), .B(G113), .C1(KEYINPUT5), .C2(new_n279), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n419), .A2(new_n284), .A3(new_n401), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n435), .A2(new_n286), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n447), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G110), .B(G122), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n478), .B(new_n475), .C1(new_n447), .C2(new_n476), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(KEYINPUT6), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT6), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n477), .A2(new_n483), .A3(new_n479), .ZN(new_n484));
  AOI21_X1  g298(.A(G125), .B1(new_n313), .B2(new_n250), .ZN(new_n485));
  INV_X1    g299(.A(G224), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(G953), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n298), .A2(G125), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n487), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n257), .A2(new_n192), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n491), .B1(new_n492), .B2(new_n488), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n482), .A2(new_n484), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT83), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n482), .A2(new_n494), .A3(KEYINPUT83), .A4(new_n484), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n491), .A2(KEYINPUT7), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n485), .B2(new_n489), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n492), .A2(new_n488), .A3(new_n499), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n478), .B(KEYINPUT8), .ZN(new_n503));
  INV_X1    g317(.A(new_n475), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n419), .A2(new_n401), .B1(new_n284), .B2(new_n474), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n501), .A2(new_n502), .A3(new_n481), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n226), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n497), .A2(new_n498), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G210), .B1(G237), .B2(G902), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT84), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n508), .B1(new_n495), .B2(new_n496), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n513), .A3(new_n498), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n472), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n304), .A2(new_n305), .A3(G214), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(new_n234), .ZN(new_n520));
  NAND2_X1  g334(.A1(KEYINPUT18), .A2(G131), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n519), .B(G143), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n521), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n190), .B(new_n195), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT85), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n523), .A2(new_n525), .A3(KEYINPUT85), .A4(new_n526), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n520), .A2(KEYINPUT17), .A3(G131), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n531), .A2(new_n213), .A3(new_n194), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n520), .A2(G131), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n524), .A2(new_n264), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n529), .A2(new_n530), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G113), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(new_n394), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT87), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n226), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n529), .A2(new_n530), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n532), .A2(new_n536), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n544), .A2(new_n545), .A3(new_n542), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT88), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n545), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n541), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT88), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n537), .A2(new_n542), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .A4(new_n226), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n547), .A2(G475), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n212), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n533), .A2(new_n534), .B1(new_n554), .B2(G146), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT86), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n190), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT19), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n195), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n539), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n544), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(G475), .A2(G902), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n562), .B(new_n563), .C1(new_n537), .C2(new_n540), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT20), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n548), .A2(new_n539), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT20), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n562), .A4(new_n563), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n553), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G952), .ZN(new_n571));
  AOI211_X1 g385(.A(G953), .B(new_n571), .C1(G234), .C2(G237), .ZN(new_n572));
  AOI211_X1 g386(.A(new_n226), .B(new_n305), .C1(G234), .C2(G237), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT21), .B(G898), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n234), .A2(G128), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n205), .A2(G143), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n288), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n234), .A2(KEYINPUT13), .A3(G128), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT90), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n581), .A3(new_n577), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT13), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n582), .B1(new_n583), .B2(new_n576), .ZN(new_n584));
  OAI21_X1  g398(.A(G134), .B1(new_n580), .B2(new_n581), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT89), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(G122), .ZN(new_n587));
  INV_X1    g401(.A(G122), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(KEYINPUT89), .ZN(new_n589));
  OAI21_X1  g403(.A(G116), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n280), .A2(G122), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n590), .A2(new_n399), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n399), .B1(new_n590), .B2(new_n591), .ZN(new_n593));
  OAI221_X1 g407(.A(new_n579), .B1(new_n584), .B2(new_n585), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n592), .ZN(new_n595));
  INV_X1    g409(.A(new_n590), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n591), .B(KEYINPUT14), .ZN(new_n597));
  OAI21_X1  g411(.A(G107), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n288), .B(new_n578), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n385), .A2(G217), .A3(new_n305), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n602), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(new_n594), .A3(new_n600), .ZN(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(G478), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(KEYINPUT15), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n606), .B(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n570), .A2(new_n575), .A3(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n470), .A2(new_n518), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n383), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  OAI21_X1  g428(.A(KEYINPUT91), .B1(new_n372), .B2(G902), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT91), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n379), .A2(new_n616), .A3(new_n226), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(new_n617), .A3(G472), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT92), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n379), .B2(new_n373), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n615), .A2(new_n617), .A3(new_n619), .A4(G472), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n461), .A2(new_n469), .ZN(new_n624));
  INV_X1    g438(.A(new_n386), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n232), .ZN(new_n627));
  INV_X1    g441(.A(new_n575), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n510), .A2(KEYINPUT93), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT93), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n516), .A2(new_n630), .A3(new_n498), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n629), .A2(new_n512), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n630), .B1(new_n516), .B2(new_n498), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n472), .B1(new_n633), .B2(new_n511), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n553), .A2(new_n569), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n607), .A2(G902), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n605), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n604), .B1(new_n594), .B2(new_n600), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT33), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n603), .A2(new_n641), .A3(new_n605), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n637), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT94), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT94), .B1(new_n606), .B2(G478), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n645), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n635), .A2(new_n647), .ZN(new_n648));
  AND4_X1   g462(.A1(new_n628), .A2(new_n632), .A3(new_n634), .A4(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n623), .A2(new_n627), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n394), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT95), .B(KEYINPUT34), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  INV_X1    g467(.A(KEYINPUT96), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n565), .A2(new_n568), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n564), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n655), .A2(new_n553), .A3(new_n610), .A4(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n575), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n632), .A2(new_n634), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT97), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n623), .A3(new_n627), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(new_n399), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT98), .B(KEYINPUT35), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  NOR2_X1   g479(.A1(new_n222), .A2(KEYINPUT36), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n217), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n230), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n229), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n623), .A2(new_n612), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  NOR2_X1   g486(.A1(new_n361), .A2(new_n362), .ZN(new_n673));
  AOI211_X1 g487(.A(KEYINPUT73), .B(new_n344), .C1(new_n349), .C2(new_n360), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n382), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n470), .A3(new_n669), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n632), .A2(new_n634), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n573), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n572), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n657), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n676), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(new_n205), .ZN(G30));
  XOR2_X1   g501(.A(new_n682), .B(KEYINPUT39), .Z(new_n688));
  NOR2_X1   g502(.A1(new_n626), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT40), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT99), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT40), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n689), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT99), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n331), .A2(new_n309), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n336), .A2(new_n322), .A3(new_n337), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n226), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G472), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n669), .B1(new_n382), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n610), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n635), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n700), .A2(new_n471), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n515), .A2(new_n517), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT38), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n692), .A2(new_n695), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G143), .ZN(G45));
  NOR3_X1   g523(.A1(new_n635), .A2(new_n647), .A3(new_n683), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n632), .A2(new_n634), .A3(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(new_n675), .A3(new_n470), .A4(new_n669), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  NAND2_X1  g527(.A1(new_n456), .A2(new_n443), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n430), .A2(new_n455), .B1(new_n714), .B2(new_n389), .ZN(new_n715));
  OAI21_X1  g529(.A(G469), .B1(new_n715), .B2(G902), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n466), .A2(new_n467), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n462), .A3(new_n226), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n716), .A2(new_n625), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT100), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT100), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n716), .A2(new_n718), .A3(new_n721), .A4(new_n625), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n383), .A2(new_n649), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND3_X1  g540(.A1(new_n661), .A2(new_n383), .A3(new_n723), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT101), .B(G116), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G18));
  INV_X1    g543(.A(new_n669), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n364), .B2(new_n382), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n723), .A3(new_n611), .A4(new_n678), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  AND3_X1   g547(.A1(new_n632), .A2(new_n634), .A3(new_n702), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n723), .A2(new_n628), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n369), .A2(new_n371), .ZN(new_n737));
  INV_X1    g551(.A(new_n302), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n322), .B1(new_n338), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n374), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(G472), .B1(new_n372), .B2(G902), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n740), .B1(new_n741), .B2(KEYINPUT102), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT102), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n743), .B(G472), .C1(new_n372), .C2(G902), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n736), .B1(new_n745), .B2(new_n232), .ZN(new_n746));
  INV_X1    g560(.A(new_n232), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n742), .A2(new_n747), .A3(KEYINPUT103), .A4(new_n744), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n735), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n588), .ZN(G24));
  NAND4_X1  g564(.A1(new_n742), .A2(new_n669), .A3(new_n710), .A4(new_n744), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n720), .A2(new_n632), .A3(new_n634), .A4(new_n722), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n192), .ZN(G27));
  OR2_X1    g568(.A1(new_n383), .A2(KEYINPUT107), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n383), .A2(KEYINPUT107), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n515), .A2(new_n471), .A3(new_n517), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n457), .B(G469), .C1(new_n459), .C2(new_n390), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n463), .B(KEYINPUT104), .Z(new_n759));
  NAND3_X1  g573(.A1(new_n718), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n625), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT105), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n757), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n760), .A2(KEYINPUT105), .A3(new_n625), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n710), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n755), .A2(new_n756), .A3(new_n765), .A4(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n383), .A2(new_n710), .A3(new_n764), .A4(new_n763), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n770), .A2(KEYINPUT106), .A3(new_n767), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT106), .B1(new_n770), .B2(new_n767), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G131), .ZN(G33));
  NAND3_X1  g588(.A1(new_n765), .A2(new_n383), .A3(new_n684), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  AOI21_X1  g590(.A(KEYINPUT45), .B1(new_n453), .B2(new_n460), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n444), .A2(new_n452), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n462), .B1(new_n779), .B2(KEYINPUT45), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n759), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT46), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n781), .A2(KEYINPUT46), .A3(new_n759), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n718), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n625), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n688), .ZN(new_n788));
  INV_X1    g602(.A(new_n623), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n643), .A2(new_n646), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n644), .B2(new_n643), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n635), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n790), .B1(new_n793), .B2(KEYINPUT108), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT43), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n795), .B1(new_n793), .B2(new_n790), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n794), .A2(KEYINPUT43), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n789), .B(new_n669), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n757), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n788), .B(new_n801), .C1(new_n800), .C2(new_n799), .ZN(new_n802));
  XOR2_X1   g616(.A(KEYINPUT110), .B(G137), .Z(new_n803));
  XNOR2_X1  g617(.A(new_n802), .B(new_n803), .ZN(G39));
  XNOR2_X1  g618(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n787), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n786), .A2(new_n625), .A3(new_n805), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n343), .A2(new_n363), .B1(new_n375), .B2(new_n381), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n747), .A2(new_n766), .A3(new_n757), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  NAND2_X1  g627(.A1(new_n716), .A2(new_n718), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n807), .B(new_n808), .C1(new_n625), .C2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n572), .B1(new_n798), .B2(new_n797), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(new_n746), .B2(new_n748), .ZN(new_n817));
  INV_X1    g631(.A(new_n757), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT116), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n706), .A2(new_n723), .A3(new_n472), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n706), .A2(new_n723), .A3(KEYINPUT117), .A4(new_n472), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(KEYINPUT50), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n817), .A2(new_n823), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n723), .A2(new_n818), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n816), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n745), .A2(new_n730), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n382), .A2(new_n699), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n828), .A2(new_n232), .A3(new_n681), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n792), .A2(new_n570), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n829), .A2(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n794), .A2(new_n796), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n794), .A2(KEYINPUT43), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n681), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n746), .A2(new_n748), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n823), .A2(new_n837), .A3(new_n838), .A4(new_n824), .ZN(new_n839));
  INV_X1    g653(.A(new_n826), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n825), .A2(KEYINPUT50), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n827), .A2(new_n834), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n820), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n815), .A2(KEYINPUT116), .A3(new_n819), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT51), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n815), .B2(new_n819), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n827), .A2(new_n834), .A3(new_n842), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n752), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n817), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n755), .A2(new_n756), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n853), .A2(new_n816), .A3(new_n828), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT48), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT119), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n855), .A2(KEYINPUT119), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n854), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  AOI211_X1 g674(.A(new_n571), .B(G953), .C1(new_n832), .C2(new_n648), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n850), .A2(new_n852), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT120), .B1(new_n846), .B2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n857), .A2(new_n852), .A3(new_n861), .A4(new_n859), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n849), .B2(new_n848), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n866));
  INV_X1    g680(.A(new_n845), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n867), .A2(new_n820), .A3(new_n843), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n865), .B(new_n866), .C1(new_n868), .C2(KEYINPUT51), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n863), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n655), .A2(new_n553), .A3(new_n656), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n818), .A2(new_n701), .A3(new_n871), .A4(new_n682), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n872), .A2(KEYINPUT113), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n810), .A2(new_n626), .A3(new_n730), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(KEYINPUT113), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n751), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n765), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n775), .A3(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n763), .A2(new_n675), .A3(new_n747), .A4(new_n764), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n767), .B1(new_n880), .B2(new_n766), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT106), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n770), .A2(KEYINPUT106), .A3(new_n767), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n879), .B1(new_n885), .B2(new_n769), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n659), .B(KEYINPUT97), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n383), .A2(new_n723), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n732), .B(new_n724), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n569), .A2(new_n553), .A3(new_n610), .A4(new_n628), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n516), .A2(new_n513), .A3(new_n498), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n513), .B1(new_n516), .B2(new_n498), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n890), .B(new_n471), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT112), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n518), .A2(new_n648), .A3(new_n628), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n518), .A2(KEYINPUT112), .A3(new_n890), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(new_n623), .A3(new_n627), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n613), .A3(new_n670), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n889), .A2(new_n900), .A3(new_n749), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n677), .A2(new_n657), .A3(new_n683), .ZN(new_n902));
  AOI22_X1  g716(.A1(new_n874), .A2(new_n902), .B1(new_n877), .B2(new_n851), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n761), .A2(new_n683), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n734), .A2(new_n700), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n712), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n903), .A2(new_n906), .A3(KEYINPUT52), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT114), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT52), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n676), .A2(new_n685), .B1(new_n752), .B2(new_n751), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n712), .A2(new_n905), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n907), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n908), .B1(new_n907), .B2(new_n912), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n886), .B(new_n901), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT53), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n907), .A2(new_n912), .ZN(new_n917));
  INV_X1    g731(.A(new_n879), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n900), .A2(new_n916), .ZN(new_n919));
  AND4_X1   g733(.A1(new_n773), .A2(new_n917), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n838), .A2(new_n628), .A3(new_n723), .A4(new_n734), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n732), .A2(new_n724), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT115), .A4(new_n727), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT115), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n889), .B2(new_n749), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  AOI22_X1  g740(.A1(new_n915), .A2(new_n916), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT54), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n901), .A2(new_n773), .A3(new_n918), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(new_n916), .A3(new_n917), .ZN(new_n931));
  INV_X1    g745(.A(new_n915), .ZN(new_n932));
  OAI211_X1 g746(.A(KEYINPUT54), .B(new_n931), .C1(new_n932), .C2(new_n916), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  OAI22_X1  g748(.A1(new_n870), .A2(new_n934), .B1(G952), .B2(G953), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n814), .B(KEYINPUT49), .Z(new_n936));
  NOR4_X1   g750(.A1(new_n232), .A2(new_n793), .A3(new_n386), .A4(new_n472), .ZN(new_n937));
  INV_X1    g751(.A(new_n831), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n936), .A2(new_n706), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n935), .A2(new_n939), .ZN(G75));
  NOR2_X1   g754(.A1(new_n305), .A2(G952), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n913), .A2(new_n914), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n901), .A2(new_n773), .A3(new_n918), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n916), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n920), .A2(new_n926), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n226), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT56), .B1(new_n947), .B2(G210), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n482), .A2(new_n484), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(new_n494), .Z(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT55), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n942), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n948), .A2(new_n951), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT121), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT121), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n948), .A2(new_n955), .A3(new_n951), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n952), .B1(new_n954), .B2(new_n956), .ZN(G51));
  XOR2_X1   g771(.A(new_n759), .B(KEYINPUT57), .Z(new_n958));
  NAND4_X1  g772(.A1(new_n945), .A2(KEYINPUT122), .A3(new_n946), .A4(new_n928), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT52), .B1(new_n903), .B2(new_n906), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n910), .A2(new_n911), .A3(new_n909), .ZN(new_n961));
  OAI21_X1  g775(.A(KEYINPUT114), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n907), .A2(new_n908), .A3(new_n912), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT53), .B1(new_n930), .B2(new_n964), .ZN(new_n965));
  AND4_X1   g779(.A1(new_n886), .A2(new_n926), .A3(new_n917), .A4(new_n919), .ZN(new_n966));
  OAI21_X1  g780(.A(KEYINPUT54), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n959), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT122), .B1(new_n927), .B2(new_n928), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n958), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n717), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n947), .A2(new_n778), .A3(new_n780), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n941), .B1(new_n971), .B2(new_n972), .ZN(G54));
  AND2_X1   g787(.A1(KEYINPUT58), .A2(G475), .ZN(new_n974));
  OAI211_X1 g788(.A(G902), .B(new_n974), .C1(new_n965), .C2(new_n966), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n566), .A2(new_n562), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n945), .A2(new_n946), .ZN(new_n978));
  INV_X1    g792(.A(new_n976), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n978), .A2(G902), .A3(new_n979), .A4(new_n974), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n977), .A2(new_n980), .A3(new_n942), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT123), .ZN(G60));
  NOR2_X1   g796(.A1(new_n968), .A2(new_n969), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n640), .A2(new_n642), .ZN(new_n984));
  NAND2_X1  g798(.A1(G478), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT59), .Z(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n986), .B1(new_n929), .B2(new_n933), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n942), .B1(new_n990), .B2(new_n984), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n989), .A2(new_n991), .ZN(G63));
  NAND2_X1  g806(.A1(G217), .A2(G902), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT124), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT60), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n978), .A2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n225), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n978), .A2(new_n667), .A3(new_n995), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n998), .A2(new_n942), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT61), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n998), .A2(KEYINPUT61), .A3(new_n942), .A4(new_n999), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(G66));
  NOR3_X1   g818(.A1(new_n574), .A2(new_n486), .A3(new_n305), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(new_n901), .B2(new_n305), .ZN(new_n1006));
  INV_X1    g820(.A(G898), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n949), .B1(new_n1007), .B2(G953), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1006), .B(new_n1008), .Z(G69));
  NAND2_X1  g823(.A1(new_n355), .A2(new_n325), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(new_n559), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1011), .B1(G900), .B2(G953), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n910), .B1(new_n874), .B2(new_n711), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n775), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n755), .A2(new_n734), .A3(new_n756), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1014), .B1(new_n788), .B2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1016), .A2(new_n812), .A3(new_n802), .A4(new_n773), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1012), .B1(new_n1017), .B2(G953), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n305), .B1(G227), .B2(G900), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT62), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n708), .A2(new_n1023), .A3(new_n1013), .ZN(new_n1024));
  INV_X1    g838(.A(new_n648), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1025), .B1(new_n570), .B2(new_n701), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n383), .A2(new_n689), .A3(new_n818), .A4(new_n1026), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n812), .A2(new_n1024), .A3(new_n802), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n708), .A2(new_n1013), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT125), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1029), .A2(new_n1030), .A3(KEYINPUT62), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1029), .A2(KEYINPUT62), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(KEYINPUT125), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1028), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1011), .B1(new_n1034), .B2(G953), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1022), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g852(.A(new_n1036), .B(new_n1038), .ZN(G72));
  NOR2_X1   g853(.A1(new_n331), .A2(new_n309), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(new_n696), .ZN(new_n1042));
  NAND2_X1  g856(.A1(G472), .A2(G902), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(KEYINPUT63), .Z(new_n1044));
  XNOR2_X1  g858(.A(new_n1044), .B(KEYINPUT127), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(new_n942), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n931), .B1(new_n932), .B2(new_n916), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1044), .ZN(new_n1049));
  NOR3_X1   g863(.A1(new_n1048), .A2(new_n1049), .A3(new_n1042), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n1034), .A2(new_n309), .A3(new_n331), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1051), .B1(new_n1017), .B2(new_n1041), .ZN(new_n1052));
  AOI211_X1 g866(.A(new_n1047), .B(new_n1050), .C1(new_n1052), .C2(new_n901), .ZN(G57));
endmodule


