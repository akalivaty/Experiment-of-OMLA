//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n463), .A2(G137), .A3(new_n462), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n462), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  OR2_X1    g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n462), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  AND2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  OAI211_X1 g058(.A(G138), .B(new_n462), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n463), .A2(new_n486), .A3(G138), .A4(new_n462), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n482), .C2(new_n483), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n492), .A3(G2104), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n489), .A2(KEYINPUT67), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(KEYINPUT67), .B1(new_n489), .B2(new_n493), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n488), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT68), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n488), .B(new_n498), .C1(new_n494), .C2(new_n495), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(G164));
  NOR2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT69), .B(G651), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT69), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n504), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(new_n501), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT70), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  INV_X1    g097(.A(new_n503), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n519), .A2(G62), .ZN(new_n524));
  AND2_X1   g099(.A1(G75), .A2(G543), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n508), .A2(new_n522), .A3(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  XOR2_X1   g103(.A(KEYINPUT72), .B(G89), .Z(new_n529));
  NAND3_X1  g104(.A1(new_n505), .A2(new_n519), .A3(new_n529), .ZN(new_n530));
  AND3_X1   g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  OAI221_X1 g107(.A(new_n530), .B1(KEYINPUT7), .B2(new_n531), .C1(new_n506), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n519), .A2(KEYINPUT71), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n517), .A2(new_n535), .A3(new_n518), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n534), .A2(G63), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n509), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n533), .A2(new_n539), .ZN(G168));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n534), .A2(new_n536), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(new_n523), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n505), .A2(G52), .A3(G543), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n505), .A2(G90), .A3(new_n519), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n548), .B1(new_n546), .B2(new_n547), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n545), .B1(new_n549), .B2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  AOI22_X1  g127(.A1(G43), .A2(new_n507), .B1(new_n521), .B2(G81), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n542), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(new_n523), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT74), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND3_X1  g139(.A1(new_n505), .A2(G53), .A3(G543), .ZN(new_n565));
  XNOR2_X1  g140(.A(KEYINPUT75), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  XOR2_X1   g143(.A(KEYINPUT77), .B(G65), .Z(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n520), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(KEYINPUT75), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n505), .A2(G53), .A3(G543), .A4(new_n573), .ZN(new_n574));
  AND3_X1   g149(.A1(new_n567), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n505), .A2(G91), .A3(new_n519), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G168), .ZN(G286));
  NAND3_X1  g155(.A1(new_n505), .A2(G49), .A3(G543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n505), .A2(new_n519), .ZN(new_n582));
  INV_X1    g157(.A(G87), .ZN(new_n583));
  AOI21_X1  g158(.A(G74), .B1(new_n534), .B2(new_n536), .ZN(new_n584));
  OAI221_X1 g159(.A(new_n581), .B1(new_n582), .B2(new_n583), .C1(new_n584), .C2(new_n509), .ZN(G288));
  OAI211_X1 g160(.A(G86), .B(new_n519), .C1(new_n513), .C2(new_n501), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT78), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n505), .A2(new_n588), .A3(G86), .A4(new_n519), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n591));
  OAI211_X1 g166(.A(G48), .B(G543), .C1(new_n513), .C2(new_n501), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n517), .B2(new_n518), .ZN(new_n594));
  AND2_X1   g169(.A1(G73), .A2(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n523), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n590), .A2(new_n591), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n591), .B1(new_n590), .B2(new_n597), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(G305));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n602), .A2(new_n506), .B1(new_n582), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n534), .A2(G60), .A3(new_n536), .ZN(new_n606));
  NAND2_X1  g181(.A1(G72), .A2(G543), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n503), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(G290));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n582), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n505), .A2(KEYINPUT10), .A3(G92), .A4(new_n519), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G54), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n519), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n617));
  OAI22_X1  g192(.A1(new_n506), .A2(new_n616), .B1(new_n509), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G171), .B2(new_n621), .ZN(G284));
  OAI21_X1  g198(.A(new_n622), .B1(G171), .B2(new_n621), .ZN(G321));
  NAND2_X1  g199(.A1(G299), .A2(new_n621), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n621), .B2(G168), .ZN(G280));
  XOR2_X1   g201(.A(G280), .B(KEYINPUT80), .Z(G297));
  AOI21_X1  g202(.A(new_n618), .B1(new_n613), .B2(new_n614), .ZN(new_n628));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n553), .A2(new_n557), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(new_n621), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n620), .A2(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(new_n621), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n463), .A2(new_n468), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n474), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n476), .A2(G123), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n462), .A2(G111), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  NAND3_X1  g222(.A1(new_n640), .A2(new_n641), .A3(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT81), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2430), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n655), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2443), .B(G2446), .Z(new_n661));
  OAI21_X1  g236(.A(G14), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT82), .ZN(G401));
  XNOR2_X1  g239(.A(G2084), .B(G2090), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT83), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  AOI21_X1  g245(.A(KEYINPUT18), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2100), .ZN(new_n672));
  NOR2_X1   g247(.A1(G2072), .A2(G2078), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n442), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n668), .B2(KEYINPUT18), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(G2096), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n672), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n680), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT84), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(new_n683), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT20), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NOR2_X1   g273(.A1(G171), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G5), .B2(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(G1961), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G27), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G164), .B2(new_n703), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n702), .B1(new_n705), .B2(G2078), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G2078), .B2(new_n705), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n700), .A2(new_n701), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT92), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n703), .A2(G33), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT89), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT25), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n474), .A2(G139), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n713), .B(new_n714), .C1(new_n462), .C2(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n710), .B1(new_n716), .B2(G29), .ZN(new_n717));
  INV_X1    g292(.A(G2072), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT90), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n698), .A2(G21), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G168), .B2(new_n698), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT91), .B(G1966), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n474), .A2(G141), .B1(G105), .B2(new_n468), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n476), .A2(G129), .ZN(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT26), .Z(new_n728));
  NAND3_X1  g303(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G32), .B(new_n729), .S(G29), .Z(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT27), .B(G1996), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G2084), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT24), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(G34), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(G34), .ZN(new_n736));
  AOI21_X1  g311(.A(G29), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G160), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G29), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n732), .B1(new_n733), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT31), .B(G11), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n742), .A2(G28), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n703), .B1(new_n742), .B2(G28), .ZN(new_n744));
  OAI221_X1 g319(.A(new_n741), .B1(new_n743), .B2(new_n744), .C1(new_n646), .C2(new_n703), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n739), .B2(new_n733), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n717), .B2(new_n718), .ZN(new_n747));
  NOR4_X1   g322(.A1(new_n720), .A2(new_n724), .A3(new_n740), .A4(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n707), .A2(new_n709), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(KEYINPUT93), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n698), .A2(G20), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT23), .Z(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G299), .B2(G16), .ZN(new_n753));
  INV_X1    g328(.A(G1956), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n628), .A2(new_n698), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G4), .B2(new_n698), .ZN(new_n757));
  INV_X1    g332(.A(G1348), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n703), .A2(G26), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT28), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n474), .A2(G140), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n476), .A2(G128), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n462), .A2(G116), .ZN(new_n765));
  OAI21_X1  g340(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n763), .B(new_n764), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n762), .B1(new_n767), .B2(G29), .ZN(new_n768));
  INV_X1    g343(.A(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n703), .A2(G35), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G162), .B2(new_n703), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT29), .B(G2090), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OR4_X1    g349(.A1(new_n759), .A2(new_n760), .A3(new_n770), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n698), .A2(G19), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n558), .B2(new_n698), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1341), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n750), .A2(new_n755), .A3(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n698), .A2(G6), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G305), .B2(G16), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT32), .B(G1981), .Z(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n698), .A2(G22), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G166), .B2(new_n698), .ZN(new_n787));
  INV_X1    g362(.A(G1971), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n698), .A2(G23), .ZN(new_n790));
  INV_X1    g365(.A(G288), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n698), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT33), .B(G1976), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT87), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n792), .B(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n784), .A2(new_n785), .A3(new_n789), .A4(new_n795), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n796), .A2(KEYINPUT34), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(KEYINPUT34), .ZN(new_n798));
  OR2_X1    g373(.A1(G16), .A2(G24), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G290), .B2(new_n698), .ZN(new_n800));
  INV_X1    g375(.A(G1986), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(G95), .A2(G2105), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n803), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT85), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n474), .A2(G131), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n476), .A2(G119), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  MUX2_X1   g383(.A(G25), .B(new_n808), .S(G29), .Z(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT35), .B(G1991), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT86), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n809), .B(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n800), .A2(new_n801), .ZN(new_n813));
  AND2_X1   g388(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n814));
  OR4_X1    g389(.A1(new_n802), .A2(new_n812), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n797), .A2(new_n798), .A3(new_n815), .ZN(new_n816));
  OR3_X1    g391(.A1(new_n816), .A2(KEYINPUT88), .A3(KEYINPUT36), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(KEYINPUT88), .B2(KEYINPUT36), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n749), .A2(KEYINPUT93), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n780), .A2(new_n817), .A3(new_n818), .A4(new_n819), .ZN(G150));
  INV_X1    g395(.A(G150), .ZN(G311));
  XNOR2_X1  g396(.A(KEYINPUT96), .B(G860), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  AOI22_X1  g398(.A1(G55), .A2(new_n507), .B1(new_n521), .B2(G93), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n534), .A2(G67), .A3(new_n536), .ZN(new_n825));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n825), .A2(KEYINPUT94), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(new_n523), .ZN(new_n828));
  AOI21_X1  g403(.A(KEYINPUT94), .B1(new_n825), .B2(new_n826), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n824), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT95), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n824), .B(KEYINPUT95), .C1(new_n828), .C2(new_n829), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n832), .A2(new_n558), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n830), .A2(new_n831), .A3(new_n631), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n628), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT39), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n823), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n840), .B2(new_n839), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n830), .A2(new_n823), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(G145));
  AND2_X1   g420(.A1(new_n489), .A2(new_n493), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n486), .B1(new_n474), .B2(G138), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n767), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n729), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT97), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n716), .B(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n716), .A2(new_n852), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(new_n851), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n808), .B(KEYINPUT98), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n637), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n476), .A2(G130), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n462), .A2(G118), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(G142), .B2(new_n474), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n858), .B(new_n863), .Z(new_n864));
  AOI21_X1  g439(.A(new_n856), .B1(new_n864), .B2(KEYINPUT100), .ZN(new_n865));
  XNOR2_X1  g440(.A(G160), .B(new_n646), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G162), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n864), .A2(KEYINPUT100), .A3(new_n856), .ZN(new_n869));
  AOI21_X1  g444(.A(G37), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n856), .A2(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n856), .A2(new_n871), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n864), .A2(new_n872), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n873), .B(new_n867), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n879));
  AOI22_X1  g454(.A1(G49), .A2(new_n507), .B1(new_n521), .B2(G87), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n584), .A2(new_n509), .ZN(new_n881));
  AOI22_X1  g456(.A1(new_n609), .A2(new_n605), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR3_X1   g457(.A1(G288), .A2(new_n608), .A3(new_n604), .ZN(new_n883));
  INV_X1    g458(.A(new_n600), .ZN(new_n884));
  AOI21_X1  g459(.A(G166), .B1(new_n884), .B2(new_n598), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n599), .A2(G303), .A3(new_n600), .ZN(new_n886));
  OAI221_X1 g461(.A(new_n879), .B1(new_n882), .B2(new_n883), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n879), .B1(new_n882), .B2(new_n883), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n791), .A2(new_n609), .A3(new_n605), .ZN(new_n890));
  NAND2_X1  g465(.A1(G290), .A2(G288), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT102), .ZN(new_n892));
  OAI21_X1  g467(.A(G303), .B1(new_n599), .B2(new_n600), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n888), .A2(new_n889), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n887), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT42), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n836), .B(new_n633), .Z(new_n897));
  XNOR2_X1  g472(.A(new_n576), .B(KEYINPUT76), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n567), .A2(new_n571), .A3(new_n574), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n620), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n628), .A2(new_n578), .A3(new_n575), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT101), .B1(new_n902), .B2(KEYINPUT41), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(KEYINPUT41), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n900), .A2(new_n901), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n905), .B1(new_n909), .B2(KEYINPUT101), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n904), .B1(new_n897), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT103), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n904), .B(new_n913), .C1(new_n897), .C2(new_n910), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n896), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n914), .A2(new_n896), .ZN(new_n916));
  OAI21_X1  g491(.A(G868), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n830), .A2(new_n621), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(G295));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n918), .ZN(G331));
  INV_X1    g495(.A(new_n908), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n907), .B1(new_n900), .B2(new_n901), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT101), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n905), .ZN(new_n924));
  NAND2_X1  g499(.A1(G171), .A2(G168), .ZN(new_n925));
  NAND2_X1  g500(.A1(G286), .A2(G301), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n833), .A2(new_n558), .ZN(new_n928));
  INV_X1    g503(.A(new_n829), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n523), .A3(new_n827), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT95), .B1(new_n930), .B2(new_n824), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n835), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n834), .A2(new_n835), .A3(new_n926), .A4(new_n925), .ZN(new_n935));
  AOI22_X1  g510(.A1(new_n923), .A2(new_n924), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n934), .A2(new_n903), .A3(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n895), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n887), .A2(new_n894), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n903), .A3(new_n935), .ZN(new_n940));
  INV_X1    g515(.A(new_n935), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n834), .A2(new_n835), .B1(new_n926), .B2(new_n925), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n939), .B(new_n940), .C1(new_n943), .C2(new_n910), .ZN(new_n944));
  INV_X1    g519(.A(G37), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n938), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n950), .B(new_n909), .C1(new_n941), .C2(new_n942), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n940), .A2(KEYINPUT105), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n934), .A2(new_n935), .B1(new_n906), .B2(new_n908), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n895), .B(new_n951), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n954), .A2(new_n955), .A3(new_n945), .A4(new_n944), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n944), .A2(new_n945), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n959), .A2(KEYINPUT106), .A3(new_n955), .A4(new_n954), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n946), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n949), .A2(new_n958), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n959), .A2(KEYINPUT43), .A3(new_n954), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n946), .A2(new_n955), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT44), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n964), .A2(new_n967), .ZN(G397));
  AOI21_X1  g543(.A(G1384), .B1(new_n488), .B2(new_n846), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n969), .A2(KEYINPUT45), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n474), .A2(G137), .B1(G101), .B2(new_n468), .ZN(new_n971));
  INV_X1    g546(.A(G125), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n472), .B2(new_n473), .ZN(new_n973));
  INV_X1    g548(.A(new_n465), .ZN(new_n974));
  OAI21_X1  g549(.A(G2105), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT107), .B(G40), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n971), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n970), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n767), .B(new_n769), .ZN(new_n981));
  OR3_X1    g556(.A1(new_n980), .A2(KEYINPUT108), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT108), .B1(new_n980), .B2(new_n981), .ZN(new_n983));
  INV_X1    g558(.A(new_n980), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n729), .B(G1996), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n982), .A2(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n808), .A2(new_n810), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n808), .A2(new_n810), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(G290), .B(G1986), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n990), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT60), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n620), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT119), .ZN(new_n995));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n497), .A2(new_n996), .A3(new_n499), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n849), .A2(new_n999), .A3(new_n996), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(KEYINPUT109), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(new_n969), .B2(new_n999), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n979), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n758), .B1(new_n998), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n979), .A2(new_n969), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(G2067), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n995), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1000), .A2(KEYINPUT109), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n969), .A2(new_n1002), .A3(new_n999), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n978), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1348), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1014), .A2(KEYINPUT119), .A3(new_n1007), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n994), .B1(new_n1009), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n620), .A2(new_n993), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT122), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT61), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT121), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT57), .B1(new_n898), .B2(new_n899), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n575), .A2(new_n1023), .A3(new_n578), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT56), .B(G2072), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n849), .A2(KEYINPUT45), .A3(new_n996), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n979), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n1027), .B(new_n1029), .C1(new_n997), .C2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n497), .A2(new_n999), .A3(new_n996), .A4(new_n499), .ZN(new_n1032));
  INV_X1    g607(.A(new_n969), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n978), .B1(new_n1033), .B2(KEYINPUT50), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1956), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1025), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1029), .B1(new_n997), .B2(new_n1030), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n1026), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n754), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1021), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1044));
  NOR2_X1   g619(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1006), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT58), .B(G1341), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G1996), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1049), .B1(new_n1037), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1046), .B1(new_n1051), .B2(new_n631), .ZN(new_n1052));
  AOI211_X1 g627(.A(G1996), .B(new_n1029), .C1(new_n997), .C2(new_n1030), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n558), .B(new_n1044), .C1(new_n1053), .C2(new_n1049), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1043), .A2(new_n1055), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1020), .A2(KEYINPUT121), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1031), .A2(new_n1025), .A3(new_n1035), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1039), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1021), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1018), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1062), .B(new_n994), .C1(new_n1009), .C2(new_n1015), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1019), .A2(new_n1056), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1009), .A2(new_n1015), .A3(new_n620), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1042), .B1(new_n1066), .B2(new_n1059), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1065), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n701), .B1(new_n998), .B2(new_n1004), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n996), .A4(new_n499), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n978), .B1(new_n1033), .B2(new_n1030), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(G2078), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1071), .A2(new_n1072), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(G1961), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT124), .B1(new_n1080), .B2(new_n1077), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n997), .A2(new_n1030), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1029), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1075), .B1(new_n1085), .B2(G2078), .ZN(new_n1086));
  AOI21_X1  g661(.A(G301), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n1088));
  NAND3_X1  g663(.A1(G160), .A2(new_n1088), .A3(G40), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n971), .A2(new_n975), .A3(G40), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT125), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1089), .A2(new_n1091), .B1(KEYINPUT45), .B2(new_n969), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT126), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1076), .B1(new_n969), .B2(KEYINPUT45), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1092), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1093), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1086), .A2(new_n1098), .A3(new_n1071), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(G171), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1070), .B1(new_n1087), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1082), .A2(G301), .A3(new_n1086), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1070), .B1(new_n1099), .B2(G171), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1012), .A2(new_n1013), .A3(new_n733), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1105));
  INV_X1    g680(.A(G1966), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1104), .A2(new_n1107), .A3(G168), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G8), .ZN(new_n1109));
  AOI21_X1  g684(.A(G168), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT51), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1112), .A3(G8), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1102), .A2(new_n1103), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(G303), .A2(G8), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT55), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n1117));
  AOI21_X1  g692(.A(G2090), .B1(new_n1040), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1032), .A2(new_n1034), .A3(KEYINPUT115), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1118), .A2(new_n1119), .B1(new_n788), .B2(new_n1085), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT116), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(G8), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1116), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1085), .A2(new_n788), .ZN(new_n1125));
  INV_X1    g700(.A(G2090), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1012), .A2(new_n1013), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1116), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(G8), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT110), .ZN(new_n1131));
  INV_X1    g706(.A(G8), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT110), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(new_n1134), .A3(new_n1129), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT112), .B(G1981), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n590), .A2(new_n597), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n592), .A2(new_n586), .A3(new_n596), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT113), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1138), .A2(new_n1139), .A3(G1981), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1138), .B2(G1981), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1137), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT49), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1137), .B(KEYINPUT49), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1047), .A2(new_n1132), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(G1976), .ZN(new_n1148));
  OAI211_X1 g723(.A(G8), .B(new_n1006), .C1(G288), .C2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(KEYINPUT111), .A2(KEYINPUT52), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n880), .A2(G1976), .A3(new_n881), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1150), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1152), .A2(G8), .A3(new_n1006), .A4(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT52), .ZN(new_n1155));
  NAND3_X1  g730(.A1(G288), .A2(new_n1155), .A3(new_n1148), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1151), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1147), .A2(new_n1157), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1158), .A2(KEYINPUT117), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(KEYINPUT117), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1131), .A2(new_n1135), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1101), .A2(new_n1114), .A3(new_n1124), .A4(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1068), .A2(new_n1069), .A3(new_n1162), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1147), .A2(new_n1148), .A3(new_n791), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1137), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1146), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1131), .A2(new_n1135), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1147), .A2(new_n1157), .A3(KEYINPUT114), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT114), .B1(new_n1147), .B2(new_n1157), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1168), .A2(new_n1169), .A3(KEYINPUT63), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1166), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  OAI22_X1  g746(.A1(new_n1168), .A2(new_n1169), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT118), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI221_X1 g749(.A(KEYINPUT118), .B1(new_n1133), .B2(new_n1129), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1132), .B(G286), .C1(new_n1104), .C2(new_n1107), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1171), .B1(new_n1177), .B2(KEYINPUT63), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT63), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1072), .B1(new_n1071), .B2(new_n1078), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1080), .A2(KEYINPUT124), .A3(new_n1077), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1086), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(G171), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1184), .B1(KEYINPUT62), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1111), .A2(new_n1187), .A3(new_n1113), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1180), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1161), .A2(new_n1124), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1178), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n992), .B1(new_n1163), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n981), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n984), .B1(new_n729), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT46), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1195), .B1(new_n984), .B2(new_n1050), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n980), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  XOR2_X1   g773(.A(new_n1198), .B(KEYINPUT47), .Z(new_n1199));
  NOR3_X1   g774(.A1(new_n980), .A2(G290), .A3(G1986), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT127), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT48), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1202), .A2(new_n990), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n986), .A2(new_n988), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1204), .B1(G2067), .B2(new_n767), .ZN(new_n1205));
  AOI211_X1 g780(.A(new_n1199), .B(new_n1203), .C1(new_n984), .C2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1192), .A2(new_n1206), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g782(.A(G319), .ZN(new_n1209));
  NOR4_X1   g783(.A1(G229), .A2(new_n1209), .A3(new_n663), .A4(G227), .ZN(new_n1210));
  NAND3_X1  g784(.A1(new_n962), .A2(new_n877), .A3(new_n1210), .ZN(G225));
  INV_X1    g785(.A(G225), .ZN(G308));
endmodule


