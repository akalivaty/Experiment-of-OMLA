

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764;

  BUF_X1 U366 ( .A(n718), .Z(n346) );
  XNOR2_X1 U367 ( .A(n597), .B(KEYINPUT33), .ZN(n718) );
  XNOR2_X1 U368 ( .A(n440), .B(n347), .ZN(n697) );
  NOR2_X1 U369 ( .A1(n738), .A2(G902), .ZN(n523) );
  XNOR2_X1 U370 ( .A(n467), .B(n466), .ZN(n554) );
  OR2_X1 U371 ( .A1(n731), .A2(n625), .ZN(n467) );
  XNOR2_X1 U372 ( .A(n397), .B(n651), .ZN(n731) );
  NOR2_X2 U373 ( .A1(n612), .A2(n502), .ZN(n503) );
  NOR2_X2 U374 ( .A1(G953), .A2(G237), .ZN(n509) );
  XNOR2_X1 U375 ( .A(G113), .B(G143), .ZN(n489) );
  AND2_X1 U376 ( .A1(n408), .A2(n413), .ZN(n558) );
  NAND2_X2 U377 ( .A1(n401), .A2(n605), .ZN(n685) );
  INV_X2 U378 ( .A(G143), .ZN(n445) );
  NAND2_X4 U379 ( .A1(n380), .A2(n376), .ZN(n704) );
  NAND2_X1 U380 ( .A1(n665), .A2(n681), .ZN(n370) );
  AND2_X1 U381 ( .A1(n550), .A2(KEYINPUT110), .ZN(n409) );
  NOR2_X1 U382 ( .A1(n567), .A2(n566), .ZN(n675) );
  INV_X1 U383 ( .A(n369), .ZN(n741) );
  AND2_X1 U384 ( .A1(n634), .A2(n627), .ZN(n356) );
  XNOR2_X1 U385 ( .A(n558), .B(KEYINPUT36), .ZN(n401) );
  XNOR2_X1 U386 ( .A(n373), .B(n372), .ZN(n763) );
  XNOR2_X1 U387 ( .A(n537), .B(n536), .ZN(n701) );
  XNOR2_X1 U388 ( .A(n439), .B(n438), .ZN(n530) );
  XNOR2_X1 U389 ( .A(n454), .B(G104), .ZN(n521) );
  XNOR2_X1 U390 ( .A(G110), .B(G107), .ZN(n454) );
  NOR2_X2 U391 ( .A1(n718), .A2(n426), .ZN(n598) );
  OR2_X1 U392 ( .A1(n637), .A2(n367), .ZN(n657) );
  NAND2_X1 U393 ( .A1(n701), .A2(n700), .ZN(n698) );
  INV_X1 U394 ( .A(G134), .ZN(n475) );
  NAND2_X1 U395 ( .A1(n468), .A2(G214), .ZN(n687) );
  NAND2_X1 U396 ( .A1(n548), .A2(n700), .ZN(n564) );
  NOR2_X1 U397 ( .A1(n560), .A2(n701), .ZN(n548) );
  INV_X1 U398 ( .A(G469), .ZN(n388) );
  NAND2_X1 U399 ( .A1(n603), .A2(n759), .ZN(n622) );
  XNOR2_X1 U400 ( .A(G902), .B(KEYINPUT92), .ZN(n462) );
  INV_X1 U401 ( .A(G237), .ZN(n463) );
  INV_X1 U402 ( .A(G131), .ZN(n488) );
  XNOR2_X1 U403 ( .A(G104), .B(G122), .ZN(n492) );
  XNOR2_X1 U404 ( .A(n405), .B(G140), .ZN(n493) );
  INV_X1 U405 ( .A(KEYINPUT12), .ZN(n405) );
  XOR2_X1 U406 ( .A(KEYINPUT11), .B(KEYINPUT101), .Z(n487) );
  XNOR2_X1 U407 ( .A(G146), .B(G125), .ZN(n494) );
  XNOR2_X1 U408 ( .A(n419), .B(n417), .ZN(n562) );
  XNOR2_X1 U409 ( .A(n497), .B(n418), .ZN(n417) );
  OR2_X1 U410 ( .A1(n655), .A2(G902), .ZN(n419) );
  INV_X1 U411 ( .A(G475), .ZN(n418) );
  XNOR2_X1 U412 ( .A(n353), .B(n633), .ZN(n637) );
  NOR2_X1 U413 ( .A1(n693), .A2(n690), .ZN(n577) );
  XNOR2_X1 U414 ( .A(n386), .B(n581), .ZN(n587) );
  NOR2_X1 U415 ( .A1(n580), .A2(n579), .ZN(n386) );
  NOR2_X1 U416 ( .A1(n564), .A2(n615), .ZN(n442) );
  AND2_X1 U417 ( .A1(n382), .A2(n381), .ZN(n380) );
  NAND2_X1 U418 ( .A1(n379), .A2(n378), .ZN(n377) );
  AND2_X1 U419 ( .A1(n613), .A2(KEYINPUT97), .ZN(n430) );
  AND2_X1 U420 ( .A1(n428), .A2(n615), .ZN(n427) );
  OR2_X1 U421 ( .A1(n613), .A2(KEYINPUT97), .ZN(n428) );
  INV_X1 U422 ( .A(n614), .ZN(n426) );
  XNOR2_X1 U423 ( .A(n483), .B(n482), .ZN(n742) );
  XNOR2_X1 U424 ( .A(n481), .B(n480), .ZN(n483) );
  XNOR2_X1 U425 ( .A(n522), .B(n399), .ZN(n398) );
  INV_X1 U426 ( .A(n521), .ZN(n399) );
  XNOR2_X1 U427 ( .A(n728), .B(KEYINPUT87), .ZN(n360) );
  NOR2_X1 U428 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U429 ( .A1(n616), .A2(n433), .ZN(n432) );
  XNOR2_X1 U430 ( .A(n619), .B(KEYINPUT107), .ZN(n620) );
  INV_X1 U431 ( .A(KEYINPUT90), .ZN(n395) );
  INV_X1 U432 ( .A(KEYINPUT44), .ZN(n392) );
  XNOR2_X1 U433 ( .A(n635), .B(KEYINPUT80), .ZN(n355) );
  XNOR2_X1 U434 ( .A(n436), .B(G140), .ZN(n526) );
  INV_X1 U435 ( .A(G137), .ZN(n436) );
  NAND2_X1 U436 ( .A1(n688), .A2(n687), .ZN(n693) );
  NAND2_X1 U437 ( .A1(G234), .A2(G237), .ZN(n470) );
  XNOR2_X1 U438 ( .A(n575), .B(n371), .ZN(n688) );
  INV_X1 U439 ( .A(KEYINPUT38), .ZN(n371) );
  NAND2_X1 U440 ( .A1(n564), .A2(KEYINPUT110), .ZN(n412) );
  NAND2_X1 U441 ( .A1(G902), .A2(G472), .ZN(n381) );
  XNOR2_X1 U442 ( .A(KEYINPUT4), .B(G131), .ZN(n504) );
  XOR2_X1 U443 ( .A(KEYINPUT3), .B(G116), .Z(n458) );
  XNOR2_X1 U444 ( .A(G113), .B(G101), .ZN(n457) );
  XNOR2_X1 U445 ( .A(G110), .B(KEYINPUT81), .ZN(n527) );
  INV_X1 U446 ( .A(KEYINPUT8), .ZN(n438) );
  NAND2_X1 U447 ( .A1(n755), .A2(G234), .ZN(n439) );
  XNOR2_X1 U448 ( .A(G116), .B(G107), .ZN(n477) );
  XOR2_X1 U449 ( .A(KEYINPUT104), .B(G122), .Z(n478) );
  XNOR2_X1 U450 ( .A(n495), .B(n496), .ZN(n655) );
  XNOR2_X1 U451 ( .A(n491), .B(n490), .ZN(n496) );
  XOR2_X1 U452 ( .A(G146), .B(G101), .Z(n520) );
  XNOR2_X1 U453 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n446) );
  OR2_X1 U454 ( .A1(n550), .A2(n414), .ZN(n413) );
  NAND2_X1 U455 ( .A1(n415), .A2(n416), .ZN(n414) );
  INV_X1 U456 ( .A(KEYINPUT0), .ZN(n421) );
  NOR2_X1 U457 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U458 ( .A(n383), .B(KEYINPUT30), .ZN(n559) );
  NAND2_X1 U459 ( .A1(n704), .A2(n687), .ZN(n383) );
  BUF_X1 U460 ( .A(n697), .Z(n404) );
  XNOR2_X1 U461 ( .A(KEYINPUT105), .B(G478), .ZN(n484) );
  BUF_X1 U462 ( .A(n701), .Z(n403) );
  NAND2_X1 U463 ( .A1(n365), .A2(n362), .ZN(n361) );
  INV_X1 U464 ( .A(G210), .ZN(n364) );
  XNOR2_X1 U465 ( .A(KEYINPUT42), .B(KEYINPUT113), .ZN(n372) );
  NAND2_X1 U466 ( .A1(n375), .A2(n374), .ZN(n373) );
  INV_X1 U467 ( .A(n578), .ZN(n374) );
  XNOR2_X1 U468 ( .A(n385), .B(n384), .ZN(n761) );
  INV_X1 U469 ( .A(KEYINPUT40), .ZN(n384) );
  NAND2_X1 U470 ( .A1(n587), .A2(n675), .ZN(n385) );
  NAND2_X1 U471 ( .A1(n607), .A2(n541), .ZN(n542) );
  NAND2_X1 U472 ( .A1(n424), .A2(n423), .ZN(n665) );
  AND2_X1 U473 ( .A1(n429), .A2(n427), .ZN(n424) );
  INV_X1 U474 ( .A(KEYINPUT97), .ZN(n425) );
  INV_X1 U475 ( .A(G217), .ZN(n368) );
  XNOR2_X1 U476 ( .A(n744), .B(n743), .ZN(n352) );
  XNOR2_X1 U477 ( .A(n740), .B(n739), .ZN(n351) );
  XNOR2_X1 U478 ( .A(n358), .B(n357), .ZN(G75) );
  INV_X1 U479 ( .A(KEYINPUT53), .ZN(n357) );
  AND2_X1 U480 ( .A1(n729), .A2(n643), .ZN(n359) );
  XOR2_X1 U481 ( .A(n525), .B(n524), .Z(n347) );
  AND2_X1 U482 ( .A1(n570), .A2(n676), .ZN(n348) );
  BUF_X1 U483 ( .A(n554), .Z(n575) );
  XOR2_X1 U484 ( .A(G119), .B(G128), .Z(n349) );
  AND2_X1 U485 ( .A1(n404), .A2(n592), .ZN(n350) );
  INV_X1 U486 ( .A(G902), .ZN(n378) );
  INV_X1 U487 ( .A(n411), .ZN(n410) );
  NAND2_X1 U488 ( .A1(n412), .A2(n687), .ZN(n411) );
  INV_X1 U489 ( .A(KEYINPUT110), .ZN(n416) );
  INV_X1 U490 ( .A(KEYINPUT47), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n518), .B(n526), .ZN(n749) );
  INV_X1 U492 ( .A(G472), .ZN(n379) );
  XNOR2_X1 U493 ( .A(n391), .B(KEYINPUT74), .ZN(n390) );
  NOR2_X1 U494 ( .A1(n348), .A2(n435), .ZN(n571) );
  NAND2_X1 U495 ( .A1(n360), .A2(n359), .ZN(n358) );
  NOR2_X1 U496 ( .A1(n674), .A2(n432), .ZN(n431) );
  NOR2_X1 U497 ( .A1(n351), .A2(n748), .ZN(G54) );
  NOR2_X1 U498 ( .A1(n352), .A2(n748), .ZN(G63) );
  XNOR2_X1 U499 ( .A(n396), .B(n395), .ZN(n394) );
  NAND2_X1 U500 ( .A1(n354), .A2(n632), .ZN(n353) );
  NAND2_X1 U501 ( .A1(n621), .A2(n620), .ZN(n396) );
  NAND2_X1 U502 ( .A1(n356), .A2(n355), .ZN(n354) );
  XNOR2_X1 U503 ( .A(n361), .B(n640), .ZN(n641) );
  NOR2_X1 U504 ( .A1(n727), .A2(n379), .ZN(n362) );
  NAND2_X1 U505 ( .A1(n365), .A2(n363), .ZN(n733) );
  NOR2_X1 U506 ( .A1(n727), .A2(n364), .ZN(n363) );
  INV_X1 U507 ( .A(n637), .ZN(n365) );
  NAND2_X1 U508 ( .A1(n366), .A2(G475), .ZN(n367) );
  INV_X1 U509 ( .A(n727), .ZN(n366) );
  OR2_X1 U510 ( .A1(n637), .A2(n727), .ZN(n369) );
  NOR2_X1 U511 ( .A1(n369), .A2(n368), .ZN(n746) );
  NAND2_X1 U512 ( .A1(n426), .A2(n425), .ZN(n423) );
  XNOR2_X1 U513 ( .A(n370), .B(KEYINPUT100), .ZN(n617) );
  NAND2_X1 U514 ( .A1(n607), .A2(n350), .ZN(n669) );
  XNOR2_X2 U515 ( .A(n503), .B(n444), .ZN(n607) );
  XNOR2_X2 U516 ( .A(n602), .B(n601), .ZN(n759) );
  NOR2_X2 U517 ( .A1(n596), .A2(n604), .ZN(n597) );
  XOR2_X2 U518 ( .A(n704), .B(n517), .Z(n604) );
  NOR2_X2 U519 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U520 ( .A(n389), .B(KEYINPUT45), .ZN(n634) );
  INV_X1 U521 ( .A(n688), .ZN(n579) );
  NOR2_X1 U522 ( .A1(n761), .A2(n763), .ZN(n583) );
  INV_X1 U523 ( .A(n717), .ZN(n375) );
  OR2_X1 U524 ( .A1(n639), .A2(n377), .ZN(n376) );
  NAND2_X1 U525 ( .A1(n639), .A2(G472), .ZN(n382) );
  NOR2_X1 U526 ( .A1(n698), .A2(n387), .ZN(n613) );
  INV_X1 U527 ( .A(n440), .ZN(n387) );
  XNOR2_X2 U528 ( .A(n523), .B(n388), .ZN(n440) );
  NAND2_X1 U529 ( .A1(n394), .A2(n390), .ZN(n389) );
  NAND2_X1 U530 ( .A1(n393), .A2(n392), .ZN(n391) );
  INV_X1 U531 ( .A(n622), .ZN(n393) );
  XNOR2_X1 U532 ( .A(n453), .B(n452), .ZN(n397) );
  XNOR2_X1 U533 ( .A(n749), .B(n398), .ZN(n738) );
  XNOR2_X1 U534 ( .A(n400), .B(n437), .ZN(n532) );
  XNOR2_X1 U535 ( .A(n402), .B(n529), .ZN(n400) );
  NAND2_X1 U536 ( .A1(n410), .A2(n575), .ZN(n406) );
  NAND2_X1 U537 ( .A1(n755), .A2(G227), .ZN(n519) );
  XNOR2_X2 U538 ( .A(n449), .B(G953), .ZN(n755) );
  NOR2_X2 U539 ( .A1(n697), .A2(n698), .ZN(n610) );
  XNOR2_X1 U540 ( .A(n349), .B(n526), .ZN(n402) );
  NOR2_X1 U541 ( .A1(n409), .A2(n406), .ZN(n408) );
  NAND2_X1 U542 ( .A1(n407), .A2(n413), .ZN(n557) );
  NOR2_X1 U543 ( .A1(n409), .A2(n411), .ZN(n407) );
  INV_X1 U544 ( .A(n564), .ZN(n415) );
  XNOR2_X2 U545 ( .A(n420), .B(n421), .ZN(n612) );
  NOR2_X2 U546 ( .A1(n565), .A2(n474), .ZN(n420) );
  XNOR2_X2 U547 ( .A(n422), .B(n469), .ZN(n565) );
  NAND2_X1 U548 ( .A1(n554), .A2(n687), .ZN(n422) );
  NAND2_X1 U549 ( .A1(n614), .A2(n430), .ZN(n429) );
  NAND2_X1 U550 ( .A1(n434), .A2(n431), .ZN(n435) );
  OR2_X1 U551 ( .A1(n676), .A2(n433), .ZN(n434) );
  NAND2_X1 U552 ( .A1(n530), .A2(G221), .ZN(n437) );
  NAND2_X1 U553 ( .A1(n441), .A2(n440), .ZN(n578) );
  XNOR2_X1 U554 ( .A(n442), .B(KEYINPUT28), .ZN(n441) );
  BUF_X1 U555 ( .A(n634), .Z(n721) );
  XNOR2_X2 U556 ( .A(n542), .B(KEYINPUT32), .ZN(n593) );
  OR2_X1 U557 ( .A1(n755), .A2(G952), .ZN(n734) );
  XOR2_X1 U558 ( .A(n493), .B(n492), .Z(n443) );
  XOR2_X1 U559 ( .A(KEYINPUT67), .B(KEYINPUT22), .Z(n444) );
  INV_X1 U560 ( .A(KEYINPUT73), .ZN(n573) );
  XNOR2_X1 U561 ( .A(n574), .B(n573), .ZN(n585) );
  INV_X1 U562 ( .A(KEYINPUT108), .ZN(n595) );
  XNOR2_X1 U563 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U564 ( .A(n443), .B(n750), .ZN(n495) );
  INV_X1 U565 ( .A(KEYINPUT1), .ZN(n524) );
  XNOR2_X1 U566 ( .A(n485), .B(n484), .ZN(n567) );
  XNOR2_X1 U567 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X2 U568 ( .A(n445), .B(G128), .ZN(n476) );
  XNOR2_X1 U569 ( .A(n476), .B(n494), .ZN(n448) );
  XNOR2_X1 U570 ( .A(n446), .B(KEYINPUT82), .ZN(n447) );
  XNOR2_X1 U571 ( .A(n448), .B(n447), .ZN(n453) );
  XOR2_X1 U572 ( .A(KEYINPUT93), .B(KEYINPUT4), .Z(n451) );
  INV_X1 U573 ( .A(KEYINPUT64), .ZN(n449) );
  NAND2_X1 U574 ( .A1(n755), .A2(G224), .ZN(n450) );
  XNOR2_X1 U575 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U576 ( .A(KEYINPUT76), .B(KEYINPUT16), .ZN(n455) );
  XNOR2_X1 U577 ( .A(n455), .B(G122), .ZN(n456) );
  XNOR2_X1 U578 ( .A(n521), .B(n456), .ZN(n460) );
  XNOR2_X1 U579 ( .A(n457), .B(G119), .ZN(n459) );
  XNOR2_X1 U580 ( .A(n459), .B(n458), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n460), .B(n513), .ZN(n651) );
  INV_X1 U582 ( .A(KEYINPUT15), .ZN(n461) );
  XNOR2_X1 U583 ( .A(n462), .B(n461), .ZN(n625) );
  NAND2_X1 U584 ( .A1(n378), .A2(n463), .ZN(n468) );
  NAND2_X1 U585 ( .A1(n468), .A2(G210), .ZN(n465) );
  INV_X1 U586 ( .A(KEYINPUT84), .ZN(n464) );
  XNOR2_X1 U587 ( .A(n465), .B(n464), .ZN(n466) );
  INV_X1 U588 ( .A(KEYINPUT19), .ZN(n469) );
  XNOR2_X1 U589 ( .A(n470), .B(KEYINPUT94), .ZN(n471) );
  XNOR2_X1 U590 ( .A(KEYINPUT14), .B(n471), .ZN(n472) );
  NAND2_X1 U591 ( .A1(G952), .A2(n472), .ZN(n716) );
  NOR2_X1 U592 ( .A1(n716), .A2(G953), .ZN(n547) );
  NAND2_X1 U593 ( .A1(G902), .A2(n472), .ZN(n543) );
  INV_X1 U594 ( .A(G898), .ZN(n647) );
  NAND2_X1 U595 ( .A1(G953), .A2(n647), .ZN(n650) );
  NOR2_X1 U596 ( .A1(n543), .A2(n650), .ZN(n473) );
  NOR2_X1 U597 ( .A1(n547), .A2(n473), .ZN(n474) );
  XNOR2_X2 U598 ( .A(n476), .B(n475), .ZN(n505) );
  XNOR2_X1 U599 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U600 ( .A(n505), .B(n479), .ZN(n481) );
  XOR2_X1 U601 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n480) );
  NAND2_X1 U602 ( .A1(G217), .A2(n530), .ZN(n482) );
  NOR2_X1 U603 ( .A1(G902), .A2(n742), .ZN(n485) );
  NAND2_X1 U604 ( .A1(G214), .A2(n509), .ZN(n486) );
  XNOR2_X1 U605 ( .A(n487), .B(n486), .ZN(n491) );
  XNOR2_X1 U606 ( .A(n494), .B(KEYINPUT10), .ZN(n750) );
  XNOR2_X1 U607 ( .A(KEYINPUT13), .B(KEYINPUT102), .ZN(n497) );
  NOR2_X1 U608 ( .A1(n567), .A2(n562), .ZN(n576) );
  INV_X1 U609 ( .A(n625), .ZN(n498) );
  NAND2_X1 U610 ( .A1(G234), .A2(n498), .ZN(n499) );
  XNOR2_X1 U611 ( .A(n499), .B(KEYINPUT20), .ZN(n533) );
  NAND2_X1 U612 ( .A1(n533), .A2(G221), .ZN(n501) );
  XOR2_X1 U613 ( .A(KEYINPUT21), .B(KEYINPUT96), .Z(n500) );
  XNOR2_X1 U614 ( .A(n501), .B(n500), .ZN(n700) );
  NAND2_X1 U615 ( .A1(n576), .A2(n700), .ZN(n502) );
  XNOR2_X2 U616 ( .A(n505), .B(n504), .ZN(n518) );
  XOR2_X1 U617 ( .A(KEYINPUT98), .B(KEYINPUT79), .Z(n507) );
  XNOR2_X1 U618 ( .A(KEYINPUT99), .B(KEYINPUT78), .ZN(n506) );
  XNOR2_X1 U619 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U620 ( .A(n518), .B(n508), .ZN(n516) );
  XOR2_X1 U621 ( .A(G146), .B(KEYINPUT5), .Z(n511) );
  NAND2_X1 U622 ( .A1(n509), .A2(G210), .ZN(n510) );
  XNOR2_X1 U623 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U624 ( .A(n512), .B(G137), .Z(n514) );
  XNOR2_X1 U625 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U626 ( .A(n516), .B(n515), .ZN(n639) );
  XOR2_X1 U627 ( .A(KEYINPUT106), .B(KEYINPUT6), .Z(n517) );
  XNOR2_X1 U628 ( .A(n604), .B(KEYINPUT83), .ZN(n540) );
  XNOR2_X1 U629 ( .A(n520), .B(n519), .ZN(n522) );
  INV_X1 U630 ( .A(KEYINPUT68), .ZN(n525) );
  INV_X1 U631 ( .A(n404), .ZN(n605) );
  XOR2_X1 U632 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n528) );
  XNOR2_X1 U633 ( .A(n528), .B(n527), .ZN(n529) );
  INV_X1 U634 ( .A(n750), .ZN(n531) );
  XNOR2_X1 U635 ( .A(n532), .B(n531), .ZN(n745) );
  NAND2_X1 U636 ( .A1(n745), .A2(n378), .ZN(n537) );
  NAND2_X1 U637 ( .A1(n533), .A2(G217), .ZN(n535) );
  XNOR2_X1 U638 ( .A(KEYINPUT25), .B(KEYINPUT95), .ZN(n534) );
  XNOR2_X1 U639 ( .A(n535), .B(n534), .ZN(n536) );
  INV_X1 U640 ( .A(n403), .ZN(n538) );
  NAND2_X1 U641 ( .A1(n605), .A2(n538), .ZN(n539) );
  NOR2_X1 U642 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U643 ( .A(n593), .B(G119), .ZN(G21) );
  NOR2_X1 U644 ( .A1(n755), .A2(n543), .ZN(n544) );
  XNOR2_X1 U645 ( .A(n544), .B(KEYINPUT109), .ZN(n545) );
  NOR2_X1 U646 ( .A1(G900), .A2(n545), .ZN(n546) );
  NOR2_X1 U647 ( .A1(n547), .A2(n546), .ZN(n560) );
  XNOR2_X1 U648 ( .A(n562), .B(KEYINPUT103), .ZN(n566) );
  INV_X1 U649 ( .A(n604), .ZN(n549) );
  NAND2_X1 U650 ( .A1(n675), .A2(n549), .ZN(n550) );
  NOR2_X1 U651 ( .A1(n605), .A2(n557), .ZN(n553) );
  XNOR2_X1 U652 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n551) );
  XNOR2_X1 U653 ( .A(n551), .B(KEYINPUT43), .ZN(n552) );
  XNOR2_X1 U654 ( .A(n553), .B(n552), .ZN(n555) );
  INV_X1 U655 ( .A(n575), .ZN(n556) );
  AND2_X1 U656 ( .A1(n555), .A2(n556), .ZN(n589) );
  XOR2_X1 U657 ( .A(n589), .B(G140), .Z(G42) );
  XNOR2_X1 U658 ( .A(n685), .B(KEYINPUT88), .ZN(n572) );
  NAND2_X1 U659 ( .A1(n613), .A2(n561), .ZN(n580) );
  AND2_X1 U660 ( .A1(n567), .A2(n562), .ZN(n599) );
  NAND2_X1 U661 ( .A1(n575), .A2(n599), .ZN(n563) );
  NOR2_X1 U662 ( .A1(n580), .A2(n563), .ZN(n674) );
  INV_X1 U663 ( .A(n704), .ZN(n615) );
  NOR2_X1 U664 ( .A1(n578), .A2(n565), .ZN(n676) );
  NAND2_X1 U665 ( .A1(n567), .A2(n566), .ZN(n682) );
  INV_X1 U666 ( .A(n675), .ZN(n678) );
  NAND2_X1 U667 ( .A1(n682), .A2(n678), .ZN(n616) );
  INV_X1 U668 ( .A(n616), .ZN(n692) );
  XNOR2_X1 U669 ( .A(KEYINPUT72), .B(KEYINPUT47), .ZN(n568) );
  NOR2_X1 U670 ( .A1(n692), .A2(n568), .ZN(n569) );
  XOR2_X1 U671 ( .A(KEYINPUT77), .B(n569), .Z(n570) );
  NAND2_X1 U672 ( .A1(n572), .A2(n571), .ZN(n574) );
  INV_X1 U673 ( .A(n576), .ZN(n690) );
  XNOR2_X1 U674 ( .A(KEYINPUT41), .B(n577), .ZN(n717) );
  XNOR2_X1 U675 ( .A(KEYINPUT75), .B(KEYINPUT39), .ZN(n581) );
  XNOR2_X1 U676 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n582) );
  XNOR2_X1 U677 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U678 ( .A(n586), .B(KEYINPUT48), .ZN(n591) );
  INV_X1 U679 ( .A(n682), .ZN(n670) );
  NAND2_X1 U680 ( .A1(n587), .A2(n670), .ZN(n588) );
  XOR2_X1 U681 ( .A(KEYINPUT114), .B(n588), .Z(n762) );
  NOR2_X1 U682 ( .A1(n762), .A2(n589), .ZN(n590) );
  AND2_X2 U683 ( .A1(n591), .A2(n590), .ZN(n635) );
  NOR2_X1 U684 ( .A1(n704), .A2(n403), .ZN(n592) );
  NAND2_X1 U685 ( .A1(n593), .A2(n669), .ZN(n594) );
  XNOR2_X1 U686 ( .A(n594), .B(KEYINPUT91), .ZN(n603) );
  XNOR2_X1 U687 ( .A(n610), .B(n595), .ZN(n596) );
  XNOR2_X1 U688 ( .A(n598), .B(KEYINPUT34), .ZN(n600) );
  NAND2_X1 U689 ( .A1(n600), .A2(n599), .ZN(n602) );
  INV_X1 U690 ( .A(KEYINPUT35), .ZN(n601) );
  NAND2_X1 U691 ( .A1(n622), .A2(KEYINPUT44), .ZN(n621) );
  NOR2_X1 U692 ( .A1(n549), .A2(n605), .ZN(n606) );
  NAND2_X1 U693 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U694 ( .A(n608), .B(KEYINPUT89), .ZN(n609) );
  NAND2_X1 U695 ( .A1(n609), .A2(n403), .ZN(n662) );
  NAND2_X1 U696 ( .A1(n704), .A2(n610), .ZN(n707) );
  NOR2_X1 U697 ( .A1(n707), .A2(n612), .ZN(n611) );
  XNOR2_X1 U698 ( .A(n611), .B(KEYINPUT31), .ZN(n681) );
  INV_X1 U699 ( .A(n612), .ZN(n614) );
  NAND2_X1 U700 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n662), .A2(n618), .ZN(n619) );
  NAND2_X1 U702 ( .A1(n625), .A2(KEYINPUT2), .ZN(n624) );
  INV_X1 U703 ( .A(KEYINPUT70), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n628) );
  INV_X1 U705 ( .A(n628), .ZN(n626) );
  OR2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n627) );
  INV_X1 U707 ( .A(n627), .ZN(n631) );
  NAND2_X1 U708 ( .A1(KEYINPUT2), .A2(KEYINPUT70), .ZN(n629) );
  AND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n630) );
  OR2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n632) );
  INV_X1 U711 ( .A(KEYINPUT66), .ZN(n633) );
  AND2_X1 U712 ( .A1(n635), .A2(KEYINPUT2), .ZN(n636) );
  AND2_X1 U713 ( .A1(n636), .A2(n721), .ZN(n727) );
  XNOR2_X1 U714 ( .A(KEYINPUT115), .B(KEYINPUT62), .ZN(n638) );
  XNOR2_X1 U715 ( .A(n639), .B(n638), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n641), .A2(n734), .ZN(n642) );
  XNOR2_X1 U717 ( .A(n642), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U718 ( .A(G953), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n721), .A2(n643), .ZN(n644) );
  XOR2_X1 U720 ( .A(KEYINPUT124), .B(n644), .Z(n649) );
  NAND2_X1 U721 ( .A1(G953), .A2(G224), .ZN(n645) );
  XOR2_X1 U722 ( .A(KEYINPUT61), .B(n645), .Z(n646) );
  NOR2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U724 ( .A1(n649), .A2(n648), .ZN(n653) );
  NAND2_X1 U725 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n653), .B(n652), .ZN(G69) );
  XOR2_X1 U727 ( .A(KEYINPUT69), .B(KEYINPUT59), .Z(n654) );
  XNOR2_X1 U728 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n657), .B(n656), .ZN(n658) );
  NAND2_X1 U730 ( .A1(n658), .A2(n734), .ZN(n661) );
  XNOR2_X1 U731 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n659), .B(KEYINPUT71), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n661), .B(n660), .ZN(G60) );
  XNOR2_X1 U734 ( .A(G101), .B(KEYINPUT116), .ZN(n663) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(G3) );
  NOR2_X1 U736 ( .A1(n678), .A2(n665), .ZN(n664) );
  XOR2_X1 U737 ( .A(G104), .B(n664), .Z(G6) );
  NOR2_X1 U738 ( .A1(n682), .A2(n665), .ZN(n667) );
  XNOR2_X1 U739 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n666) );
  XNOR2_X1 U740 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U741 ( .A(G107), .B(n668), .ZN(G9) );
  XNOR2_X1 U742 ( .A(n669), .B(G110), .ZN(G12) );
  XOR2_X1 U743 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n672) );
  NAND2_X1 U744 ( .A1(n676), .A2(n670), .ZN(n671) );
  XNOR2_X1 U745 ( .A(n672), .B(n671), .ZN(n673) );
  XOR2_X1 U746 ( .A(G128), .B(n673), .Z(G30) );
  XOR2_X1 U747 ( .A(G143), .B(n674), .Z(G45) );
  NAND2_X1 U748 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n677), .B(G146), .ZN(G48) );
  NOR2_X1 U750 ( .A1(n678), .A2(n681), .ZN(n679) );
  XOR2_X1 U751 ( .A(KEYINPUT118), .B(n679), .Z(n680) );
  XNOR2_X1 U752 ( .A(G113), .B(n680), .ZN(G15) );
  NOR2_X1 U753 ( .A1(n682), .A2(n681), .ZN(n684) );
  XNOR2_X1 U754 ( .A(G116), .B(KEYINPUT119), .ZN(n683) );
  XNOR2_X1 U755 ( .A(n684), .B(n683), .ZN(G18) );
  XOR2_X1 U756 ( .A(G125), .B(KEYINPUT37), .Z(n686) );
  XNOR2_X1 U757 ( .A(n685), .B(n686), .ZN(G27) );
  NOR2_X1 U758 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U760 ( .A(n691), .B(KEYINPUT120), .ZN(n695) );
  NOR2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U763 ( .A1(n696), .A2(n346), .ZN(n712) );
  NAND2_X1 U764 ( .A1(n698), .A2(n404), .ZN(n699) );
  XNOR2_X1 U765 ( .A(n699), .B(KEYINPUT50), .ZN(n706) );
  NOR2_X1 U766 ( .A1(n403), .A2(n700), .ZN(n702) );
  XOR2_X1 U767 ( .A(KEYINPUT49), .B(n702), .Z(n703) );
  NOR2_X1 U768 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U769 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U770 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U771 ( .A(KEYINPUT51), .B(n709), .ZN(n710) );
  NOR2_X1 U772 ( .A1(n710), .A2(n717), .ZN(n711) );
  NOR2_X1 U773 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U774 ( .A(n713), .B(KEYINPUT52), .Z(n714) );
  XNOR2_X1 U775 ( .A(KEYINPUT121), .B(n714), .ZN(n715) );
  NOR2_X1 U776 ( .A1(n716), .A2(n715), .ZN(n720) );
  NOR2_X1 U777 ( .A1(n346), .A2(n717), .ZN(n719) );
  NOR2_X1 U778 ( .A1(n720), .A2(n719), .ZN(n729) );
  NAND2_X1 U779 ( .A1(n721), .A2(n635), .ZN(n724) );
  INV_X1 U780 ( .A(KEYINPUT2), .ZN(n722) );
  XNOR2_X1 U781 ( .A(KEYINPUT86), .B(n722), .ZN(n723) );
  NAND2_X1 U782 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U783 ( .A(KEYINPUT85), .B(n725), .ZN(n726) );
  XOR2_X1 U784 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n730) );
  XNOR2_X1 U785 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U786 ( .A(n733), .B(n732), .ZN(n735) );
  INV_X1 U787 ( .A(n734), .ZN(n748) );
  NOR2_X1 U788 ( .A1(n735), .A2(n748), .ZN(n736) );
  XNOR2_X1 U789 ( .A(KEYINPUT56), .B(n736), .ZN(G51) );
  NAND2_X1 U790 ( .A1(n741), .A2(G469), .ZN(n740) );
  XOR2_X1 U791 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n737) );
  NAND2_X1 U792 ( .A1(n741), .A2(G478), .ZN(n744) );
  XOR2_X1 U793 ( .A(n742), .B(KEYINPUT123), .Z(n743) );
  XNOR2_X1 U794 ( .A(n746), .B(n745), .ZN(n747) );
  NOR2_X1 U795 ( .A1(n748), .A2(n747), .ZN(G66) );
  XNOR2_X1 U796 ( .A(n750), .B(n749), .ZN(n753) );
  XNOR2_X1 U797 ( .A(G227), .B(n753), .ZN(n751) );
  NAND2_X1 U798 ( .A1(n751), .A2(G900), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n752), .A2(G953), .ZN(n758) );
  XNOR2_X1 U800 ( .A(n635), .B(n753), .ZN(n754) );
  XNOR2_X1 U801 ( .A(n754), .B(KEYINPUT125), .ZN(n756) );
  NAND2_X1 U802 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U803 ( .A1(n758), .A2(n757), .ZN(G72) );
  XNOR2_X1 U804 ( .A(G122), .B(KEYINPUT126), .ZN(n760) );
  XNOR2_X1 U805 ( .A(n760), .B(n759), .ZN(G24) );
  XOR2_X1 U806 ( .A(G131), .B(n761), .Z(G33) );
  XOR2_X1 U807 ( .A(G134), .B(n762), .Z(G36) );
  XNOR2_X1 U808 ( .A(G137), .B(KEYINPUT127), .ZN(n764) );
  XNOR2_X1 U809 ( .A(n764), .B(n763), .ZN(G39) );
endmodule

