//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n570, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT66), .B1(new_n465), .B2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n465), .A2(G2104), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n466), .A2(new_n469), .A3(new_n461), .A4(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n464), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(new_n470), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n461), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n473), .A2(new_n477), .ZN(G160));
  NAND4_X1  g053(.A1(new_n466), .A2(new_n469), .A3(G2105), .A4(new_n470), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  OR2_X1    g059(.A1(new_n471), .A2(KEYINPUT67), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n471), .A2(KEYINPUT67), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n481), .B(new_n484), .C1(new_n487), .C2(G136), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  NOR3_X1   g065(.A1(new_n465), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n493), .A2(G126), .A3(G2105), .A4(new_n466), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n490), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n490), .B(new_n496), .C1(new_n479), .C2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n474), .A2(new_n470), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR4_X1   g078(.A1(new_n502), .A2(KEYINPUT4), .A3(new_n503), .A4(G2105), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(G2105), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n466), .A2(new_n469), .A3(new_n470), .A4(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n506), .A2(KEYINPUT69), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n508), .B1(new_n506), .B2(KEYINPUT69), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n504), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n489), .B1(new_n501), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n496), .B1(new_n479), .B2(new_n498), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT68), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(new_n499), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n507), .A2(new_n509), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n514), .B(KEYINPUT70), .C1(new_n515), .C2(new_n504), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n511), .A2(new_n516), .ZN(G164));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n521), .B1(new_n522), .B2(G543), .ZN(new_n523));
  NOR3_X1   g098(.A1(new_n519), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n518), .B(new_n520), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT72), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT71), .B1(new_n519), .B2(KEYINPUT5), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n521), .A2(new_n522), .A3(G543), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n527), .A2(new_n528), .B1(KEYINPUT5), .B2(new_n519), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n529), .A2(new_n530), .A3(new_n518), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G88), .ZN(new_n534));
  NAND2_X1  g109(.A1(G75), .A2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n536));
  INV_X1    g111(.A(G62), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n518), .A2(G543), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n538), .A2(G651), .B1(G50), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n534), .A2(new_n540), .ZN(G303));
  INV_X1    g116(.A(G303), .ZN(G166));
  NAND2_X1  g117(.A1(new_n533), .A2(G89), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n529), .A2(KEYINPUT73), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n547), .A2(G63), .A3(G651), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n549));
  NAND3_X1  g124(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n549), .B(new_n550), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(G51), .B2(new_n539), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n543), .A2(new_n548), .A3(new_n552), .ZN(G286));
  INV_X1    g128(.A(G286), .ZN(G168));
  INV_X1    g129(.A(G651), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n547), .A2(G64), .ZN(new_n556));
  NAND2_X1  g131(.A1(G77), .A2(G543), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n539), .A2(G52), .ZN(new_n559));
  INV_X1    g134(.A(G90), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n532), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n558), .A2(new_n561), .ZN(G171));
  AOI22_X1  g137(.A1(new_n533), .A2(G81), .B1(G43), .B2(new_n539), .ZN(new_n563));
  AND3_X1   g138(.A1(new_n545), .A2(G56), .A3(new_n546), .ZN(new_n564));
  AND2_X1   g139(.A1(G68), .A2(G543), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT75), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  AND2_X1   g148(.A1(new_n533), .A2(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n539), .A2(G53), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n575), .A2(KEYINPUT9), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(KEYINPUT9), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n529), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n576), .A2(new_n577), .B1(new_n555), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  NAND3_X1  g157(.A1(new_n526), .A2(G87), .A3(new_n531), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n539), .A2(G49), .ZN(new_n584));
  AOI21_X1  g159(.A(G74), .B1(new_n545), .B2(new_n546), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n555), .ZN(G288));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT76), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n536), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G48), .B2(new_n539), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n526), .A2(G86), .A3(new_n531), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(new_n547), .A2(G60), .ZN(new_n594));
  NAND2_X1  g169(.A1(G72), .A2(G543), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n555), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n539), .A2(G47), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n532), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n533), .A2(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n539), .A2(G54), .ZN(new_n606));
  AND2_X1   g181(.A1(G79), .A2(G543), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(new_n529), .B2(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(G651), .B1(new_n608), .B2(KEYINPUT77), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n610));
  AOI211_X1 g185(.A(new_n610), .B(new_n607), .C1(new_n529), .C2(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n606), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n605), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n602), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n602), .B1(new_n617), .B2(G868), .ZN(G321));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  OR3_X1    g195(.A1(G168), .A2(KEYINPUT79), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(KEYINPUT79), .B1(G168), .B2(new_n620), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n621), .B(new_n622), .C1(G868), .C2(new_n580), .ZN(G297));
  OAI211_X1 g198(.A(new_n621), .B(new_n622), .C1(G868), .C2(new_n580), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n617), .B1(new_n625), .B2(G860), .ZN(G148));
  OR3_X1    g201(.A1(new_n616), .A2(KEYINPUT80), .A3(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(KEYINPUT80), .B1(new_n616), .B2(G559), .ZN(new_n628));
  AND3_X1   g203(.A1(new_n627), .A2(G868), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(new_n620), .B2(new_n567), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g206(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT12), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2100), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n480), .A2(G123), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n461), .A2(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n485), .A2(new_n486), .ZN(new_n639));
  INV_X1    g214(.A(G135), .ZN(new_n640));
  OAI221_X1 g215(.A(new_n636), .B1(new_n637), .B2(new_n638), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n635), .A2(new_n642), .A3(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  INV_X1    g220(.A(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2430), .Z(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT82), .B(KEYINPUT14), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n652), .A2(new_n653), .ZN(new_n658));
  AND3_X1   g233(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n657), .B1(new_n654), .B2(new_n658), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  OAI21_X1  g237(.A(G14), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n653), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n652), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n657), .ZN(new_n666));
  INV_X1    g241(.A(new_n662), .ZN(new_n667));
  OAI21_X1  g242(.A(KEYINPUT83), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT83), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n661), .A2(new_n669), .A3(new_n662), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n663), .B1(new_n668), .B2(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n672), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(KEYINPUT17), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n672), .A2(new_n673), .ZN(new_n679));
  OAI221_X1 g254(.A(new_n674), .B1(new_n673), .B2(new_n677), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n674), .A2(new_n676), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT18), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT84), .B(G2096), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT87), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1956), .B(G2474), .Z(new_n692));
  XOR2_X1   g267(.A(G1961), .B(G1966), .Z(new_n693));
  AND2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT20), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n692), .A2(new_n693), .ZN(new_n698));
  OR3_X1    g273(.A1(new_n691), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n691), .A2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n697), .A2(new_n701), .A3(KEYINPUT85), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n703));
  OAI21_X1  g278(.A(KEYINPUT85), .B1(new_n697), .B2(new_n701), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n703), .B1(new_n702), .B2(new_n704), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n688), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n707), .ZN(new_n709));
  INV_X1    g284(.A(new_n688), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n709), .A2(new_n710), .A3(new_n705), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT88), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n714), .B(new_n715), .Z(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n708), .A2(new_n711), .A3(new_n716), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(G229));
  NAND2_X1  g296(.A1(G166), .A2(G16), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G16), .B2(G22), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT93), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT92), .B(G1971), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n723), .B(KEYINPUT93), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(new_n726), .ZN(new_n730));
  MUX2_X1   g305(.A(G23), .B(G288), .S(G16), .Z(new_n731));
  XOR2_X1   g306(.A(KEYINPUT33), .B(G1976), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(G6), .A2(G16), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(G305), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT32), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n733), .B1(G1981), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G1981), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n728), .A2(new_n730), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT34), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(KEYINPUT34), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n487), .A2(G131), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(KEYINPUT89), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(KEYINPUT89), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n749));
  INV_X1    g324(.A(G107), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G2105), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT90), .ZN(new_n752));
  INV_X1    g327(.A(G119), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(new_n479), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n748), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G29), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G25), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT35), .B(G1991), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT91), .Z(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n759), .A2(new_n762), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n600), .A2(new_n735), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n735), .B2(G24), .ZN(new_n766));
  INV_X1    g341(.A(G1986), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NOR4_X1   g344(.A1(new_n763), .A2(new_n764), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n743), .A2(new_n744), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT36), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n735), .A2(G5), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G171), .B2(new_n735), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(G1961), .Z(new_n775));
  INV_X1    g350(.A(G29), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(G32), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n480), .A2(G129), .ZN(new_n778));
  NAND3_X1  g353(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT26), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G105), .B2(new_n463), .ZN(new_n781));
  INV_X1    g356(.A(G141), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n778), .B(new_n781), .C1(new_n639), .C2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT96), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n777), .B1(new_n784), .B2(new_n776), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT27), .B(G1996), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G27), .A2(G29), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G164), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT98), .B(G2078), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n775), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n735), .A2(G21), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G168), .B2(new_n735), .ZN(new_n794));
  INV_X1    g369(.A(G2072), .ZN(new_n795));
  NOR2_X1   g370(.A1(G29), .A2(G33), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT95), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n487), .A2(G139), .ZN(new_n798));
  NAND2_X1  g373(.A1(G115), .A2(G2104), .ZN(new_n799));
  INV_X1    g374(.A(G127), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n502), .B2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT25), .ZN(new_n802));
  NAND2_X1  g377(.A1(G103), .A2(G2104), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G2105), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n801), .A2(G2105), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n798), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n797), .B1(new_n807), .B2(new_n776), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n794), .A2(G1966), .B1(new_n795), .B2(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n795), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G16), .A2(G19), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n567), .B2(G16), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(G1341), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT24), .ZN(new_n815));
  INV_X1    g390(.A(G34), .ZN(new_n816));
  AOI21_X1  g391(.A(G29), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n815), .B2(new_n816), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G160), .B2(new_n776), .ZN(new_n819));
  INV_X1    g394(.A(G2084), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n794), .B2(G1966), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n811), .A2(new_n814), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n735), .A2(G20), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT23), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n580), .B2(new_n735), .ZN(new_n827));
  INV_X1    g402(.A(G1956), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT30), .B(G28), .ZN(new_n830));
  OR2_X1    g405(.A1(KEYINPUT31), .A2(G11), .ZN(new_n831));
  NAND2_X1  g406(.A1(KEYINPUT31), .A2(G11), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n830), .A2(new_n776), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n641), .B2(new_n776), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT97), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n813), .A2(G1341), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n776), .A2(G26), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT28), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n487), .A2(G140), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n840));
  INV_X1    g415(.A(G116), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n840), .B1(new_n841), .B2(G2105), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n480), .B2(G128), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n838), .B1(new_n844), .B2(G29), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G2067), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n829), .A2(new_n835), .A3(new_n836), .A4(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n824), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(G4), .A2(G16), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT94), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n616), .B2(new_n735), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(G1348), .Z(new_n852));
  NOR2_X1   g427(.A1(G29), .A2(G35), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(G162), .B2(G29), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT29), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G2090), .ZN(new_n856));
  NOR4_X1   g431(.A1(new_n792), .A2(new_n848), .A3(new_n852), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n772), .A2(new_n857), .ZN(G150));
  INV_X1    g433(.A(G150), .ZN(G311));
  NOR2_X1   g434(.A1(new_n616), .A2(new_n625), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n547), .A2(G67), .ZN(new_n862));
  NAND2_X1  g437(.A1(G80), .A2(G543), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n555), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n539), .A2(G55), .ZN(new_n865));
  INV_X1    g440(.A(G93), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n532), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n563), .A2(new_n566), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n861), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n872));
  AOI21_X1  g447(.A(G860), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n872), .B2(new_n871), .ZN(new_n874));
  OAI21_X1  g449(.A(G860), .B1(new_n864), .B2(new_n867), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT37), .Z(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(G145));
  NAND2_X1  g452(.A1(new_n756), .A2(new_n633), .ZN(new_n878));
  INV_X1    g453(.A(new_n633), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n748), .A2(new_n879), .A3(new_n755), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT96), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n783), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n844), .ZN(new_n884));
  INV_X1    g459(.A(new_n844), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n784), .A2(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(G106), .A2(G2105), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n887), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n888));
  INV_X1    g463(.A(G130), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n479), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(new_n487), .B2(G142), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n884), .A2(new_n886), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n892), .B1(new_n884), .B2(new_n886), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n881), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n510), .A2(new_n512), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n784), .A2(new_n885), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n883), .A2(new_n844), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n891), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n879), .B1(new_n748), .B2(new_n755), .ZN(new_n901));
  AOI211_X1 g476(.A(new_n633), .B(new_n754), .C1(new_n746), .C2(new_n747), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n884), .A2(new_n886), .A3(new_n892), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n895), .A2(new_n897), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n897), .B1(new_n895), .B2(new_n905), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n807), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n900), .A2(new_n903), .A3(new_n904), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n903), .B1(new_n900), .B2(new_n904), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n896), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n807), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n895), .A2(new_n905), .A3(new_n897), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n641), .B(G160), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(G162), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n908), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT99), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n908), .A2(new_n914), .A3(KEYINPUT99), .A4(new_n916), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n916), .B1(new_n908), .B2(new_n914), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(G37), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n921), .A2(KEYINPUT40), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT40), .B1(new_n921), .B2(new_n923), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(G395));
  NAND2_X1  g501(.A1(new_n627), .A2(new_n628), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(new_n870), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n616), .A2(G299), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n605), .B(new_n580), .C1(new_n615), .C2(new_n614), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(new_n931), .B2(KEYINPUT41), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT41), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n929), .A2(KEYINPUT100), .A3(new_n935), .A4(new_n930), .ZN(new_n936));
  XOR2_X1   g511(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n931), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n928), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n600), .B(G305), .ZN(new_n942));
  XOR2_X1   g517(.A(G303), .B(G288), .Z(new_n943));
  XOR2_X1   g518(.A(new_n942), .B(new_n943), .Z(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(KEYINPUT42), .Z(new_n945));
  AND3_X1   g520(.A1(new_n932), .A2(new_n941), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(new_n932), .B2(new_n941), .ZN(new_n947));
  OAI21_X1  g522(.A(G868), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(G868), .B2(new_n868), .ZN(G295));
  OAI21_X1  g524(.A(new_n948), .B1(G868), .B2(new_n868), .ZN(G331));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n951));
  XNOR2_X1  g526(.A(G171), .B(G286), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n870), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n870), .A2(new_n952), .A3(KEYINPUT104), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n868), .B(new_n567), .ZN(new_n957));
  XNOR2_X1  g532(.A(G171), .B(G168), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n957), .A2(new_n958), .A3(KEYINPUT103), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT103), .B1(new_n957), .B2(new_n958), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n955), .B(new_n956), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n957), .A2(new_n958), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n953), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n937), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n931), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n963), .A2(KEYINPUT41), .A3(new_n931), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n944), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G37), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n963), .A2(new_n931), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n940), .B2(new_n961), .ZN(new_n970));
  INV_X1    g545(.A(new_n944), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n967), .A2(new_n968), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n970), .A2(new_n971), .ZN(new_n975));
  XOR2_X1   g550(.A(KEYINPUT102), .B(KEYINPUT43), .Z(new_n976));
  NAND4_X1  g551(.A1(new_n975), .A2(new_n968), .A3(new_n972), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n951), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n976), .ZN(new_n979));
  INV_X1    g554(.A(new_n972), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n967), .A2(new_n968), .A3(new_n972), .A4(new_n976), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n982), .A2(new_n951), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n978), .A2(new_n984), .ZN(G397));
  INV_X1    g560(.A(G1384), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n510), .B2(new_n512), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(G40), .B(new_n464), .C1(new_n471), .C2(new_n472), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(new_n477), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1996), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT106), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n784), .A2(new_n994), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n844), .B(G2067), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n996), .A2(new_n784), .B1(new_n999), .B2(new_n993), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n757), .A2(new_n762), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n756), .A2(new_n761), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n993), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n600), .A2(new_n767), .ZN(new_n1005));
  XOR2_X1   g580(.A(new_n1005), .B(KEYINPUT105), .Z(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n767), .B2(new_n600), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1004), .B1(new_n993), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(G303), .A2(G8), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT55), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1013), .B(new_n986), .C1(new_n510), .C2(new_n512), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n511), .A2(new_n986), .A3(new_n516), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(KEYINPUT50), .ZN(new_n1017));
  INV_X1    g592(.A(G2090), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n991), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n991), .B1(new_n987), .B2(new_n988), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(new_n1016), .B2(new_n988), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(G1971), .ZN(new_n1022));
  OAI211_X1 g597(.A(G8), .B(new_n1012), .C1(new_n1019), .C2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n591), .A2(new_n740), .A3(new_n592), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT110), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT110), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n591), .A2(new_n592), .A3(new_n1026), .A4(new_n740), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n740), .B1(new_n591), .B2(new_n592), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(KEYINPUT49), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n986), .B(new_n991), .C1(new_n510), .C2(new_n512), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT107), .B(G8), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1029), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1033), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1034), .A2(new_n1041), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n583), .A2(new_n584), .ZN(new_n1043));
  OAI21_X1  g618(.A(G651), .B1(new_n547), .B2(G74), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1043), .A2(new_n1044), .A3(KEYINPUT108), .A4(G1976), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n1046));
  INV_X1    g621(.A(G1976), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(G288), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT52), .B1(new_n1049), .B2(new_n1038), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1047), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1051), .A2(new_n1048), .A3(new_n1052), .A4(new_n1045), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT109), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1042), .B(new_n1050), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1023), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1042), .A2(new_n1047), .A3(new_n1044), .A4(new_n1043), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT112), .B1(new_n1059), .B2(new_n1028), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(new_n1038), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(KEYINPUT112), .A3(new_n1028), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1058), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT56), .B(G2072), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n511), .A2(new_n1013), .A3(new_n986), .A4(new_n516), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n992), .B1(new_n987), .B2(KEYINPUT50), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1021), .A2(new_n1065), .B1(new_n1068), .B2(new_n828), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n580), .B(KEYINPUT57), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1064), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1070), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1065), .ZN(new_n1073));
  AOI211_X1 g648(.A(new_n1073), .B(new_n1020), .C1(new_n1016), .C2(new_n988), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1956), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1072), .B(KEYINPUT117), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1348), .B1(new_n1017), .B2(new_n991), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1035), .B(KEYINPUT116), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(G2067), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n617), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1071), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1068), .A2(new_n828), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1016), .A2(new_n988), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1020), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1082), .B(new_n1070), .C1(new_n1085), .C2(new_n1073), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT115), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1069), .A2(new_n1088), .A3(new_n1070), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1081), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT118), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1081), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1082), .B1(new_n1085), .B2(new_n1073), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(new_n1072), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1069), .A2(KEYINPUT119), .A3(new_n1070), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT61), .B1(new_n1099), .B2(new_n1090), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT61), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1071), .A2(new_n1102), .A3(new_n1076), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1079), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n992), .B(new_n1015), .C1(new_n1016), .C2(KEYINPUT50), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1106), .B(KEYINPUT60), .C1(new_n1107), .C2(G1348), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1108), .A3(new_n617), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(KEYINPUT60), .A3(new_n616), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT58), .B(G1341), .Z(new_n1112));
  AOI22_X1  g687(.A1(new_n1021), .A2(new_n994), .B1(new_n1078), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT59), .B1(new_n1113), .B2(new_n869), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n1115));
  AOI211_X1 g690(.A(G1996), .B(new_n1020), .C1(new_n1016), .C2(new_n988), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1078), .A2(new_n1112), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1115), .B(new_n567), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1103), .A2(new_n1109), .A3(new_n1111), .A4(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1092), .B(new_n1094), .C1(new_n1100), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1051), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1050), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1068), .A2(G2090), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1037), .B1(new_n1022), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n1011), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1130), .A3(new_n1023), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n1133));
  INV_X1    g708(.A(G2078), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1021), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1017), .A2(new_n991), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT121), .B(G1961), .Z(new_n1137));
  AOI22_X1  g712(.A1(new_n1133), .A2(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n475), .A2(new_n476), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n1140));
  OAI21_X1  g715(.A(G2105), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n1140), .B2(new_n1139), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1142), .A2(KEYINPUT123), .A3(new_n990), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT124), .B(G2078), .Z(new_n1144));
  NOR3_X1   g719(.A1(new_n1143), .A2(new_n1133), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n987), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT45), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT123), .B1(new_n1142), .B2(new_n990), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1145), .A2(new_n1147), .A3(new_n989), .A4(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1138), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1132), .B1(new_n1150), .B2(G171), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n511), .A2(KEYINPUT45), .A3(new_n986), .A4(new_n516), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n992), .B1(new_n987), .B2(new_n988), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1152), .A2(KEYINPUT53), .A3(new_n1134), .A4(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1138), .A2(G301), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1131), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1017), .A2(new_n820), .A3(new_n991), .ZN(new_n1157));
  AOI21_X1  g732(.A(G1966), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n991), .A2(new_n820), .ZN(new_n1162));
  AOI211_X1 g737(.A(new_n1015), .B(new_n1162), .C1(new_n1016), .C2(KEYINPUT50), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT120), .B1(new_n1163), .B2(new_n1158), .ZN(new_n1164));
  NOR2_X1   g739(.A1(G168), .A2(new_n1036), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1161), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT51), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1161), .A2(new_n1164), .A3(G8), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1165), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1171));
  AOI211_X1 g746(.A(KEYINPUT51), .B(new_n1165), .C1(new_n1171), .C2(new_n1037), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1166), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1135), .A2(new_n1133), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1174), .A2(new_n1175), .A3(G301), .A4(new_n1149), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT125), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1138), .A2(new_n1178), .A3(G301), .A4(new_n1149), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1174), .A2(new_n1175), .A3(new_n1154), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(G171), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1177), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1156), .B(new_n1173), .C1(KEYINPUT54), .C2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1063), .B1(new_n1122), .B2(new_n1183), .ZN(new_n1184));
  AOI211_X1 g759(.A(G286), .B(new_n1036), .C1(new_n1157), .C2(new_n1159), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(KEYINPUT113), .B1(new_n1131), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(G8), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n1021), .A2(G1971), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1017), .A2(new_n1018), .A3(new_n991), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1057), .B1(new_n1012), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT113), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1192), .A2(new_n1193), .A3(new_n1130), .A4(new_n1185), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT63), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1187), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1185), .B(KEYINPUT63), .C1(new_n1012), .C2(new_n1191), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1127), .A2(new_n1023), .ZN(new_n1198));
  OAI21_X1  g773(.A(KEYINPUT114), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OR3_X1    g774(.A1(new_n1197), .A2(new_n1198), .A3(KEYINPUT114), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1196), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1173), .A2(KEYINPUT62), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n1203));
  OAI211_X1 g778(.A(new_n1203), .B(new_n1166), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1131), .A2(new_n1181), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1201), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1009), .B1(new_n1184), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1209));
  OR2_X1    g784(.A1(new_n844), .A2(G2067), .ZN(new_n1210));
  AOI211_X1 g785(.A(new_n992), .B(new_n989), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT46), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n996), .B(new_n1212), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n993), .B1(new_n998), .B2(new_n883), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT47), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n1215), .B(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1004), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1006), .A2(new_n993), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1219), .B(KEYINPUT48), .ZN(new_n1220));
  AOI211_X1 g795(.A(new_n1211), .B(new_n1217), .C1(new_n1218), .C2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1208), .A2(new_n1221), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g797(.A(G14), .ZN(new_n1224));
  AOI21_X1  g798(.A(new_n1224), .B1(new_n666), .B2(new_n667), .ZN(new_n1225));
  AOI21_X1  g799(.A(new_n669), .B1(new_n661), .B2(new_n662), .ZN(new_n1226));
  NOR4_X1   g800(.A1(new_n659), .A2(new_n660), .A3(KEYINPUT83), .A4(new_n667), .ZN(new_n1227));
  OAI21_X1  g801(.A(new_n1225), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g802(.A1(G227), .A2(new_n459), .ZN(new_n1229));
  NAND2_X1  g803(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n1231));
  AOI22_X1  g805(.A1(new_n1230), .A2(new_n1231), .B1(new_n719), .B2(new_n718), .ZN(new_n1232));
  NAND3_X1  g806(.A1(new_n1228), .A2(KEYINPUT126), .A3(new_n1229), .ZN(new_n1233));
  AOI21_X1  g807(.A(KEYINPUT127), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  OR2_X1    g808(.A1(G227), .A2(new_n459), .ZN(new_n1235));
  OAI21_X1  g809(.A(new_n1231), .B1(G401), .B2(new_n1235), .ZN(new_n1236));
  AND4_X1   g810(.A1(KEYINPUT127), .A2(new_n1236), .A3(new_n720), .A4(new_n1233), .ZN(new_n1237));
  NOR2_X1   g811(.A1(new_n1234), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g812(.A(new_n1238), .B1(new_n921), .B2(new_n923), .ZN(new_n1239));
  NAND2_X1  g813(.A1(new_n982), .A2(new_n983), .ZN(new_n1240));
  AND2_X1   g814(.A1(new_n1239), .A2(new_n1240), .ZN(G308));
  NAND2_X1  g815(.A1(new_n1239), .A2(new_n1240), .ZN(G225));
endmodule


