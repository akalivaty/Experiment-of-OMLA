

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762;

  NOR2_X1 U377 ( .A1(n594), .A2(n601), .ZN(n673) );
  XNOR2_X1 U378 ( .A(n631), .B(n630), .ZN(n642) );
  AND2_X4 U379 ( .A1(n402), .A2(n401), .ZN(n724) );
  AND2_X2 U380 ( .A1(n451), .A2(n363), .ZN(n456) );
  XNOR2_X2 U381 ( .A(n746), .B(n513), .ZN(n571) );
  NOR2_X2 U382 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X2 U383 ( .A1(n435), .A2(n456), .ZN(n650) );
  NOR2_X1 U384 ( .A1(n695), .A2(n597), .ZN(n598) );
  NOR2_X1 U385 ( .A1(G953), .A2(G237), .ZN(n531) );
  INV_X1 U386 ( .A(n710), .ZN(n354) );
  AND2_X1 U387 ( .A1(n638), .A2(n455), .ZN(n450) );
  XNOR2_X1 U388 ( .A(n598), .B(n392), .ZN(n757) );
  NOR2_X1 U389 ( .A1(n715), .A2(G902), .ZN(n573) );
  XNOR2_X1 U390 ( .A(n557), .B(n556), .ZN(n558) );
  INV_X1 U391 ( .A(KEYINPUT87), .ZN(n546) );
  NAND2_X1 U392 ( .A1(n395), .A2(n393), .ZN(n710) );
  XNOR2_X1 U393 ( .A(n626), .B(n625), .ZN(n759) );
  NAND2_X1 U394 ( .A1(n406), .A2(n404), .ZN(n637) );
  XNOR2_X1 U395 ( .A(n441), .B(n440), .ZN(n627) );
  AND2_X1 U396 ( .A1(n620), .A2(n687), .ZN(n441) );
  NOR2_X1 U397 ( .A1(n597), .A2(n618), .ZN(n668) );
  AND2_X1 U398 ( .A1(n646), .A2(n434), .ZN(n620) );
  XNOR2_X1 U399 ( .A(n436), .B(n596), .ZN(n695) );
  OR2_X1 U400 ( .A1(n696), .A2(n701), .ZN(n436) );
  XNOR2_X1 U401 ( .A(n579), .B(KEYINPUT19), .ZN(n618) );
  OR2_X1 U402 ( .A1(n629), .A2(n684), .ZN(n631) );
  XNOR2_X1 U403 ( .A(n693), .B(KEYINPUT6), .ZN(n640) );
  XNOR2_X1 U404 ( .A(n587), .B(KEYINPUT67), .ZN(n684) );
  AND2_X1 U405 ( .A1(n586), .A2(n687), .ZN(n587) );
  XNOR2_X1 U406 ( .A(n416), .B(n415), .ZN(n643) );
  XNOR2_X1 U407 ( .A(n547), .B(n546), .ZN(n549) );
  INV_X2 U408 ( .A(G953), .ZN(n750) );
  INV_X1 U409 ( .A(G143), .ZN(n414) );
  NOR2_X2 U410 ( .A1(n734), .A2(n749), .ZN(n681) );
  INV_X1 U411 ( .A(KEYINPUT33), .ZN(n444) );
  INV_X1 U412 ( .A(G469), .ZN(n373) );
  XNOR2_X1 U413 ( .A(n650), .B(KEYINPUT45), .ZN(n734) );
  NAND2_X1 U414 ( .A1(n762), .A2(n757), .ZN(n391) );
  XNOR2_X1 U415 ( .A(KEYINPUT15), .B(G902), .ZN(n651) );
  INV_X1 U416 ( .A(G472), .ZN(n415) );
  OR2_X1 U417 ( .A1(n654), .A2(G902), .ZN(n416) );
  AND2_X1 U418 ( .A1(n683), .A2(n359), .ZN(n395) );
  XNOR2_X1 U419 ( .A(n681), .B(n483), .ZN(n394) );
  INV_X1 U420 ( .A(KEYINPUT1), .ZN(n371) );
  INV_X1 U421 ( .A(KEYINPUT22), .ZN(n440) );
  NOR2_X1 U422 ( .A1(n374), .A2(n695), .ZN(n706) );
  XNOR2_X1 U423 ( .A(n375), .B(KEYINPUT51), .ZN(n374) );
  OR2_X1 U424 ( .A1(n694), .A2(n376), .ZN(n375) );
  NAND2_X1 U425 ( .A1(G234), .A2(G237), .ZN(n496) );
  XNOR2_X1 U426 ( .A(G116), .B(G137), .ZN(n519) );
  AND2_X1 U427 ( .A1(n600), .A2(n389), .ZN(n388) );
  NOR2_X1 U428 ( .A1(n599), .A2(n605), .ZN(n389) );
  XNOR2_X1 U429 ( .A(n517), .B(n518), .ZN(n561) );
  XNOR2_X1 U430 ( .A(n514), .B(G113), .ZN(n518) );
  INV_X1 U431 ( .A(KEYINPUT86), .ZN(n515) );
  NOR2_X1 U432 ( .A1(n458), .A2(KEYINPUT70), .ZN(n453) );
  XNOR2_X1 U433 ( .A(n569), .B(n568), .ZN(n570) );
  INV_X1 U434 ( .A(KEYINPUT89), .ZN(n568) );
  XNOR2_X1 U435 ( .A(n567), .B(KEYINPUT74), .ZN(n446) );
  INV_X1 U436 ( .A(G137), .ZN(n448) );
  XNOR2_X1 U437 ( .A(n378), .B(n377), .ZN(n709) );
  INV_X1 U438 ( .A(KEYINPUT116), .ZN(n377) );
  NAND2_X1 U439 ( .A1(n380), .A2(n379), .ZN(n378) );
  INV_X1 U440 ( .A(n708), .ZN(n379) );
  NAND2_X1 U441 ( .A1(n400), .A2(n398), .ZN(n576) );
  NOR2_X1 U442 ( .A1(n399), .A2(n590), .ZN(n398) );
  INV_X1 U443 ( .A(n687), .ZN(n399) );
  OR2_X1 U444 ( .A1(n576), .A2(n643), .ZN(n397) );
  XOR2_X1 U445 ( .A(n545), .B(n544), .Z(n595) );
  AND2_X1 U446 ( .A1(n484), .A2(n670), .ZN(n606) );
  NOR2_X1 U447 ( .A1(n640), .A2(n417), .ZN(n484) );
  NAND2_X1 U448 ( .A1(n418), .A2(n698), .ZN(n417) );
  INV_X1 U449 ( .A(n576), .ZN(n418) );
  NOR2_X1 U450 ( .A1(n634), .A2(n364), .ZN(n410) );
  AND2_X1 U451 ( .A1(n407), .A2(n408), .ZN(n406) );
  AND2_X1 U452 ( .A1(n409), .A2(n430), .ZN(n408) );
  AND2_X1 U453 ( .A1(n622), .A2(n412), .ZN(n623) );
  AND2_X1 U454 ( .A1(n621), .A2(n400), .ZN(n412) );
  XNOR2_X1 U455 ( .A(n428), .B(n427), .ZN(n589) );
  NOR2_X1 U456 ( .A1(n602), .A2(n595), .ZN(n592) );
  NOR2_X1 U457 ( .A1(n628), .A2(n627), .ZN(n639) );
  XNOR2_X1 U458 ( .A(n488), .B(n485), .ZN(n725) );
  XNOR2_X1 U459 ( .A(n527), .B(n486), .ZN(n485) );
  XNOR2_X1 U460 ( .A(n524), .B(n525), .ZN(n488) );
  XNOR2_X1 U461 ( .A(n528), .B(n487), .ZN(n486) );
  NAND2_X1 U462 ( .A1(n403), .A2(n365), .ZN(n402) );
  NOR2_X1 U463 ( .A1(n463), .A2(n470), .ZN(n462) );
  INV_X1 U464 ( .A(n466), .ZN(n463) );
  AND2_X1 U465 ( .A1(n459), .A2(n470), .ZN(n383) );
  NAND2_X1 U466 ( .A1(n354), .A2(n466), .ZN(n384) );
  NAND2_X1 U467 ( .A1(n354), .A2(n355), .ZN(n467) );
  INV_X1 U468 ( .A(KEYINPUT46), .ZN(n432) );
  XNOR2_X1 U469 ( .A(G119), .B(KEYINPUT69), .ZN(n514) );
  XNOR2_X1 U470 ( .A(KEYINPUT68), .B(KEYINPUT3), .ZN(n516) );
  XNOR2_X1 U471 ( .A(n707), .B(n381), .ZN(n380) );
  XNOR2_X1 U472 ( .A(KEYINPUT115), .B(KEYINPUT52), .ZN(n381) );
  INV_X1 U473 ( .A(KEYINPUT48), .ZN(n425) );
  XOR2_X1 U474 ( .A(KEYINPUT98), .B(KEYINPUT96), .Z(n537) );
  XNOR2_X1 U475 ( .A(G143), .B(G140), .ZN(n536) );
  XNOR2_X1 U476 ( .A(n532), .B(n442), .ZN(n535) );
  XNOR2_X1 U477 ( .A(n533), .B(n443), .ZN(n442) );
  INV_X1 U478 ( .A(G131), .ZN(n443) );
  XNOR2_X1 U479 ( .A(KEYINPUT11), .B(KEYINPUT95), .ZN(n538) );
  XOR2_X1 U480 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n539) );
  XOR2_X1 U481 ( .A(G125), .B(G146), .Z(n551) );
  INV_X1 U482 ( .A(KEYINPUT77), .ZN(n483) );
  INV_X1 U483 ( .A(n701), .ZN(n434) );
  NOR2_X1 U484 ( .A1(n643), .A2(n588), .ZN(n428) );
  INV_X1 U485 ( .A(KEYINPUT30), .ZN(n427) );
  OR2_X1 U486 ( .A1(G902), .A2(G237), .ZN(n563) );
  AND2_X1 U487 ( .A1(G953), .A2(G902), .ZN(n497) );
  XNOR2_X1 U488 ( .A(n411), .B(n561), .ZN(n522) );
  XNOR2_X1 U489 ( .A(n358), .B(n521), .ZN(n411) );
  XOR2_X1 U490 ( .A(G110), .B(KEYINPUT16), .Z(n559) );
  XNOR2_X1 U491 ( .A(n477), .B(KEYINPUT24), .ZN(n476) );
  INV_X1 U492 ( .A(KEYINPUT23), .ZN(n477) );
  XNOR2_X1 U493 ( .A(n482), .B(n481), .ZN(n523) );
  INV_X1 U494 ( .A(KEYINPUT8), .ZN(n481) );
  NAND2_X1 U495 ( .A1(n750), .A2(G234), .ZN(n482) );
  INV_X1 U496 ( .A(G134), .ZN(n487) );
  NAND2_X1 U497 ( .A1(n681), .A2(n652), .ZN(n403) );
  XNOR2_X1 U498 ( .A(n447), .B(n413), .ZN(n572) );
  XNOR2_X1 U499 ( .A(n446), .B(G110), .ZN(n413) );
  XNOR2_X1 U500 ( .A(n570), .B(n357), .ZN(n447) );
  NOR2_X1 U501 ( .A1(G953), .A2(n360), .ZN(n466) );
  INV_X1 U502 ( .A(KEYINPUT53), .ZN(n470) );
  NOR2_X1 U503 ( .A1(n608), .A2(n588), .ZN(n579) );
  XNOR2_X1 U504 ( .A(n397), .B(n396), .ZN(n578) );
  INV_X1 U505 ( .A(KEYINPUT28), .ZN(n396) );
  NOR2_X1 U506 ( .A1(n684), .A2(n370), .ZN(n647) );
  XNOR2_X1 U507 ( .A(n593), .B(n489), .ZN(n762) );
  XNOR2_X1 U508 ( .A(KEYINPUT81), .B(KEYINPUT36), .ZN(n431) );
  INV_X1 U509 ( .A(KEYINPUT35), .ZN(n636) );
  NAND2_X1 U510 ( .A1(n405), .A2(n410), .ZN(n404) );
  XNOR2_X1 U511 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n625) );
  NOR2_X1 U512 ( .A1(n627), .A2(n624), .ZN(n626) );
  XNOR2_X1 U513 ( .A(n645), .B(KEYINPUT31), .ZN(n674) );
  NOR2_X1 U514 ( .A1(n693), .A2(n686), .ZN(n429) );
  XNOR2_X1 U515 ( .A(n592), .B(KEYINPUT102), .ZN(n670) );
  AND2_X1 U516 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U517 ( .A(n725), .B(KEYINPUT119), .ZN(n479) );
  INV_X1 U518 ( .A(KEYINPUT60), .ZN(n419) );
  INV_X1 U519 ( .A(KEYINPUT56), .ZN(n421) );
  AND2_X1 U520 ( .A1(n468), .A2(n462), .ZN(n461) );
  INV_X1 U521 ( .A(n643), .ZN(n693) );
  NOR2_X1 U522 ( .A1(n709), .A2(n469), .ZN(n355) );
  AND2_X1 U523 ( .A1(n639), .A2(n429), .ZN(n356) );
  XOR2_X1 U524 ( .A(n448), .B(G140), .Z(n357) );
  XOR2_X1 U525 ( .A(n520), .B(n519), .Z(n358) );
  XNOR2_X1 U526 ( .A(n608), .B(KEYINPUT38), .ZN(n699) );
  OR2_X1 U527 ( .A1(n695), .A2(n680), .ZN(n359) );
  AND2_X1 U528 ( .A1(n709), .A2(n469), .ZN(n360) );
  XOR2_X1 U529 ( .A(G131), .B(G134), .Z(n361) );
  BUF_X1 U530 ( .A(n586), .Z(n686) );
  INV_X1 U531 ( .A(n686), .ZN(n400) );
  AND2_X1 U532 ( .A1(n355), .A2(n470), .ZN(n362) );
  OR2_X1 U533 ( .A1(n457), .A2(KEYINPUT44), .ZN(n363) );
  XOR2_X1 U534 ( .A(KEYINPUT71), .B(KEYINPUT34), .Z(n364) );
  XOR2_X1 U535 ( .A(n491), .B(KEYINPUT65), .Z(n365) );
  XNOR2_X1 U536 ( .A(n532), .B(n357), .ZN(n745) );
  XOR2_X1 U537 ( .A(n654), .B(KEYINPUT62), .Z(n366) );
  INV_X1 U538 ( .A(KEYINPUT70), .ZN(n457) );
  XNOR2_X1 U539 ( .A(n713), .B(n712), .ZN(n367) );
  XOR2_X1 U540 ( .A(n722), .B(n721), .Z(n368) );
  NOR2_X1 U541 ( .A1(G952), .A2(n750), .ZN(n729) );
  INV_X1 U542 ( .A(n729), .ZN(n437) );
  XOR2_X1 U543 ( .A(KEYINPUT63), .B(KEYINPUT85), .Z(n369) );
  INV_X1 U544 ( .A(KEYINPUT117), .ZN(n469) );
  XNOR2_X2 U545 ( .A(n591), .B(KEYINPUT39), .ZN(n612) );
  NAND2_X1 U546 ( .A1(n394), .A2(n653), .ZN(n393) );
  INV_X1 U547 ( .A(n372), .ZN(n370) );
  XNOR2_X2 U548 ( .A(n372), .B(n371), .ZN(n629) );
  XNOR2_X1 U549 ( .A(n372), .B(KEYINPUT106), .ZN(n577) );
  XNOR2_X2 U550 ( .A(n573), .B(n373), .ZN(n372) );
  XNOR2_X2 U551 ( .A(n554), .B(n361), .ZN(n746) );
  XNOR2_X2 U552 ( .A(n526), .B(KEYINPUT4), .ZN(n554) );
  NOR2_X1 U553 ( .A1(n692), .A2(n693), .ZN(n376) );
  XNOR2_X1 U554 ( .A(n644), .B(KEYINPUT94), .ZN(n694) );
  AND2_X1 U555 ( .A1(n465), .A2(n382), .ZN(n464) );
  NAND2_X1 U556 ( .A1(n384), .A2(n383), .ZN(n382) );
  XNOR2_X1 U557 ( .A(n385), .B(n745), .ZN(n727) );
  XNOR2_X1 U558 ( .A(n386), .B(n507), .ZN(n385) );
  XNOR2_X1 U559 ( .A(n387), .B(n506), .ZN(n386) );
  XNOR2_X1 U560 ( .A(n476), .B(n505), .ZN(n387) );
  NAND2_X1 U561 ( .A1(n390), .A2(n388), .ZN(n426) );
  XNOR2_X1 U562 ( .A(n391), .B(n432), .ZN(n390) );
  INV_X1 U563 ( .A(KEYINPUT42), .ZN(n392) );
  NAND2_X1 U564 ( .A1(n681), .A2(KEYINPUT2), .ZN(n401) );
  INV_X1 U565 ( .A(n680), .ZN(n405) );
  NAND2_X1 U566 ( .A1(n680), .A2(n364), .ZN(n407) );
  XNOR2_X2 U567 ( .A(n445), .B(n444), .ZN(n680) );
  NAND2_X1 U568 ( .A1(n634), .A2(n364), .ZN(n409) );
  INV_X1 U569 ( .A(n635), .ZN(n430) );
  XNOR2_X1 U570 ( .A(n571), .B(n572), .ZN(n715) );
  XNOR2_X2 U571 ( .A(n414), .B(G128), .ZN(n526) );
  NAND2_X1 U572 ( .A1(n449), .A2(n452), .ZN(n435) );
  XNOR2_X1 U573 ( .A(n426), .B(n425), .ZN(n475) );
  XNOR2_X1 U574 ( .A(n566), .B(n431), .ZN(n574) );
  XNOR2_X1 U575 ( .A(n420), .B(n419), .ZN(G60) );
  NAND2_X1 U576 ( .A1(n424), .A2(n437), .ZN(n420) );
  XNOR2_X1 U577 ( .A(n422), .B(n421), .ZN(G51) );
  NAND2_X1 U578 ( .A1(n438), .A2(n437), .ZN(n422) );
  XNOR2_X1 U579 ( .A(n423), .B(n369), .ZN(G57) );
  NAND2_X1 U580 ( .A1(n433), .A2(n437), .ZN(n423) );
  NOR2_X2 U581 ( .A1(n759), .A2(n356), .ZN(n638) );
  XNOR2_X1 U582 ( .A(n723), .B(n368), .ZN(n424) );
  NAND2_X1 U583 ( .A1(n490), .A2(n657), .ZN(n454) );
  INV_X1 U584 ( .A(n604), .ZN(n471) );
  NAND2_X1 U585 ( .A1(n472), .A2(n474), .ZN(n604) );
  XNOR2_X1 U586 ( .A(n512), .B(n511), .ZN(n586) );
  XNOR2_X1 U587 ( .A(n655), .B(n366), .ZN(n433) );
  NOR2_X1 U588 ( .A1(n454), .A2(n453), .ZN(n452) );
  NOR2_X1 U589 ( .A1(n642), .A2(n643), .ZN(n644) );
  INV_X1 U590 ( .A(n646), .ZN(n634) );
  XNOR2_X2 U591 ( .A(n619), .B(KEYINPUT0), .ZN(n646) );
  NAND2_X1 U592 ( .A1(n471), .A2(n699), .ZN(n591) );
  XNOR2_X1 U593 ( .A(n714), .B(n367), .ZN(n438) );
  NOR2_X1 U594 ( .A1(n589), .A2(n590), .ZN(n474) );
  XNOR2_X2 U595 ( .A(n439), .B(n564), .ZN(n608) );
  NAND2_X1 U596 ( .A1(n711), .A2(n651), .ZN(n439) );
  XNOR2_X1 U597 ( .A(n549), .B(n548), .ZN(n553) );
  XOR2_X2 U598 ( .A(G122), .B(G104), .Z(n557) );
  NAND2_X1 U599 ( .A1(n633), .A2(n632), .ZN(n445) );
  NAND2_X1 U600 ( .A1(n450), .A2(n760), .ZN(n449) );
  NAND2_X1 U601 ( .A1(n760), .A2(n638), .ZN(n451) );
  AND2_X1 U602 ( .A1(KEYINPUT70), .A2(n458), .ZN(n455) );
  INV_X1 U603 ( .A(KEYINPUT44), .ZN(n458) );
  NAND2_X1 U604 ( .A1(n710), .A2(n469), .ZN(n468) );
  NAND2_X1 U605 ( .A1(n466), .A2(KEYINPUT117), .ZN(n459) );
  NAND2_X1 U606 ( .A1(n354), .A2(n362), .ZN(n465) );
  NAND2_X1 U607 ( .A1(n464), .A2(n460), .ZN(G75) );
  NAND2_X1 U608 ( .A1(n467), .A2(n461), .ZN(n460) );
  XNOR2_X1 U609 ( .A(n647), .B(n473), .ZN(n472) );
  INV_X1 U610 ( .A(KEYINPUT105), .ZN(n473) );
  NAND2_X1 U611 ( .A1(n475), .A2(n761), .ZN(n611) );
  NAND2_X1 U612 ( .A1(n504), .A2(n503), .ZN(n532) );
  AND2_X1 U613 ( .A1(n478), .A2(n437), .ZN(G63) );
  XNOR2_X1 U614 ( .A(n480), .B(n479), .ZN(n478) );
  NAND2_X1 U615 ( .A1(n724), .A2(G478), .ZN(n480) );
  XOR2_X2 U616 ( .A(G116), .B(G107), .Z(n556) );
  XOR2_X1 U617 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n489) );
  OR2_X1 U618 ( .A1(n697), .A2(n649), .ZN(n490) );
  INV_X1 U619 ( .A(KEYINPUT73), .ZN(n630) );
  INV_X1 U620 ( .A(n608), .ZN(n565) );
  INV_X1 U621 ( .A(KEYINPUT2), .ZN(n653) );
  OR2_X1 U622 ( .A1(n653), .A2(n651), .ZN(n491) );
  NAND2_X1 U623 ( .A1(G214), .A2(n563), .ZN(n492) );
  XNOR2_X1 U624 ( .A(KEYINPUT88), .B(n492), .ZN(n698) );
  INV_X1 U625 ( .A(n698), .ZN(n588) );
  XOR2_X1 U626 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n495) );
  NAND2_X1 U627 ( .A1(n651), .A2(G234), .ZN(n493) );
  XNOR2_X1 U628 ( .A(n493), .B(KEYINPUT20), .ZN(n508) );
  NAND2_X1 U629 ( .A1(G221), .A2(n508), .ZN(n494) );
  XNOR2_X1 U630 ( .A(n495), .B(n494), .ZN(n687) );
  XNOR2_X1 U631 ( .A(n496), .B(KEYINPUT14), .ZN(n498) );
  NAND2_X1 U632 ( .A1(n498), .A2(G952), .ZN(n708) );
  NOR2_X1 U633 ( .A1(G953), .A2(n708), .ZN(n616) );
  NAND2_X1 U634 ( .A1(n498), .A2(n497), .ZN(n614) );
  XOR2_X1 U635 ( .A(n614), .B(KEYINPUT103), .Z(n499) );
  NOR2_X1 U636 ( .A1(G900), .A2(n499), .ZN(n500) );
  NOR2_X1 U637 ( .A1(n616), .A2(n500), .ZN(n590) );
  INV_X1 U638 ( .A(KEYINPUT10), .ZN(n501) );
  NAND2_X1 U639 ( .A1(n551), .A2(n501), .ZN(n504) );
  XNOR2_X1 U640 ( .A(G125), .B(G146), .ZN(n502) );
  NAND2_X1 U641 ( .A1(n502), .A2(KEYINPUT10), .ZN(n503) );
  XOR2_X1 U642 ( .A(KEYINPUT90), .B(G128), .Z(n506) );
  XNOR2_X1 U643 ( .A(G119), .B(G110), .ZN(n505) );
  NAND2_X1 U644 ( .A1(n523), .A2(G221), .ZN(n507) );
  NOR2_X1 U645 ( .A1(n727), .A2(G902), .ZN(n512) );
  XOR2_X1 U646 ( .A(KEYINPUT91), .B(KEYINPUT25), .Z(n510) );
  NAND2_X1 U647 ( .A1(G217), .A2(n508), .ZN(n509) );
  XNOR2_X1 U648 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U649 ( .A(KEYINPUT66), .B(G101), .Z(n550) );
  XNOR2_X1 U650 ( .A(G146), .B(n550), .ZN(n513) );
  XNOR2_X1 U651 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U652 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n520) );
  NAND2_X1 U653 ( .A1(n531), .A2(G210), .ZN(n521) );
  XNOR2_X1 U654 ( .A(n571), .B(n522), .ZN(n654) );
  XOR2_X1 U655 ( .A(n556), .B(KEYINPUT9), .Z(n525) );
  NAND2_X1 U656 ( .A1(G217), .A2(n523), .ZN(n524) );
  XNOR2_X1 U657 ( .A(n526), .B(G122), .ZN(n527) );
  XOR2_X1 U658 ( .A(KEYINPUT99), .B(KEYINPUT7), .Z(n528) );
  NOR2_X1 U659 ( .A1(G902), .A2(n725), .ZN(n530) );
  XNOR2_X1 U660 ( .A(KEYINPUT100), .B(G478), .ZN(n529) );
  XOR2_X1 U661 ( .A(n530), .B(n529), .Z(n602) );
  NAND2_X1 U662 ( .A1(G214), .A2(n531), .ZN(n533) );
  XNOR2_X1 U663 ( .A(G113), .B(n557), .ZN(n534) );
  XNOR2_X1 U664 ( .A(n535), .B(n534), .ZN(n543) );
  XNOR2_X1 U665 ( .A(n537), .B(n536), .ZN(n541) );
  XNOR2_X1 U666 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U667 ( .A(n541), .B(n540), .Z(n542) );
  XNOR2_X1 U668 ( .A(n543), .B(n542), .ZN(n722) );
  NOR2_X1 U669 ( .A1(G902), .A2(n722), .ZN(n545) );
  XNOR2_X1 U670 ( .A(KEYINPUT13), .B(G475), .ZN(n544) );
  NAND2_X1 U671 ( .A1(G224), .A2(n750), .ZN(n547) );
  XOR2_X1 U672 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n548) );
  XNOR2_X1 U673 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U674 ( .A(n553), .B(n552), .ZN(n555) );
  XNOR2_X1 U675 ( .A(n555), .B(n554), .ZN(n562) );
  XNOR2_X1 U676 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U677 ( .A(n561), .B(n560), .ZN(n738) );
  XNOR2_X1 U678 ( .A(n562), .B(n738), .ZN(n711) );
  NAND2_X1 U679 ( .A1(n563), .A2(G210), .ZN(n564) );
  NAND2_X1 U680 ( .A1(n606), .A2(n565), .ZN(n566) );
  XNOR2_X1 U681 ( .A(G104), .B(G107), .ZN(n567) );
  NAND2_X1 U682 ( .A1(G227), .A2(n750), .ZN(n569) );
  XNOR2_X1 U683 ( .A(n629), .B(KEYINPUT83), .ZN(n621) );
  NAND2_X1 U684 ( .A1(n574), .A2(n621), .ZN(n676) );
  XNOR2_X1 U685 ( .A(KEYINPUT80), .B(n676), .ZN(n600) );
  INV_X1 U686 ( .A(n602), .ZN(n594) );
  INV_X1 U687 ( .A(n595), .ZN(n601) );
  NOR2_X1 U688 ( .A1(n673), .A2(n592), .ZN(n697) );
  INV_X1 U689 ( .A(KEYINPUT72), .ZN(n575) );
  NOR2_X1 U690 ( .A1(n697), .A2(n575), .ZN(n580) );
  NAND2_X1 U691 ( .A1(n578), .A2(n577), .ZN(n597) );
  NAND2_X1 U692 ( .A1(n580), .A2(n668), .ZN(n581) );
  NAND2_X1 U693 ( .A1(n581), .A2(KEYINPUT47), .ZN(n585) );
  XNOR2_X1 U694 ( .A(KEYINPUT72), .B(n697), .ZN(n582) );
  NOR2_X1 U695 ( .A1(KEYINPUT47), .A2(n582), .ZN(n583) );
  NAND2_X1 U696 ( .A1(n583), .A2(n668), .ZN(n584) );
  NAND2_X1 U697 ( .A1(n585), .A2(n584), .ZN(n599) );
  NAND2_X1 U698 ( .A1(n612), .A2(n592), .ZN(n593) );
  XOR2_X1 U699 ( .A(KEYINPUT41), .B(KEYINPUT108), .Z(n596) );
  NAND2_X1 U700 ( .A1(n699), .A2(n698), .ZN(n696) );
  NAND2_X1 U701 ( .A1(n595), .A2(n594), .ZN(n701) );
  NAND2_X1 U702 ( .A1(n602), .A2(n601), .ZN(n635) );
  OR2_X1 U703 ( .A1(n608), .A2(n635), .ZN(n603) );
  NOR2_X1 U704 ( .A1(n604), .A2(n603), .ZN(n667) );
  XNOR2_X1 U705 ( .A(n667), .B(KEYINPUT78), .ZN(n605) );
  NAND2_X1 U706 ( .A1(n606), .A2(n629), .ZN(n607) );
  XNOR2_X1 U707 ( .A(n607), .B(KEYINPUT43), .ZN(n609) );
  NAND2_X1 U708 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U709 ( .A(KEYINPUT104), .B(n610), .ZN(n761) );
  XNOR2_X1 U710 ( .A(n611), .B(KEYINPUT79), .ZN(n613) );
  NAND2_X1 U711 ( .A1(n612), .A2(n673), .ZN(n679) );
  NAND2_X1 U712 ( .A1(n613), .A2(n679), .ZN(n749) );
  NOR2_X1 U713 ( .A1(G898), .A2(n614), .ZN(n615) );
  NOR2_X1 U714 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U715 ( .A(KEYINPUT76), .B(n640), .ZN(n622) );
  XNOR2_X1 U716 ( .A(n623), .B(KEYINPUT75), .ZN(n624) );
  INV_X1 U717 ( .A(n629), .ZN(n628) );
  XNOR2_X1 U718 ( .A(n642), .B(KEYINPUT101), .ZN(n633) );
  INV_X1 U719 ( .A(n640), .ZN(n632) );
  XNOR2_X2 U720 ( .A(n637), .B(n636), .ZN(n760) );
  NAND2_X1 U721 ( .A1(n641), .A2(n686), .ZN(n657) );
  NAND2_X1 U722 ( .A1(n694), .A2(n646), .ZN(n645) );
  NAND2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U724 ( .A1(n693), .A2(n648), .ZN(n659) );
  NOR2_X1 U725 ( .A1(n674), .A2(n659), .ZN(n649) );
  INV_X1 U726 ( .A(n651), .ZN(n652) );
  NAND2_X1 U727 ( .A1(G472), .A2(n724), .ZN(n655) );
  XOR2_X1 U728 ( .A(G101), .B(KEYINPUT109), .Z(n656) );
  XNOR2_X1 U729 ( .A(n657), .B(n656), .ZN(G3) );
  NAND2_X1 U730 ( .A1(n670), .A2(n659), .ZN(n658) );
  XNOR2_X1 U731 ( .A(n658), .B(G104), .ZN(G6) );
  XNOR2_X1 U732 ( .A(G107), .B(KEYINPUT110), .ZN(n663) );
  XOR2_X1 U733 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n661) );
  NAND2_X1 U734 ( .A1(n659), .A2(n673), .ZN(n660) );
  XNOR2_X1 U735 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U736 ( .A(n663), .B(n662), .ZN(G9) );
  XOR2_X1 U737 ( .A(n356), .B(G110), .Z(G12) );
  XOR2_X1 U738 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n665) );
  NAND2_X1 U739 ( .A1(n668), .A2(n673), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n665), .B(n664), .ZN(n666) );
  XOR2_X1 U741 ( .A(G128), .B(n666), .Z(G30) );
  XOR2_X1 U742 ( .A(G143), .B(n667), .Z(G45) );
  NAND2_X1 U743 ( .A1(n670), .A2(n668), .ZN(n669) );
  XNOR2_X1 U744 ( .A(n669), .B(G146), .ZN(G48) );
  NAND2_X1 U745 ( .A1(n670), .A2(n674), .ZN(n671) );
  XNOR2_X1 U746 ( .A(n671), .B(KEYINPUT112), .ZN(n672) );
  XNOR2_X1 U747 ( .A(G113), .B(n672), .ZN(G15) );
  NAND2_X1 U748 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U749 ( .A(n675), .B(G116), .ZN(G18) );
  XNOR2_X1 U750 ( .A(KEYINPUT113), .B(KEYINPUT37), .ZN(n677) );
  XNOR2_X1 U751 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U752 ( .A(G125), .B(n678), .ZN(G27) );
  XNOR2_X1 U753 ( .A(G134), .B(n679), .ZN(G36) );
  NOR2_X1 U754 ( .A1(n681), .A2(KEYINPUT77), .ZN(n682) );
  NAND2_X1 U755 ( .A1(KEYINPUT2), .A2(n682), .ZN(n683) );
  NAND2_X1 U756 ( .A1(n629), .A2(n684), .ZN(n685) );
  XNOR2_X1 U757 ( .A(KEYINPUT50), .B(n685), .ZN(n691) );
  NOR2_X1 U758 ( .A1(n687), .A2(n686), .ZN(n689) );
  XNOR2_X1 U759 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n688) );
  XNOR2_X1 U760 ( .A(n689), .B(n688), .ZN(n690) );
  NAND2_X1 U761 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n703) );
  NOR2_X1 U763 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U764 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U766 ( .A1(n704), .A2(n680), .ZN(n705) );
  NOR2_X1 U767 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U768 ( .A1(n724), .A2(G210), .ZN(n714) );
  XOR2_X1 U769 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n713) );
  XNOR2_X1 U770 ( .A(n711), .B(KEYINPUT82), .ZN(n712) );
  XOR2_X1 U771 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n717) );
  XNOR2_X1 U772 ( .A(n715), .B(KEYINPUT118), .ZN(n716) );
  XNOR2_X1 U773 ( .A(n717), .B(n716), .ZN(n719) );
  NAND2_X1 U774 ( .A1(n724), .A2(G469), .ZN(n718) );
  XNOR2_X1 U775 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U776 ( .A1(n729), .A2(n720), .ZN(G54) );
  NAND2_X1 U777 ( .A1(n724), .A2(G475), .ZN(n723) );
  XOR2_X1 U778 ( .A(KEYINPUT59), .B(KEYINPUT84), .Z(n721) );
  NAND2_X1 U779 ( .A1(G217), .A2(n724), .ZN(n726) );
  XNOR2_X1 U780 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U781 ( .A1(n729), .A2(n728), .ZN(G66) );
  NAND2_X1 U782 ( .A1(G224), .A2(G953), .ZN(n730) );
  XNOR2_X1 U783 ( .A(n730), .B(KEYINPUT120), .ZN(n731) );
  XNOR2_X1 U784 ( .A(KEYINPUT61), .B(n731), .ZN(n732) );
  NAND2_X1 U785 ( .A1(n732), .A2(G898), .ZN(n733) );
  XNOR2_X1 U786 ( .A(KEYINPUT121), .B(n733), .ZN(n737) );
  NOR2_X1 U787 ( .A1(G953), .A2(n734), .ZN(n735) );
  XNOR2_X1 U788 ( .A(n735), .B(KEYINPUT122), .ZN(n736) );
  NOR2_X1 U789 ( .A1(n737), .A2(n736), .ZN(n744) );
  XNOR2_X1 U790 ( .A(G101), .B(KEYINPUT123), .ZN(n739) );
  XNOR2_X1 U791 ( .A(n739), .B(n738), .ZN(n741) );
  NOR2_X1 U792 ( .A1(G898), .A2(n750), .ZN(n740) );
  NOR2_X1 U793 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U794 ( .A(KEYINPUT124), .B(n742), .Z(n743) );
  XNOR2_X1 U795 ( .A(n744), .B(n743), .ZN(G69) );
  XOR2_X1 U796 ( .A(KEYINPUT125), .B(n745), .Z(n748) );
  XNOR2_X1 U797 ( .A(n746), .B(KEYINPUT89), .ZN(n747) );
  XNOR2_X1 U798 ( .A(n748), .B(n747), .ZN(n752) );
  XNOR2_X1 U799 ( .A(n749), .B(n752), .ZN(n751) );
  NAND2_X1 U800 ( .A1(n751), .A2(n750), .ZN(n756) );
  XNOR2_X1 U801 ( .A(G227), .B(n752), .ZN(n753) );
  NAND2_X1 U802 ( .A1(n753), .A2(G900), .ZN(n754) );
  NAND2_X1 U803 ( .A1(n754), .A2(G953), .ZN(n755) );
  NAND2_X1 U804 ( .A1(n756), .A2(n755), .ZN(G72) );
  XNOR2_X1 U805 ( .A(G137), .B(n757), .ZN(n758) );
  XNOR2_X1 U806 ( .A(n758), .B(KEYINPUT126), .ZN(G39) );
  XOR2_X1 U807 ( .A(n759), .B(G119), .Z(G21) );
  XNOR2_X1 U808 ( .A(n760), .B(G122), .ZN(G24) );
  XNOR2_X1 U809 ( .A(G140), .B(n761), .ZN(G42) );
  XNOR2_X1 U810 ( .A(n762), .B(G131), .ZN(G33) );
endmodule

