//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1284, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1360, new_n1361, new_n1362, new_n1363;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(G355));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n208), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  INV_X1    g0020(.A(new_n201), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G50), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(new_n217), .A2(new_n218), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n224), .B1(new_n217), .B2(new_n218), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  INV_X1    g0026(.A(G68), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  INV_X1    g0028(.A(G87), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n208), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n231));
  INV_X1    g0031(.A(G77), .ZN(new_n232));
  INV_X1    g0032(.A(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G107), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n231), .B1(new_n232), .B2(new_n233), .C1(new_n234), .C2(new_n216), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n212), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT1), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n225), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT67), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G68), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(G58), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT66), .B(G50), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n251), .B(new_n255), .ZN(G351));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(G274), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n262), .B1(new_n264), .B2(new_n240), .ZN(new_n265));
  INV_X1    g0065(.A(G223), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G1698), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT77), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G87), .ZN(new_n273));
  OAI211_X1 g0073(.A(G226), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n267), .B(KEYINPUT77), .C1(new_n269), .C2(new_n268), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n272), .A2(new_n273), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n265), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT78), .ZN(new_n279));
  INV_X1    g0079(.A(G179), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n276), .A2(new_n277), .ZN(new_n282));
  INV_X1    g0082(.A(new_n265), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT78), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n278), .A2(G169), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n281), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT18), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT69), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G58), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n219), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n209), .B2(G20), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n294), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n268), .A2(new_n269), .A3(G20), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT7), .ZN(new_n303));
  OR2_X1    g0103(.A1(KEYINPUT3), .A2(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n210), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT76), .ZN(new_n307));
  AND2_X1   g0107(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n308));
  NOR2_X1   g0108(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n306), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n303), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n307), .B1(new_n306), .B2(new_n310), .ZN(new_n313));
  OAI21_X1  g0113(.A(G68), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(G58), .B(G68), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G20), .A2(G33), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n315), .A2(G20), .B1(G159), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT16), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n227), .B1(new_n306), .B2(KEYINPUT7), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n302), .A2(new_n310), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n317), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT16), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n296), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n301), .B1(new_n318), .B2(new_n324), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n287), .A2(new_n288), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n288), .B1(new_n287), .B2(new_n325), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT79), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n278), .A2(G169), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n279), .B1(new_n278), .B2(new_n280), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n314), .A2(new_n317), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n323), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n295), .A2(new_n219), .ZN(new_n335));
  INV_X1    g0135(.A(new_n317), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n320), .B2(new_n319), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n335), .B1(new_n337), .B2(KEYINPUT16), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n300), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT18), .B1(new_n332), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT79), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n287), .A2(new_n288), .A3(new_n325), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n278), .A2(G200), .ZN(new_n345));
  AOI211_X1 g0145(.A(G190), .B(new_n265), .C1(new_n276), .C2(new_n277), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n344), .B1(new_n325), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g0148(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT76), .B1(new_n302), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(new_n303), .A3(new_n311), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n336), .B1(new_n351), .B2(G68), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n338), .B1(KEYINPUT16), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G190), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n278), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(G200), .B2(new_n278), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n353), .A2(new_n356), .A3(KEYINPUT17), .A4(new_n301), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT80), .B1(new_n348), .B2(new_n357), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n348), .A2(KEYINPUT80), .A3(new_n357), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n328), .B(new_n343), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n361));
  OR2_X1    g0161(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n297), .A2(G50), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(G50), .B2(new_n299), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n316), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n210), .A2(G33), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n294), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n364), .B1(new_n296), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT9), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n277), .A2(new_n261), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT68), .B(G226), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n262), .ZN(new_n373));
  INV_X1    g0173(.A(G1698), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n304), .B2(new_n305), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n268), .A2(new_n269), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n375), .A2(G223), .B1(new_n376), .B2(G77), .ZN(new_n377));
  INV_X1    g0177(.A(G222), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n304), .A2(new_n305), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n374), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n377), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n373), .B1(new_n381), .B2(new_n277), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G190), .ZN(new_n383));
  INV_X1    g0183(.A(G200), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(new_n382), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n361), .B(new_n362), .C1(new_n369), .C2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n385), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT9), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n368), .B(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n387), .A2(new_n389), .A3(KEYINPUT71), .A4(KEYINPUT10), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n382), .ZN(new_n392));
  INV_X1    g0192(.A(G169), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n368), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(G179), .B2(new_n392), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n262), .B1(new_n264), .B2(new_n233), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n375), .A2(G238), .B1(new_n376), .B2(G107), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n240), .B2(new_n380), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n396), .B1(new_n398), .B2(new_n277), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n280), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  XOR2_X1   g0201(.A(KEYINPUT15), .B(G87), .Z(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT70), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT15), .B(G87), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT70), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n403), .A2(new_n210), .A3(G33), .A4(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n289), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(new_n316), .B1(G20), .B2(G77), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n335), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n297), .A2(G77), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(G77), .B2(new_n299), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n399), .A2(G169), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n401), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n410), .A2(new_n412), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(G190), .B2(new_n399), .ZN(new_n417));
  INV_X1    g0217(.A(new_n399), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G200), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n414), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n391), .A2(new_n395), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT13), .ZN(new_n422));
  OAI211_X1 g0222(.A(G232), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT72), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT72), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n379), .A2(new_n425), .A3(G232), .A4(G1698), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G97), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n379), .A2(G226), .A3(new_n374), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n424), .A2(new_n426), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n277), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n262), .B1(new_n264), .B2(new_n228), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n422), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  AOI211_X1 g0233(.A(KEYINPUT13), .B(new_n431), .C1(new_n429), .C2(new_n277), .ZN(new_n434));
  OAI21_X1  g0234(.A(G169), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n430), .A2(new_n432), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT13), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n430), .A2(new_n422), .A3(new_n432), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(G179), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n435), .B2(KEYINPUT14), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT74), .B1(new_n435), .B2(KEYINPUT14), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n437), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n297), .A2(G68), .ZN(new_n445));
  INV_X1    g0245(.A(new_n299), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(KEYINPUT12), .A3(new_n227), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT12), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n299), .B2(G68), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n445), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT73), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n451), .ZN(new_n453));
  INV_X1    g0253(.A(new_n316), .ZN(new_n454));
  OAI22_X1  g0254(.A1(new_n454), .A2(new_n202), .B1(new_n210), .B2(G68), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n366), .A2(new_n232), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n296), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT11), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n457), .A2(new_n458), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n452), .A2(new_n453), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n444), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n439), .A2(G190), .A3(new_n440), .ZN(new_n464));
  OAI21_X1  g0264(.A(G200), .B1(new_n433), .B2(new_n434), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NOR4_X1   g0267(.A1(new_n360), .A2(new_n421), .A3(new_n463), .A4(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n299), .A2(G116), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n209), .A2(G33), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n335), .A2(new_n299), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n469), .B1(new_n471), .B2(G116), .ZN(new_n472));
  INV_X1    g0272(.A(G116), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n295), .A2(new_n219), .B1(G20), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  INV_X1    g0275(.A(G97), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n475), .B(new_n210), .C1(G33), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT20), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n474), .A2(KEYINPUT20), .A3(new_n477), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n472), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n209), .A2(G45), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  XNOR2_X1  g0285(.A(KEYINPUT5), .B(G41), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n277), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n485), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G274), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n277), .A2(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n487), .A2(G270), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(G257), .B(new_n374), .C1(new_n268), .C2(new_n269), .ZN(new_n493));
  INV_X1    g0293(.A(G303), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(new_n379), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT86), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n375), .A2(new_n496), .A3(G264), .ZN(new_n497));
  OAI211_X1 g0297(.A(G264), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT86), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n492), .B1(new_n500), .B2(new_n259), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n483), .B1(new_n501), .B2(G200), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n354), .B2(new_n501), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n393), .B1(new_n472), .B2(new_n482), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n501), .A2(new_n504), .A3(KEYINPUT21), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n497), .A2(new_n499), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n215), .B1(new_n304), .B2(new_n305), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n507), .A2(new_n374), .B1(new_n376), .B2(G303), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n277), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n510), .A2(new_n483), .A3(G179), .A4(new_n492), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n501), .A2(new_n504), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT21), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT87), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT87), .ZN(new_n516));
  AOI211_X1 g0316(.A(new_n516), .B(KEYINPUT21), .C1(new_n501), .C2(new_n504), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n503), .B(new_n512), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n210), .B(G87), .C1(new_n268), .C2(new_n269), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT22), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT22), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n379), .A2(new_n522), .A3(new_n210), .A4(G87), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g0324(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT23), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n210), .B2(G107), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n234), .A2(KEYINPUT23), .A3(G20), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT89), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G116), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(G20), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n210), .A2(KEYINPUT89), .A3(G33), .A4(G116), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n524), .A2(new_n525), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n525), .B1(new_n524), .B2(new_n534), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n296), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT25), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n299), .A2(new_n538), .A3(G107), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n299), .B2(G107), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n471), .A2(G107), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(G257), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n544));
  OAI211_X1 g0344(.A(G250), .B(new_n374), .C1(new_n268), .C2(new_n269), .ZN(new_n545));
  INV_X1    g0345(.A(G294), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n544), .B(new_n545), .C1(new_n257), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n277), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n486), .A2(new_n259), .A3(G274), .A4(new_n485), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n487), .A2(G264), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G169), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n547), .A2(new_n277), .B1(new_n487), .B2(G264), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n553), .A2(G179), .A3(new_n549), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n543), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n551), .A2(G190), .ZN(new_n557));
  AOI21_X1  g0357(.A(G200), .B1(new_n553), .B2(new_n549), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n537), .B(new_n542), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n299), .A2(G97), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n471), .B2(G97), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT6), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n563), .A2(new_n476), .A3(G107), .ZN(new_n564));
  XNOR2_X1  g0364(.A(G97), .B(G107), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n564), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n566), .A2(new_n210), .B1(new_n232), .B2(new_n454), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(G107), .B2(new_n351), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n562), .B1(new_n568), .B2(new_n335), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n488), .A2(G257), .A3(new_n259), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n549), .ZN(new_n571));
  OAI211_X1 g0371(.A(G244), .B(new_n374), .C1(new_n268), .C2(new_n269), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT81), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT4), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n375), .A2(G250), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(new_n574), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n379), .A2(G244), .A3(new_n374), .A4(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n575), .A2(new_n576), .A3(new_n578), .A4(new_n475), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n571), .B1(new_n579), .B2(new_n277), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n280), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n277), .ZN(new_n582));
  INV_X1    g0382(.A(new_n571), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n393), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n569), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n582), .A2(new_n354), .A3(new_n583), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G200), .B2(new_n580), .ZN(new_n588));
  INV_X1    g0388(.A(new_n562), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n351), .A2(G107), .ZN(new_n590));
  INV_X1    g0390(.A(new_n567), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n589), .B1(new_n592), .B2(new_n296), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT82), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n484), .A2(G250), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n277), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n259), .A2(KEYINPUT82), .A3(G250), .A4(new_n484), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n259), .A2(G274), .A3(new_n485), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n379), .A2(G238), .A3(new_n374), .ZN(new_n602));
  OAI211_X1 g0402(.A(G244), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n603), .A3(new_n531), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n277), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n393), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n600), .B1(new_n277), .B2(new_n604), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n280), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n403), .A2(new_n406), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n446), .ZN(new_n611));
  XNOR2_X1  g0411(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n427), .A2(new_n210), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n229), .A2(new_n476), .A3(new_n234), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT19), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n616), .A2(KEYINPUT83), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(KEYINPUT83), .ZN(new_n618));
  OAI22_X1  g0418(.A1(new_n617), .A2(new_n618), .B1(new_n366), .B2(new_n476), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n210), .B(G68), .C1(new_n268), .C2(new_n269), .ZN(new_n621));
  OR2_X1    g0421(.A1(new_n621), .A2(KEYINPUT84), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(KEYINPUT84), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n611), .B1(new_n624), .B2(new_n335), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n403), .A2(new_n406), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(KEYINPUT85), .A3(new_n471), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT85), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n335), .A2(new_n299), .A3(new_n470), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n628), .B1(new_n610), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n607), .B(new_n609), .C1(new_n625), .C2(new_n631), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n621), .B(KEYINPUT84), .ZN(new_n633));
  INV_X1    g0433(.A(new_n620), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n335), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n611), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n606), .A2(G200), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n608), .A2(G190), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n629), .A2(new_n229), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n637), .A2(new_n638), .A3(new_n639), .A4(new_n641), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n586), .A2(new_n594), .A3(new_n632), .A4(new_n642), .ZN(new_n643));
  AND4_X1   g0443(.A1(new_n468), .A2(new_n519), .A3(new_n560), .A4(new_n643), .ZN(G372));
  INV_X1    g0444(.A(new_n395), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n326), .A2(new_n327), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n463), .B1(new_n466), .B2(new_n414), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n359), .A2(new_n358), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n645), .B1(new_n649), .B2(new_n391), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n642), .A2(new_n632), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT26), .B1(new_n651), .B2(new_n586), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n569), .A2(new_n581), .A3(new_n585), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n600), .A2(KEYINPUT90), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT90), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n597), .A2(new_n598), .A3(new_n655), .A4(new_n599), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n605), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n393), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n633), .A2(new_n634), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n296), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n661), .A2(new_n611), .A3(new_n630), .A4(new_n627), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n659), .A2(new_n662), .A3(new_n609), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n635), .A2(new_n636), .A3(new_n640), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n654), .A2(new_n656), .B1(new_n277), .B2(new_n604), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n665), .B(new_n639), .C1(new_n384), .C2(new_n666), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n653), .A2(new_n663), .A3(new_n664), .A4(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n652), .A2(new_n668), .A3(new_n663), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n488), .A2(new_n259), .ZN(new_n671));
  INV_X1    g0471(.A(G270), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n549), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n509), .B2(new_n277), .ZN(new_n674));
  INV_X1    g0474(.A(new_n481), .ZN(new_n675));
  AOI21_X1  g0475(.A(KEYINPUT20), .B1(new_n474), .B2(new_n477), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n469), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n629), .B2(new_n473), .ZN(new_n679));
  OAI21_X1  g0479(.A(G169), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n514), .B1(new_n674), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n516), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n513), .A2(KEYINPUT87), .A3(new_n514), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n543), .A2(KEYINPUT91), .A3(new_n555), .ZN(new_n685));
  AOI21_X1  g0485(.A(KEYINPUT91), .B1(new_n543), .B2(new_n555), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n684), .B(new_n512), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n594), .A2(new_n586), .A3(new_n559), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n665), .A2(new_n639), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n666), .A2(new_n384), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n609), .B1(new_n625), .B2(new_n631), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n666), .A2(G169), .ZN(new_n692));
  OAI22_X1  g0492(.A1(new_n689), .A2(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n670), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n468), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n650), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT92), .ZN(G369));
  NAND3_X1  g0499(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G213), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G343), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n483), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n518), .B2(KEYINPUT93), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(KEYINPUT93), .B2(new_n518), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n684), .A2(new_n512), .A3(new_n707), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n543), .A2(new_n705), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n560), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n543), .A2(new_n555), .A3(new_n705), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(KEYINPUT94), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n714), .A2(KEYINPUT94), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n713), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n711), .A2(G330), .A3(new_n717), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n685), .A2(new_n686), .A3(new_n705), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n705), .B1(new_n684), .B2(new_n512), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n719), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n718), .A2(new_n721), .ZN(G399));
  NOR2_X1   g0522(.A1(new_n214), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n614), .A2(G116), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n222), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT95), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  INV_X1    g0529(.A(new_n705), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n696), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n594), .A2(new_n586), .A3(new_n559), .ZN(new_n734));
  INV_X1    g0534(.A(new_n693), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n512), .B(new_n556), .C1(new_n515), .C2(new_n517), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n664), .B1(new_n651), .B2(new_n586), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n653), .A2(new_n663), .A3(KEYINPUT26), .A4(new_n667), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(new_n740), .A3(new_n663), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n733), .B1(new_n741), .B2(new_n730), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n732), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G330), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n580), .A2(new_n553), .A3(new_n608), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n510), .A2(G179), .A3(new_n492), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n259), .B1(new_n506), .B2(new_n508), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n749), .A2(new_n280), .A3(new_n673), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n553), .A2(new_n601), .A3(new_n605), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT30), .A4(new_n580), .ZN(new_n752));
  AOI21_X1  g0552(.A(G179), .B1(new_n582), .B2(new_n583), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n658), .A2(new_n753), .A3(new_n501), .A4(new_n551), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n748), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  AND3_X1   g0555(.A1(new_n755), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n756));
  AOI21_X1  g0556(.A(KEYINPUT31), .B1(new_n755), .B2(new_n705), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n519), .A2(new_n643), .A3(new_n560), .A4(new_n730), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n744), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n743), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n729), .B1(new_n763), .B2(G1), .ZN(G364));
  NAND2_X1  g0564(.A1(new_n711), .A2(G330), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G13), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n209), .B1(new_n768), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n723), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n711), .A2(G330), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n711), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n771), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n213), .A2(new_n379), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n781), .A2(new_n206), .B1(G116), .B2(new_n213), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n255), .A2(G45), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT96), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n214), .A2(new_n379), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(new_n260), .B2(new_n223), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n782), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n219), .B1(G20), .B2(new_n393), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n777), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n210), .A2(G179), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G190), .A2(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G159), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT32), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n210), .A2(new_n280), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n794), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n376), .B(new_n799), .C1(G77), .C2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n800), .A2(G190), .A3(new_n384), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT97), .Z(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G58), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n800), .A2(G200), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G190), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n793), .A2(G190), .A3(G200), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n810), .A2(new_n227), .B1(new_n229), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n808), .A2(new_n354), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n793), .A2(new_n354), .A3(G200), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n814), .A2(new_n202), .B1(new_n815), .B2(new_n234), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n280), .A2(new_n384), .A3(G190), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(G20), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n797), .A2(new_n798), .B1(G97), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n803), .A2(new_n807), .A3(new_n817), .A4(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n802), .A2(G311), .B1(G294), .B2(new_n819), .ZN(new_n822));
  INV_X1    g0622(.A(G326), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n823), .B2(new_n814), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT98), .Z(new_n825));
  INV_X1    g0625(.A(G317), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(KEYINPUT33), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n826), .A2(KEYINPUT33), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n809), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G283), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n830), .B2(new_n815), .C1(new_n494), .C2(new_n811), .ZN(new_n831));
  INV_X1    g0631(.A(G329), .ZN(new_n832));
  INV_X1    g0632(.A(G322), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n376), .B1(new_n795), .B2(new_n832), .C1(new_n804), .C2(new_n833), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n821), .B1(new_n825), .B2(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n780), .B(new_n792), .C1(new_n789), .C2(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n772), .A2(new_n774), .B1(new_n779), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G396));
  INV_X1    g0639(.A(new_n413), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n840), .A2(KEYINPUT99), .A3(new_n400), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT99), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n401), .B2(new_n413), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n419), .B2(new_n417), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n687), .A2(new_n694), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n730), .B(new_n845), .C1(new_n846), .C2(new_n669), .ZN(new_n847));
  INV_X1    g0647(.A(new_n731), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n419), .B(new_n415), .C1(new_n354), .C2(new_n418), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n416), .A2(new_n705), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n841), .A2(new_n849), .A3(new_n843), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n414), .A2(new_n705), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n847), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n771), .B1(new_n854), .B2(new_n761), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n761), .B2(new_n854), .ZN(new_n856));
  INV_X1    g0656(.A(new_n789), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n813), .A2(G137), .B1(new_n802), .B2(G159), .ZN(new_n858));
  INV_X1    g0658(.A(G150), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n858), .B1(new_n859), .B2(new_n810), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G143), .B2(new_n806), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT34), .ZN(new_n862));
  INV_X1    g0662(.A(G132), .ZN(new_n863));
  INV_X1    g0663(.A(new_n819), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n379), .B1(new_n863), .B2(new_n795), .C1(new_n864), .C2(new_n292), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n202), .A2(new_n811), .B1(new_n815), .B2(new_n227), .ZN(new_n866));
  OR3_X1    g0666(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n811), .A2(new_n234), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n815), .A2(new_n229), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n868), .B(new_n869), .C1(G283), .C2(new_n809), .ZN(new_n870));
  INV_X1    g0670(.A(new_n795), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n379), .B1(new_n871), .B2(G311), .ZN(new_n872));
  INV_X1    g0672(.A(new_n804), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n873), .A2(G294), .B1(new_n802), .B2(G116), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n813), .A2(G303), .B1(G97), .B2(new_n819), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n870), .A2(new_n872), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n857), .B1(new_n867), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n789), .A2(new_n775), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n780), .B(new_n877), .C1(new_n232), .C2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n776), .B2(new_n853), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n856), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(G384));
  NOR2_X1   g0682(.A1(new_n768), .A2(new_n209), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n844), .A2(new_n730), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT100), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n461), .A2(new_n705), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n466), .B(new_n886), .C1(new_n444), .C2(new_n462), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n435), .A2(KEYINPUT14), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT74), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n435), .A2(KEYINPUT14), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n890), .A2(new_n891), .A3(new_n436), .A4(new_n441), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n461), .B(new_n705), .C1(new_n892), .C2(new_n467), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n847), .A2(new_n885), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n322), .A2(new_n323), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n300), .B1(new_n338), .B2(new_n896), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n325), .A2(new_n347), .B1(new_n897), .B2(new_n703), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n330), .A2(new_n331), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n897), .B1(new_n899), .B2(new_n281), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT37), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n287), .A2(new_n325), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n339), .A2(new_n356), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT37), .ZN(new_n904));
  INV_X1    g0704(.A(new_n703), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n325), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n902), .A2(new_n903), .A3(new_n904), .A4(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n897), .A2(new_n703), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n895), .B(new_n908), .C1(new_n360), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n328), .A2(new_n343), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n910), .B1(new_n912), .B2(new_n648), .ZN(new_n913));
  INV_X1    g0713(.A(new_n908), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n894), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n703), .B1(new_n326), .B2(new_n327), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n913), .A2(KEYINPUT38), .A3(new_n914), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n340), .A2(new_n348), .A3(new_n357), .A4(new_n342), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n325), .A3(new_n905), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n902), .A2(new_n903), .A3(new_n906), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT37), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n907), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT39), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n913), .A2(new_n914), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n895), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(KEYINPUT39), .A3(new_n918), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n444), .A2(new_n462), .A3(new_n705), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n916), .B(new_n917), .C1(new_n931), .C2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n468), .B1(new_n732), .B2(new_n742), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n650), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n934), .B(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n908), .B1(new_n360), .B2(new_n910), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n924), .B1(new_n938), .B2(KEYINPUT38), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n887), .A2(new_n893), .ZN(new_n940));
  INV_X1    g0740(.A(new_n853), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n758), .B2(new_n759), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT40), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n758), .A2(new_n759), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n468), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT40), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n940), .A2(new_n942), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n911), .B2(new_n915), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n944), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n944), .A2(new_n949), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(new_n468), .A3(new_n945), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n950), .A2(G330), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n883), .B1(new_n937), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n937), .B2(new_n953), .ZN(new_n955));
  INV_X1    g0755(.A(new_n566), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT35), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(KEYINPUT35), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n957), .A2(G116), .A3(new_n220), .A4(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT36), .ZN(new_n960));
  OAI21_X1  g0760(.A(G77), .B1(new_n292), .B2(new_n227), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n222), .A2(new_n961), .B1(G50), .B2(new_n227), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(G1), .A3(new_n767), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n955), .A2(new_n960), .A3(new_n963), .ZN(G367));
  OAI221_X1 g0764(.A(new_n790), .B1(new_n213), .B2(new_n610), .C1(new_n786), .C2(new_n246), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n965), .A2(new_n771), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n815), .A2(new_n232), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n811), .A2(new_n292), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(G68), .C2(new_n819), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n376), .B1(new_n873), .B2(G150), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G50), .A2(new_n802), .B1(new_n871), .B2(G137), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G143), .A2(new_n813), .B1(new_n809), .B2(G159), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n815), .A2(new_n476), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n379), .B(new_n974), .C1(G317), .C2(new_n871), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT105), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(KEYINPUT105), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n809), .A2(G294), .B1(new_n802), .B2(G283), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n813), .A2(G311), .B1(G107), .B2(new_n819), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n976), .A2(new_n977), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n811), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(KEYINPUT46), .A3(G116), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT46), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n811), .B2(new_n473), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n982), .B(new_n984), .C1(new_n805), .C2(new_n494), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n973), .B1(new_n980), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT47), .Z(new_n987));
  NOR2_X1   g0787(.A1(new_n665), .A2(new_n730), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n735), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n663), .B2(new_n988), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT101), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n966), .B1(new_n857), .B2(new_n987), .C1(new_n991), .C2(new_n778), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n594), .B(new_n586), .C1(new_n593), .C2(new_n730), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n653), .A2(new_n705), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n721), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT45), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n995), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n717), .A2(new_n720), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI211_X1 g0801(.A(KEYINPUT44), .B(new_n999), .C1(new_n1001), .C2(new_n719), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT44), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n721), .B2(new_n995), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1004), .A3(KEYINPUT103), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(KEYINPUT103), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n998), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT104), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n718), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n717), .A2(new_n720), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n1000), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n765), .A2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n711), .A2(G330), .A3(new_n1000), .A4(new_n1012), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n762), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n998), .A2(new_n1005), .A3(new_n1006), .A4(new_n718), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n718), .A2(KEYINPUT104), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n763), .B1(new_n1011), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n723), .B(KEYINPUT41), .Z(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n770), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  OR3_X1    g0826(.A1(new_n718), .A2(KEYINPUT102), .A3(new_n999), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT102), .B1(new_n718), .B2(new_n999), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n993), .A2(new_n556), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n705), .B1(new_n1032), .B2(new_n586), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1001), .A2(new_n995), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1033), .B1(new_n1034), .B2(KEYINPUT42), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(KEYINPUT42), .B2(new_n1034), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1027), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1030), .A2(new_n1031), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1031), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1037), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1039), .B1(new_n1040), .B2(new_n1029), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n992), .B1(new_n1024), .B2(new_n1042), .ZN(G387));
  AND2_X1   g0843(.A1(new_n762), .A2(new_n1016), .ZN(new_n1044));
  OR3_X1    g0844(.A1(new_n1044), .A2(new_n1017), .A3(new_n724), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1014), .A2(new_n770), .A3(new_n1015), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT106), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n781), .A2(new_n725), .B1(G107), .B2(new_n213), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT107), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n243), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n408), .A2(new_n202), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT50), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n725), .B(new_n260), .C1(new_n227), .C2(new_n232), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n785), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1050), .A2(G45), .B1(KEYINPUT108), .B2(new_n1054), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(KEYINPUT108), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1049), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n771), .B1(new_n1057), .B2(new_n791), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n809), .A2(G311), .B1(new_n802), .B2(G303), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n833), .B2(new_n814), .C1(new_n805), .C2(new_n826), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n981), .A2(G294), .B1(new_n819), .B2(G283), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n376), .B1(new_n795), .B2(new_n823), .C1(new_n473), .C2(new_n815), .ZN(new_n1069));
  OR3_X1    g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n379), .B1(new_n801), .B2(new_n227), .C1(new_n202), .C2(new_n804), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n974), .B(new_n1071), .C1(G159), .C2(new_n813), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n981), .A2(G77), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n859), .B2(new_n795), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT109), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n294), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n626), .A2(new_n819), .B1(new_n1076), .B2(new_n809), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1072), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1070), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1058), .B1(new_n1079), .B2(new_n789), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n717), .B2(new_n778), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1045), .A2(new_n1047), .A3(new_n1081), .ZN(G393));
  NAND2_X1  g0882(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT110), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n1084), .A3(new_n1018), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1007), .A2(KEYINPUT110), .A3(new_n1009), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(new_n762), .C2(new_n1016), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n724), .B1(new_n1088), .B2(new_n1010), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT113), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n769), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n999), .A2(new_n777), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n251), .A2(new_n785), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n790), .B1(new_n476), .B2(new_n213), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n771), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n809), .A2(G50), .B1(new_n802), .B2(new_n408), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1098), .A2(KEYINPUT111), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(KEYINPUT111), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n376), .B(new_n869), .C1(G143), .C2(new_n871), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n981), .A2(G68), .B1(new_n819), .B2(G77), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G150), .A2(new_n813), .B1(new_n873), .B2(G159), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT51), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n810), .A2(new_n494), .B1(new_n815), .B2(new_n234), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n376), .B1(new_n795), .B2(new_n833), .C1(new_n801), .C2(new_n546), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n864), .A2(new_n473), .B1(new_n811), .B2(new_n830), .ZN(new_n1108));
  OR3_X1    g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G317), .A2(new_n813), .B1(new_n873), .B2(G311), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1110), .B(new_n1111), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1103), .A2(new_n1105), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1096), .B1(new_n1113), .B2(new_n789), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1092), .B1(new_n1093), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT113), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1087), .A2(new_n1089), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1091), .A2(new_n1115), .A3(new_n1117), .ZN(G390));
  INV_X1    g0918(.A(new_n878), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n813), .A2(G283), .B1(new_n802), .B2(G97), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n234), .B2(new_n810), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT117), .Z(new_n1122));
  OAI22_X1  g0922(.A1(new_n227), .A2(new_n815), .B1(new_n811), .B2(new_n229), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n376), .B1(new_n795), .B2(new_n546), .C1(new_n804), .C2(new_n473), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(G77), .C2(new_n819), .ZN(new_n1125));
  INV_X1    g0925(.A(G137), .ZN(new_n1126));
  INV_X1    g0926(.A(G128), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n810), .A2(new_n1126), .B1(new_n814), .B2(new_n1127), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n864), .A2(new_n796), .B1(new_n815), .B2(new_n202), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT53), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n981), .B2(G150), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT54), .B(G143), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n804), .A2(new_n863), .B1(new_n801), .B2(new_n1133), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n811), .A2(KEYINPUT53), .A3(new_n859), .ZN(new_n1135));
  INV_X1    g0935(.A(G125), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n379), .B1(new_n795), .B2(new_n1136), .ZN(new_n1137));
  NOR4_X1   g0937(.A1(new_n1132), .A2(new_n1134), .A3(new_n1135), .A4(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1122), .A2(new_n1125), .B1(new_n1130), .B2(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n771), .B1(new_n1076), .B2(new_n1119), .C1(new_n1139), .C2(new_n857), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n931), .B2(new_n775), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n940), .A2(new_n760), .A3(new_n853), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT116), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n894), .A2(new_n932), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n927), .B2(new_n930), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n932), .A2(KEYINPUT114), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n932), .A2(KEYINPUT114), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(new_n911), .C2(new_n924), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT115), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n940), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n741), .A2(new_n730), .A3(new_n845), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n885), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n887), .A2(new_n893), .A3(KEYINPUT115), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1153), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1148), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1145), .B1(new_n1147), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT39), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n911), .A2(new_n915), .A3(new_n1160), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n1161), .A2(new_n926), .B1(new_n932), .B2(new_n894), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n939), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1153), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1164), .A2(new_n1165), .B1(new_n1144), .B2(new_n1143), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1145), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1162), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1159), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1141), .B1(new_n1169), .B2(new_n770), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1143), .A2(new_n1155), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n760), .A2(new_n853), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1153), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1156), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1172), .A2(new_n887), .A3(new_n893), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n1142), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n847), .A2(new_n885), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1171), .A2(new_n1175), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n468), .A2(new_n760), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n650), .A2(new_n935), .A3(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n723), .B1(new_n1169), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1181), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n1159), .B2(new_n1168), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1170), .B1(new_n1183), .B2(new_n1189), .ZN(G378));
  NAND3_X1  g0990(.A1(new_n386), .A2(new_n390), .A3(new_n395), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n368), .A2(new_n703), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1193), .B(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n951), .B2(G330), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n744), .B(new_n1195), .C1(new_n944), .C2(new_n949), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n934), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n918), .A2(new_n925), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n943), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n947), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n940), .A2(new_n942), .A3(new_n947), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n929), .B2(new_n918), .ZN(new_n1204));
  OAI21_X1  g1004(.A(G330), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1195), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n916), .A2(new_n917), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n911), .A2(new_n915), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n926), .B1(new_n1208), .B2(KEYINPUT39), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1207), .B1(new_n1209), .B2(new_n932), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n951), .A2(G330), .A3(new_n1196), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1206), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1199), .A2(KEYINPUT119), .A3(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT119), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1206), .A2(new_n1210), .A3(new_n1211), .A4(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n770), .A3(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n771), .B1(new_n1119), .B2(G50), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n379), .A2(G41), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G50), .B(new_n1218), .C1(new_n257), .C2(new_n258), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n815), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(G58), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n871), .A2(G283), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1073), .A2(new_n1221), .A3(new_n1218), .A4(new_n1222), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT118), .Z(new_n1224));
  AOI22_X1  g1024(.A1(G97), .A2(new_n809), .B1(new_n813), .B2(G116), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n873), .A2(G107), .B1(G68), .B2(new_n819), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(new_n610), .C2(new_n801), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1224), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1219), .B1(new_n1228), .B2(KEYINPUT58), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n804), .A2(new_n1127), .B1(new_n801), .B2(new_n1126), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n813), .A2(G125), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n811), .B2(new_n1133), .C1(new_n810), .C2(new_n863), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1230), .B(new_n1232), .C1(G150), .C2(new_n819), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1220), .A2(G159), .ZN(new_n1236));
  AOI211_X1 g1036(.A(G33), .B(G41), .C1(new_n871), .C2(G124), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1229), .B1(KEYINPUT58), .B2(new_n1228), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1217), .B1(new_n1240), .B2(new_n789), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1196), .B2(new_n776), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1216), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT57), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1189), .A2(new_n1181), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1245), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1199), .A2(KEYINPUT120), .A3(new_n1212), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT120), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1251), .B(new_n934), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT57), .B1(new_n1189), .B2(new_n1181), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n723), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1244), .B1(new_n1249), .B2(new_n1255), .ZN(G375));
  NAND2_X1  g1056(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1188), .A2(new_n1257), .A3(new_n1023), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n775), .B1(new_n1174), .B2(new_n1173), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n780), .B1(new_n227), .B2(new_n878), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n379), .B1(new_n795), .B2(new_n1127), .C1(new_n801), .C2(new_n859), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n813), .A2(G132), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT121), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1261), .B(new_n1263), .C1(G137), .C2(new_n806), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n810), .A2(new_n1133), .B1(new_n202), .B2(new_n864), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1221), .B1(new_n796), .B2(new_n811), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n810), .A2(new_n473), .B1(new_n476), .B2(new_n811), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n967), .B(new_n1268), .C1(G294), .C2(new_n813), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n376), .B1(new_n795), .B2(new_n494), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n804), .A2(new_n830), .B1(new_n801), .B2(new_n234), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1270), .B(new_n1271), .C1(new_n626), .C2(new_n819), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1264), .A2(new_n1267), .B1(new_n1269), .B2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1259), .B(new_n1260), .C1(new_n857), .C2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1179), .B2(new_n769), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1258), .A2(new_n1276), .ZN(G381));
  NAND4_X1  g1077(.A1(new_n1045), .A2(new_n838), .A3(new_n1047), .A4(new_n1081), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1278), .A2(G384), .ZN(new_n1279));
  XOR2_X1   g1079(.A(new_n1279), .B(KEYINPUT122), .Z(new_n1280));
  OR3_X1    g1080(.A1(new_n1280), .A2(G387), .A3(G381), .ZN(new_n1281));
  OR4_X1    g1081(.A1(G390), .A2(new_n1281), .A3(G378), .A4(G375), .ZN(G407));
  NAND2_X1  g1082(.A1(new_n704), .A2(G213), .ZN(new_n1283));
  OR2_X1    g1083(.A1(G378), .A2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G407), .B(G213), .C1(G375), .C2(new_n1284), .ZN(G409));
  OAI21_X1  g1085(.A(KEYINPUT60), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n724), .B1(new_n1286), .B2(new_n1257), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1179), .A2(KEYINPUT60), .A3(new_n1181), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT124), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT124), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1287), .A2(new_n1291), .A3(new_n1288), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(G384), .B1(new_n1293), .B2(new_n1276), .ZN(new_n1294));
  AOI211_X1 g1094(.A(new_n881), .B(new_n1275), .C1(new_n1290), .C2(new_n1292), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(G378), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1169), .A2(new_n1182), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1245), .B1(new_n1299), .B2(new_n1187), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n724), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n1297), .B(new_n1243), .C1(new_n1301), .C2(new_n1248), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(new_n1187), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1303), .A2(new_n1023), .A3(new_n1215), .A4(new_n1213), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1304), .A2(new_n1242), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1253), .A2(KEYINPUT123), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT123), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1250), .A2(new_n1307), .A3(new_n1252), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1306), .A2(new_n770), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(G378), .B1(new_n1305), .B2(new_n1309), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1283), .B(new_n1296), .C1(new_n1302), .C2(new_n1310), .ZN(new_n1311));
  XOR2_X1   g1111(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1283), .B1(new_n1302), .B2(new_n1310), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n704), .A2(G213), .A3(G2897), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1292), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1291), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1276), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n881), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1293), .A2(G384), .A3(new_n1276), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1315), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1316), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1314), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT61), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1306), .A2(new_n770), .A3(new_n1308), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1304), .A2(new_n1242), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1297), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  OAI211_X1 g1129(.A(G378), .B(new_n1244), .C1(new_n1249), .C2(new_n1255), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT62), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1331), .A2(new_n1332), .A3(new_n1283), .A4(new_n1296), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1313), .A2(new_n1325), .A3(new_n1326), .A4(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(G393), .A2(G396), .ZN(new_n1335));
  AOI21_X1  g1135(.A(G387), .B1(new_n1278), .B2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1278), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1042), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1088), .A2(new_n1010), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1022), .B1(new_n1339), .B2(new_n763), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1338), .B1(new_n1340), .B2(new_n770), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1337), .B1(new_n1341), .B2(new_n992), .ZN(new_n1342));
  OAI21_X1  g1142(.A(G390), .B1(new_n1336), .B2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(G390), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(G387), .A2(new_n1278), .A3(new_n1335), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1341), .A2(new_n1337), .A3(new_n992), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1344), .A2(new_n1345), .A3(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1343), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1334), .A2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT125), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1324), .A2(new_n1350), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1316), .A2(new_n1323), .A3(KEYINPUT125), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1351), .A2(new_n1314), .A3(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT63), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1311), .A2(new_n1354), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1331), .A2(KEYINPUT63), .A3(new_n1283), .A4(new_n1296), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1348), .A2(KEYINPUT61), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1353), .A2(new_n1355), .A3(new_n1356), .A4(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1349), .A2(new_n1358), .ZN(G405));
  NAND2_X1  g1159(.A1(new_n1296), .A2(KEYINPUT127), .ZN(new_n1360));
  XNOR2_X1  g1160(.A(new_n1348), .B(new_n1360), .ZN(new_n1361));
  AND2_X1   g1161(.A1(G375), .A2(new_n1297), .ZN(new_n1362));
  OAI22_X1  g1162(.A1(new_n1362), .A2(new_n1302), .B1(KEYINPUT127), .B2(new_n1296), .ZN(new_n1363));
  XNOR2_X1  g1163(.A(new_n1361), .B(new_n1363), .ZN(G402));
endmodule


