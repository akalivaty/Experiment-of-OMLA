//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT65), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G50), .A2(G226), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n202), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n208), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n206), .A2(KEYINPUT64), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT64), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n208), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  NOR3_X1   g0028(.A1(new_n218), .A2(new_n225), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G58), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G116), .ZN(new_n242));
  INV_X1    g0042(.A(G107), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G97), .ZN(new_n244));
  INV_X1    g0044(.A(G97), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G107), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n242), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  AND2_X1   g0047(.A1(G97), .A2(G107), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G97), .A2(G107), .ZN(new_n249));
  OR2_X1    g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n247), .B1(new_n242), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n241), .B(new_n251), .ZN(G351));
  XNOR2_X1  g0052(.A(KEYINPUT64), .B(G20), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  OAI21_X1  g0054(.A(KEYINPUT67), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT67), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n220), .A2(G20), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n206), .A2(KEYINPUT64), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n256), .B(G33), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  XOR2_X1   g0059(.A(KEYINPUT8), .B(G58), .Z(new_n260));
  NAND3_X1  g0060(.A1(new_n255), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G150), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n261), .B1(new_n206), .B2(new_n201), .C1(new_n262), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n223), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n266), .B1(new_n207), .B2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G50), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n267), .B1(G1), .B2(new_n206), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G50), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n269), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT9), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n265), .A2(new_n268), .B1(new_n272), .B2(new_n271), .ZN(new_n280));
  AOI21_X1  g0080(.A(KEYINPUT9), .B1(new_n280), .B2(new_n276), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT69), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(KEYINPUT10), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n205), .B(G274), .C1(G41), .C2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  OAI211_X1 g0087(.A(G1), .B(G13), .C1(new_n254), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G226), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n286), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n292), .A2(KEYINPUT66), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT3), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n254), .ZN(new_n295));
  NAND2_X1  g0095(.A1(KEYINPUT3), .A2(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G1698), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G222), .ZN(new_n299));
  INV_X1    g0099(.A(G223), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n297), .B(new_n299), .C1(new_n300), .C2(new_n298), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n301), .B(new_n302), .C1(G77), .C2(new_n297), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n292), .A2(KEYINPUT66), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n293), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n305), .A2(G200), .B1(new_n283), .B2(KEYINPUT10), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n282), .A2(new_n285), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n277), .A2(new_n278), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n280), .A2(KEYINPUT9), .A3(new_n276), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n310), .A2(new_n307), .A3(new_n311), .A4(new_n308), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n284), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n305), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n277), .B(new_n315), .C1(G179), .C2(new_n305), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n309), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  XOR2_X1   g0117(.A(KEYINPUT15), .B(G87), .Z(new_n318));
  NAND3_X1  g0118(.A1(new_n255), .A2(new_n259), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT68), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n319), .A2(new_n320), .B1(new_n260), .B2(new_n263), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n321), .B1(new_n320), .B2(new_n319), .C1(new_n202), .C2(new_n222), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n268), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n270), .A2(G77), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n275), .A2(G77), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G238), .A2(G1698), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n297), .B(new_n328), .C1(new_n231), .C2(G1698), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n329), .B(new_n302), .C1(G107), .C2(new_n297), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n330), .B(new_n286), .C1(new_n215), .C2(new_n290), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n314), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n331), .A2(G179), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n327), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n324), .B1(new_n322), .B2(new_n268), .ZN(new_n336));
  OR2_X1    g0136(.A1(new_n331), .A2(new_n306), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n331), .A2(G200), .ZN(new_n338));
  AND4_X1   g0138(.A1(new_n336), .A2(new_n326), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  OR4_X1    g0139(.A1(KEYINPUT70), .A2(new_n317), .A3(new_n335), .A4(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n255), .A2(G77), .A3(new_n259), .ZN(new_n341));
  INV_X1    g0141(.A(G68), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G20), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n263), .A2(G50), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n268), .ZN(new_n346));
  XOR2_X1   g0146(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G13), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n343), .A2(G1), .A3(new_n350), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n351), .A2(KEYINPUT12), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n345), .A2(new_n268), .A3(new_n347), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n275), .A2(G68), .B1(KEYINPUT12), .B2(new_n351), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n349), .A2(new_n352), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n291), .A2(new_n298), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n231), .A2(G1698), .ZN(new_n358));
  AND2_X1   g0158(.A1(KEYINPUT3), .A2(G33), .ZN(new_n359));
  NOR2_X1   g0159(.A1(KEYINPUT3), .A2(G33), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n357), .B(new_n358), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G97), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT71), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT71), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(G33), .A3(G97), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n302), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n288), .A2(new_n289), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G238), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n286), .B(KEYINPUT72), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT13), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT13), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n368), .A2(new_n370), .A3(new_n374), .A4(new_n371), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G200), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT74), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT73), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n373), .A2(new_n379), .A3(new_n375), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n372), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n378), .B1(new_n382), .B2(G190), .ZN(new_n383));
  AOI211_X1 g0183(.A(KEYINPUT74), .B(new_n306), .C1(new_n380), .C2(new_n381), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n356), .B(new_n377), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n355), .A2(KEYINPUT76), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n353), .A2(new_n354), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT76), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n387), .A2(new_n388), .A3(new_n352), .A4(new_n349), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n376), .A2(G169), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT14), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n375), .A2(new_n379), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n302), .A2(new_n367), .B1(new_n369), .B2(G238), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n374), .B1(new_n394), .B2(new_n371), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n381), .ZN(new_n397));
  OAI21_X1  g0197(.A(G179), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT14), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n376), .A2(new_n399), .A3(G169), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n392), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n390), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n385), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n312), .B(new_n285), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n336), .A2(new_n326), .A3(new_n337), .A4(new_n338), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n316), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT70), .B1(new_n407), .B2(new_n335), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n274), .A2(new_n260), .ZN(new_n409));
  INV_X1    g0209(.A(new_n260), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n270), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n359), .A2(new_n360), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT7), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n222), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n295), .A2(new_n206), .A3(new_n296), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT7), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n418), .A3(G68), .ZN(new_n419));
  XNOR2_X1  g0219(.A(G58), .B(G68), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(G20), .B1(G159), .B2(new_n263), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(KEYINPUT16), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n422), .A2(new_n268), .ZN(new_n423));
  XOR2_X1   g0223(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n222), .A2(new_n414), .A3(KEYINPUT7), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n417), .A2(new_n415), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n342), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n421), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n413), .B1(new_n423), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n288), .A2(G232), .A3(new_n289), .ZN(new_n432));
  INV_X1    g0232(.A(G87), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n254), .A2(new_n433), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n295), .A2(new_n296), .B1(new_n300), .B2(new_n298), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n291), .A2(G1698), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n286), .B(new_n432), .C1(new_n437), .C2(new_n288), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n438), .A2(new_n306), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(G200), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n431), .A2(KEYINPUT17), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n430), .A2(new_n268), .A3(new_n422), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n442), .A2(new_n439), .A3(new_n412), .A4(new_n440), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT17), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n438), .A2(G169), .ZN(new_n447));
  OAI221_X1 g0247(.A(new_n436), .B1(G223), .B2(G1698), .C1(new_n359), .C2(new_n360), .ZN(new_n448));
  INV_X1    g0248(.A(new_n434), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n302), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(G179), .A3(new_n286), .A4(new_n432), .ZN(new_n452));
  AOI221_X4 g0252(.A(new_n446), .B1(new_n447), .B2(new_n452), .C1(new_n442), .C2(new_n412), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n422), .A2(new_n268), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n426), .A2(new_n427), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G68), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n424), .B1(new_n456), .B2(new_n421), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n412), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n447), .A2(new_n452), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT18), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n441), .B(new_n445), .C1(new_n453), .C2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  AND4_X1   g0262(.A1(new_n340), .A2(new_n404), .A3(new_n408), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n205), .A2(G33), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n267), .A2(new_n270), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G97), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n270), .A2(new_n245), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT80), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT80), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n467), .A2(new_n471), .A3(new_n468), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT78), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(new_n263), .B2(G77), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT6), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n248), .B2(new_n249), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n476), .B2(new_n244), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n475), .B1(new_n478), .B2(new_n253), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n243), .B1(new_n426), .B2(new_n427), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT79), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n264), .A2(KEYINPUT78), .A3(new_n202), .ZN(new_n483));
  AOI211_X1 g0283(.A(KEYINPUT79), .B(new_n243), .C1(new_n426), .C2(new_n427), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n473), .B1(new_n485), .B2(new_n267), .ZN(new_n486));
  XNOR2_X1  g0286(.A(KEYINPUT5), .B(G41), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n205), .A2(G45), .A3(G274), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G45), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(G1), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT5), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G41), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n288), .ZN(new_n496));
  INV_X1    g0296(.A(G257), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n489), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G250), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n295), .B2(new_n296), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT4), .ZN(new_n501));
  OAI21_X1  g0301(.A(G1698), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G283), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n254), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(G244), .B1(new_n359), .B2(new_n360), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(new_n501), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n297), .A2(KEYINPUT4), .A3(G244), .A4(new_n298), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n502), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n498), .B1(new_n508), .B2(new_n302), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n314), .ZN(new_n511));
  INV_X1    g0311(.A(G179), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n486), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n318), .A2(new_n270), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n219), .A2(new_n221), .B1(new_n295), .B2(new_n296), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G68), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT19), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n222), .B1(new_n366), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g0319(.A(KEYINPUT81), .B(G87), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n249), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n255), .A2(G97), .A3(new_n259), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n517), .B(new_n522), .C1(new_n523), .C2(KEYINPUT19), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n515), .B1(new_n524), .B2(new_n268), .ZN(new_n525));
  INV_X1    g0325(.A(new_n466), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n318), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n215), .A2(G1698), .ZN(new_n529));
  OAI221_X1 g0329(.A(new_n529), .B1(G238), .B2(G1698), .C1(new_n359), .C2(new_n360), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G116), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n288), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n491), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n288), .A2(new_n533), .A3(G250), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n532), .A2(new_n488), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(G169), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n512), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n528), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n480), .A2(new_n481), .ZN(new_n541));
  INV_X1    g0341(.A(new_n483), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n480), .A2(new_n481), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .A4(new_n479), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n268), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n510), .A2(G200), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n509), .A2(G190), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n545), .A2(new_n473), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n466), .A2(new_n433), .ZN(new_n549));
  AOI211_X1 g0349(.A(new_n515), .B(new_n549), .C1(new_n524), .C2(new_n268), .ZN(new_n550));
  INV_X1    g0350(.A(G200), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n536), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(G190), .B2(new_n536), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  AND4_X1   g0354(.A1(new_n514), .A2(new_n540), .A3(new_n548), .A4(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G257), .B(G1698), .C1(new_n359), .C2(new_n360), .ZN(new_n556));
  OAI211_X1 g0356(.A(G250), .B(new_n298), .C1(new_n359), .C2(new_n360), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G294), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT86), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT86), .A4(new_n558), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n302), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n302), .B1(new_n491), .B2(new_n487), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G264), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n563), .A2(new_n306), .A3(new_n489), .A4(new_n565), .ZN(new_n566));
  OR2_X1    g0366(.A1(new_n566), .A2(KEYINPUT88), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n563), .A2(new_n489), .A3(new_n565), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n551), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(KEYINPUT88), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OR3_X1    g0371(.A1(new_n222), .A2(KEYINPUT23), .A3(G107), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n531), .A2(G20), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n243), .A2(G20), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n573), .B1(KEYINPUT23), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT22), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n516), .B2(G87), .ZN(new_n577));
  AND4_X1   g0377(.A1(new_n576), .A2(new_n222), .A3(new_n297), .A4(G87), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n572), .B(new_n575), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT24), .ZN(new_n580));
  INV_X1    g0380(.A(new_n575), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n222), .A2(new_n297), .A3(G87), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT22), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n516), .A2(new_n576), .A3(G87), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT24), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n572), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n267), .B1(new_n580), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n466), .A2(new_n243), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT85), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(KEYINPUT25), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n270), .A2(new_n591), .A3(G107), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(KEYINPUT25), .ZN(new_n593));
  XNOR2_X1  g0393(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n588), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n571), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n568), .A2(G169), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n563), .A2(G179), .A3(new_n489), .A4(new_n565), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT87), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n579), .A2(KEYINPUT24), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n586), .B1(new_n585), .B2(new_n572), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n268), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n589), .ZN(new_n604));
  INV_X1    g0404(.A(new_n594), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT87), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n597), .A2(new_n607), .A3(new_n598), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n600), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n564), .A2(KEYINPUT82), .A3(G270), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT82), .ZN(new_n611));
  INV_X1    g0411(.A(G270), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(new_n496), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n610), .A2(new_n613), .B1(new_n488), .B2(new_n487), .ZN(new_n614));
  AND2_X1   g0414(.A1(G264), .A2(G1698), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n359), .B2(new_n360), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT83), .ZN(new_n617));
  OAI211_X1 g0417(.A(G257), .B(new_n298), .C1(new_n359), .C2(new_n360), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n414), .A2(G303), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT83), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n620), .B(new_n615), .C1(new_n359), .C2(new_n360), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n617), .A2(new_n618), .A3(new_n619), .A4(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT84), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n622), .A2(new_n623), .A3(new_n302), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n622), .B2(new_n302), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n614), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n526), .A2(G116), .ZN(new_n627));
  INV_X1    g0427(.A(G116), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n271), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n206), .A2(G116), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n267), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n504), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n632), .B(new_n222), .C1(G33), .C2(new_n245), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n631), .A2(KEYINPUT20), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT20), .B1(new_n631), .B2(new_n633), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n627), .B(new_n629), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n626), .A2(G169), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT21), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n636), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n614), .B(G190), .C1(new_n624), .C2(new_n625), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT82), .B1(new_n564), .B2(G270), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n496), .A2(new_n611), .A3(new_n612), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n489), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n622), .A2(new_n623), .A3(new_n302), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n622), .A2(new_n302), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT84), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n644), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n640), .B(new_n641), .C1(new_n648), .C2(new_n551), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G179), .A3(new_n636), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n626), .A2(KEYINPUT21), .A3(new_n636), .A4(G169), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n639), .A2(new_n649), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n555), .A2(new_n596), .A3(new_n609), .A4(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n464), .A2(new_n653), .ZN(G372));
  NAND2_X1  g0454(.A1(new_n335), .A2(new_n385), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n402), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n656), .A2(new_n445), .A3(new_n441), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n453), .A2(new_n460), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n405), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n316), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT89), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n540), .A2(new_n554), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(new_n514), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n663), .B1(new_n665), .B2(KEYINPUT26), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  OAI211_X1 g0467(.A(KEYINPUT89), .B(new_n667), .C1(new_n664), .C2(new_n514), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT90), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n665), .B2(KEYINPUT26), .ZN(new_n670));
  NOR4_X1   g0470(.A1(new_n664), .A2(new_n514), .A3(KEYINPUT90), .A4(new_n667), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n666), .B(new_n668), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n537), .B1(new_n525), .B2(new_n527), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n673), .A2(new_n539), .B1(new_n553), .B2(new_n550), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n596), .A2(new_n674), .A3(new_n514), .A4(new_n548), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n650), .A2(new_n651), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n677), .A2(new_n639), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n606), .A2(new_n599), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n676), .A2(new_n680), .B1(new_n673), .B2(new_n539), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n672), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n662), .B1(new_n464), .B2(new_n683), .ZN(G369));
  NAND2_X1  g0484(.A1(new_n677), .A2(new_n639), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n253), .A2(new_n350), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n205), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G213), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n685), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT91), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n609), .B(new_n596), .C1(new_n595), .C2(new_n693), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n609), .B2(new_n693), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n679), .A2(new_n692), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n692), .A2(new_n636), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n652), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n678), .B2(new_n701), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n697), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n700), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n226), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G1), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n520), .A2(new_n628), .A3(new_n249), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n711), .A2(new_n712), .B1(new_n224), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n678), .A2(KEYINPUT93), .A3(new_n609), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT93), .ZN(new_n717));
  INV_X1    g0517(.A(new_n609), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n718), .B2(new_n685), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n716), .A2(new_n719), .A3(new_n676), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n664), .A2(new_n667), .A3(new_n514), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n665), .A2(KEYINPUT26), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n720), .B(new_n540), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n715), .B1(new_n723), .B2(new_n693), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n692), .B1(new_n672), .B2(new_n681), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n725), .A2(new_n715), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n614), .B(G179), .C1(new_n624), .C2(new_n625), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n509), .A2(new_n565), .A3(new_n563), .A4(new_n536), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT92), .ZN(new_n731));
  OR3_X1    g0531(.A1(new_n728), .A2(new_n729), .A3(new_n727), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n510), .A2(new_n568), .ZN(new_n733));
  OR3_X1    g0533(.A1(new_n532), .A2(new_n488), .A3(new_n535), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n733), .A2(new_n512), .A3(new_n734), .A4(new_n626), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT92), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n736), .B(new_n727), .C1(new_n728), .C2(new_n729), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n731), .A2(new_n732), .A3(new_n735), .A4(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT31), .B1(new_n738), .B2(new_n692), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n609), .A2(new_n639), .A3(new_n677), .A4(new_n649), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n675), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n739), .B1(new_n741), .B2(new_n693), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n732), .A2(new_n735), .A3(new_n730), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n724), .B(new_n726), .C1(G330), .C2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n714), .B1(new_n746), .B2(G1), .ZN(G364));
  AOI21_X1  g0547(.A(new_n711), .B1(G45), .B2(new_n686), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n306), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n512), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n253), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G97), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n222), .A2(new_n512), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n750), .ZN(new_n755));
  INV_X1    g0555(.A(G58), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n306), .A2(new_n551), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n753), .B1(new_n755), .B2(new_n756), .C1(new_n272), .C2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n757), .A2(G20), .A3(new_n512), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n253), .A2(new_n512), .A3(new_n306), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n551), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n297), .B1(new_n520), .B2(new_n760), .C1(new_n763), .C2(new_n243), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n754), .A2(new_n306), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G200), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n759), .B(new_n764), .C1(G77), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n761), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G159), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT32), .Z(new_n770));
  NOR2_X1   g0570(.A1(new_n765), .A2(new_n551), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n767), .B(new_n770), .C1(new_n342), .C2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT95), .ZN(new_n774));
  XOR2_X1   g0574(.A(KEYINPUT33), .B(G317), .Z(new_n775));
  INV_X1    g0575(.A(G322), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n772), .A2(new_n775), .B1(new_n755), .B2(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT96), .Z(new_n778));
  NAND2_X1  g0578(.A1(new_n768), .A2(G329), .ZN(new_n779));
  INV_X1    g0579(.A(G326), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n780), .B2(new_n758), .ZN(new_n781));
  INV_X1    g0581(.A(G294), .ZN(new_n782));
  INV_X1    g0582(.A(new_n752), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n414), .B1(new_n782), .B2(new_n783), .C1(new_n763), .C2(new_n503), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n781), .B(new_n784), .C1(G311), .C2(new_n766), .ZN(new_n785));
  INV_X1    g0585(.A(G303), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n778), .B(new_n785), .C1(new_n786), .C2(new_n760), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n774), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n223), .B1(G20), .B2(new_n314), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n749), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n241), .A2(G45), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n708), .A2(new_n297), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n791), .B(new_n792), .C1(G45), .C2(new_n224), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n708), .A2(new_n414), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G355), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n793), .B(new_n795), .C1(G116), .C2(new_n226), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G13), .A2(G33), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n206), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT94), .ZN(new_n799));
  INV_X1    g0599(.A(new_n789), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n796), .A2(new_n801), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n790), .B(new_n802), .C1(new_n703), .C2(new_n799), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n703), .A2(G330), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n704), .A2(new_n749), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(G396));
  AOI21_X1  g0606(.A(new_n693), .B1(new_n336), .B2(new_n326), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n334), .B1(new_n339), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n327), .A2(new_n332), .A3(new_n333), .A4(new_n693), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n725), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n745), .A2(G330), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n749), .ZN(new_n814));
  INV_X1    g0614(.A(new_n755), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n771), .A2(G150), .B1(new_n815), .B2(G143), .ZN(new_n816));
  INV_X1    g0616(.A(G137), .ZN(new_n817));
  INV_X1    g0617(.A(G159), .ZN(new_n818));
  INV_X1    g0618(.A(new_n766), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n816), .B1(new_n817), .B2(new_n758), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT34), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n297), .B1(new_n783), .B2(new_n756), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n763), .A2(new_n342), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n822), .B(new_n823), .C1(G132), .C2(new_n768), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n821), .B(new_n824), .C1(new_n272), .C2(new_n760), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n760), .A2(new_n243), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n753), .B1(new_n755), .B2(new_n782), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT97), .Z(new_n828));
  AOI22_X1  g0628(.A1(G116), .A2(new_n766), .B1(new_n771), .B2(G283), .ZN(new_n829));
  INV_X1    g0629(.A(new_n758), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n830), .A2(G303), .B1(new_n762), .B2(G87), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n297), .B1(new_n768), .B2(G311), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n828), .A2(new_n829), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n825), .B1(new_n826), .B2(new_n833), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT98), .Z(new_n835));
  AOI21_X1  g0635(.A(new_n749), .B1(new_n835), .B2(new_n789), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n789), .A2(new_n797), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n797), .ZN(new_n839));
  AND4_X1   g0639(.A1(new_n327), .A2(new_n332), .A3(new_n333), .A4(new_n693), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n327), .A2(new_n692), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n406), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n840), .B1(new_n334), .B2(new_n842), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n836), .B1(G77), .B2(new_n838), .C1(new_n839), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n814), .A2(new_n844), .ZN(G384));
  NAND2_X1  g0645(.A1(new_n390), .A2(new_n692), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n385), .A2(new_n402), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(new_n385), .B2(new_n402), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n843), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT103), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n738), .A2(KEYINPUT103), .A3(KEYINPUT31), .A4(new_n692), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n849), .B1(new_n742), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT38), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n462), .A2(new_n431), .A3(new_n690), .ZN(new_n857));
  INV_X1    g0657(.A(new_n690), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n458), .B1(new_n459), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n443), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n860), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n856), .B1(new_n857), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n424), .B1(new_n419), .B2(new_n421), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n412), .B1(new_n454), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n858), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT100), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT100), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n865), .A2(new_n868), .A3(new_n858), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n865), .A2(new_n459), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n443), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT37), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n859), .A2(new_n861), .A3(new_n443), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n461), .A2(KEYINPUT101), .A3(new_n870), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT101), .B1(new_n461), .B2(new_n870), .ZN(new_n877));
  OAI211_X1 g0677(.A(KEYINPUT38), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n863), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n855), .A2(KEYINPUT40), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT40), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n856), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n884), .A2(new_n878), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n385), .A2(new_n402), .A3(new_n846), .ZN(new_n886));
  INV_X1    g0686(.A(new_n846), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n403), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n810), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n852), .A2(new_n853), .ZN(new_n890));
  INV_X1    g0690(.A(new_n739), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n653), .B2(new_n692), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n889), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n882), .B1(new_n885), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT104), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n884), .A2(new_n878), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n855), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(KEYINPUT104), .A3(new_n882), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n881), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n742), .A2(new_n854), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n463), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n900), .B(new_n902), .Z(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(G330), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT102), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n463), .B1(new_n726), .B2(new_n724), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n662), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n905), .B(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n847), .A2(new_n848), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n725), .A2(new_n843), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n910), .B2(new_n809), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n897), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n659), .A2(new_n690), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n885), .A2(KEYINPUT39), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n402), .A2(new_n692), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n879), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n912), .A2(new_n913), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n908), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n205), .B2(new_n686), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n266), .B(new_n253), .C1(new_n478), .C2(KEYINPUT35), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n628), .B(new_n922), .C1(KEYINPUT35), .C2(new_n478), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT99), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT36), .Z(new_n925));
  OAI21_X1  g0725(.A(G77), .B1(new_n756), .B2(new_n342), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n926), .A2(new_n224), .B1(G50), .B2(new_n342), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(G1), .A3(new_n350), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n921), .A2(new_n925), .A3(new_n928), .ZN(G367));
  INV_X1    g0729(.A(G143), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n758), .A2(new_n930), .B1(new_n783), .B2(new_n342), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(G50), .B2(new_n766), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n762), .A2(G77), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n815), .A2(G150), .B1(new_n768), .B2(G137), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n297), .B1(new_n760), .B2(new_n756), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n771), .B2(G159), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n932), .A2(new_n933), .A3(new_n934), .A4(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(G311), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n786), .A2(new_n755), .B1(new_n758), .B2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT108), .Z(new_n940));
  INV_X1    g0740(.A(new_n768), .ZN(new_n941));
  INV_X1    g0741(.A(G317), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n245), .A2(new_n763), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n760), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT46), .B1(new_n944), .B2(G116), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n944), .A2(KEYINPUT46), .A3(G116), .ZN(new_n946));
  NOR4_X1   g0746(.A1(new_n943), .A2(new_n297), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  AOI22_X1  g0747(.A1(G283), .A2(new_n766), .B1(new_n771), .B2(G294), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n940), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n783), .A2(new_n243), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n937), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT47), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n749), .B1(new_n952), .B2(new_n789), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n708), .A2(new_n318), .ZN(new_n954));
  INV_X1    g0754(.A(new_n792), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n801), .B(new_n954), .C1(new_n955), .C2(new_n237), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n674), .B1(new_n550), .B2(new_n693), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(KEYINPUT105), .ZN(new_n958));
  OR3_X1    g0758(.A1(new_n540), .A2(new_n550), .A3(new_n693), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(KEYINPUT105), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n953), .B(new_n956), .C1(new_n961), .C2(new_n799), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n205), .B1(new_n686), .B2(G45), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n486), .A2(new_n692), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n514), .A2(new_n548), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n514), .B2(new_n693), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n700), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT44), .Z(new_n969));
  NAND2_X1  g0769(.A1(new_n700), .A2(new_n967), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT45), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(new_n706), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n704), .B(new_n697), .Z(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(new_n695), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n746), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n746), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n709), .B(KEYINPUT41), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n964), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n698), .A2(new_n967), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT42), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n967), .B(KEYINPUT106), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n718), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n692), .B1(new_n986), .B2(new_n514), .ZN(new_n987));
  NOR3_X1   g0787(.A1(new_n981), .A2(new_n983), .A3(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT107), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n983), .B(new_n990), .C1(new_n981), .C2(new_n987), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n706), .A2(new_n984), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n992), .B(new_n993), .Z(new_n994));
  OAI21_X1  g0794(.A(new_n962), .B1(new_n979), .B2(new_n994), .ZN(G387));
  NOR2_X1   g0795(.A1(new_n746), .A2(new_n975), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n710), .B1(new_n996), .B2(KEYINPUT111), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n997), .B(new_n976), .C1(KEYINPUT111), .C2(new_n996), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n975), .A2(new_n964), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT109), .Z(new_n1000));
  AOI21_X1  g0800(.A(new_n955), .B1(new_n234), .B2(G45), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n712), .B2(new_n794), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n260), .A2(new_n272), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT50), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n342), .A2(new_n202), .ZN(new_n1005));
  NOR4_X1   g0805(.A1(new_n1004), .A2(G45), .A3(new_n712), .A4(new_n1005), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n1002), .A2(new_n1006), .B1(G107), .B2(new_n226), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n749), .B1(new_n1007), .B2(new_n801), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT110), .Z(new_n1009));
  OAI21_X1  g0809(.A(new_n414), .B1(new_n941), .B2(new_n780), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n771), .A2(G311), .B1(new_n815), .B2(G317), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n786), .B2(new_n819), .C1(new_n776), .C2(new_n758), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT48), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n503), .B2(new_n783), .C1(new_n782), .C2(new_n760), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT49), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1010), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n1015), .B2(new_n1014), .C1(new_n628), .C2(new_n763), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n752), .A2(new_n318), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1018), .B(new_n297), .C1(new_n202), .C2(new_n760), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G68), .B2(new_n766), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n771), .A2(new_n260), .B1(G97), .B2(new_n762), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n815), .A2(G50), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n830), .A2(G159), .B1(new_n768), .B2(G150), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n1017), .A2(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1009), .B1(new_n697), .B2(new_n799), .C1(new_n1025), .C2(new_n800), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n998), .A2(new_n1000), .A3(new_n1026), .ZN(G393));
  OR2_X1    g0827(.A1(new_n973), .A2(new_n976), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n973), .A2(new_n976), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1028), .A2(new_n709), .A3(new_n1029), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n973), .A2(new_n963), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G87), .A2(new_n762), .B1(new_n768), .B2(G143), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n297), .B1(new_n760), .B2(new_n342), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G77), .B2(new_n752), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1032), .B(new_n1034), .C1(new_n772), .C2(new_n272), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n262), .A2(new_n758), .B1(new_n755), .B2(new_n818), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT51), .Z(new_n1037));
  AOI211_X1 g0837(.A(new_n1035), .B(new_n1037), .C1(new_n260), .C2(new_n766), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n762), .A2(G107), .B1(G116), .B2(new_n752), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n414), .B1(new_n760), .B2(new_n503), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n768), .B2(G322), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1039), .B(new_n1041), .C1(new_n772), .C2(new_n786), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n938), .A2(new_n755), .B1(new_n758), .B2(new_n942), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT52), .Z(new_n1044));
  AOI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(G294), .C2(new_n766), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n789), .B1(new_n1038), .B2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n792), .A2(new_n251), .B1(G97), .B2(new_n708), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n749), .B1(new_n1047), .B2(new_n801), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT112), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1046), .B(new_n1049), .C1(new_n985), .C2(new_n799), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1030), .A2(new_n1031), .A3(new_n1050), .ZN(G390));
  AND2_X1   g0851(.A1(new_n843), .A2(G330), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n745), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1053), .A2(new_n909), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n909), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n901), .B2(new_n1052), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n723), .A2(new_n693), .A3(new_n808), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1058), .A2(new_n809), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1053), .A2(new_n909), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n901), .A2(new_n1055), .A3(new_n1052), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n910), .A2(new_n809), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1057), .A2(new_n1059), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n463), .A2(G330), .A3(new_n901), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n906), .A2(new_n1065), .A3(new_n662), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n914), .A2(new_n917), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n911), .B2(new_n915), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n915), .B1(new_n863), .B2(new_n878), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1059), .B2(new_n909), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1069), .A2(new_n1071), .A3(new_n1054), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1061), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1067), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n709), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1067), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1068), .A2(new_n797), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n414), .B1(new_n433), .B2(new_n760), .C1(new_n819), .C2(new_n245), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n823), .B(new_n1081), .C1(G107), .C2(new_n771), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n830), .A2(G283), .B1(new_n768), .B2(G294), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n628), .B2(new_n755), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G77), .B2(new_n752), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n414), .B1(new_n752), .B2(G159), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT54), .B(G143), .Z(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1087), .B1(new_n772), .B2(new_n817), .C1(new_n819), .C2(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n815), .A2(G132), .B1(new_n768), .B2(G125), .ZN(new_n1091));
  INV_X1    g0891(.A(G128), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1091), .B1(new_n272), .B2(new_n763), .C1(new_n1092), .C2(new_n758), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n944), .A2(G150), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT53), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1086), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1097), .A2(new_n789), .B1(new_n410), .B2(new_n837), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1080), .A2(new_n748), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n1077), .B2(new_n963), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1079), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(G378));
  NAND3_X1  g0902(.A1(new_n912), .A2(new_n913), .A3(new_n918), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(KEYINPUT114), .B(KEYINPUT56), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n317), .A2(KEYINPUT55), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT55), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n309), .A2(new_n1107), .A3(new_n313), .A4(new_n316), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n277), .A2(new_n858), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1109), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1105), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1109), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n1104), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT115), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n900), .B2(G330), .ZN(new_n1119));
  AOI21_X1  g0919(.A(KEYINPUT104), .B1(new_n898), .B2(new_n882), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n895), .B(KEYINPUT40), .C1(new_n855), .C2(new_n897), .ZN(new_n1121));
  OAI211_X1 g0921(.A(G330), .B(new_n880), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1112), .A2(new_n1117), .A3(KEYINPUT115), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(new_n1118), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1103), .B1(new_n1119), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT116), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT115), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1112), .A2(new_n1117), .A3(KEYINPUT115), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n900), .A2(G330), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1122), .A2(new_n1130), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n919), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1126), .A2(new_n1127), .A3(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(KEYINPUT116), .B(new_n1103), .C1(new_n1119), .C2(new_n1125), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1066), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1075), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT57), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(KEYINPUT119), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1135), .A2(KEYINPUT117), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT117), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1133), .A2(new_n1134), .A3(new_n919), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT118), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1126), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n919), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(KEYINPUT118), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1147), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1152), .A2(KEYINPUT57), .A3(new_n1139), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT119), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1140), .A2(new_n1154), .A3(new_n1141), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1143), .A2(new_n709), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1136), .A2(new_n964), .A3(new_n1137), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n762), .A2(G58), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1158), .B(new_n287), .C1(new_n202), .C2(new_n760), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n297), .B(new_n1159), .C1(G283), .C2(new_n768), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT113), .Z(new_n1161));
  OAI22_X1  g0961(.A1(new_n758), .A2(new_n628), .B1(new_n783), .B2(new_n342), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n772), .A2(new_n245), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n318), .C2(new_n766), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1161), .B(new_n1164), .C1(new_n243), .C2(new_n755), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT58), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n272), .B1(new_n359), .B2(G41), .ZN(new_n1167));
  INV_X1    g0967(.A(G132), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n1168), .A2(new_n772), .B1(new_n819), .B2(new_n817), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n830), .A2(G125), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n1092), .B2(new_n755), .C1(new_n760), .C2(new_n1089), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(G150), .C2(new_n752), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT59), .ZN(new_n1173));
  AOI21_X1  g0973(.A(G41), .B1(new_n768), .B2(G124), .ZN(new_n1174));
  AOI21_X1  g0974(.A(G33), .B1(new_n762), .B2(G159), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1166), .A2(new_n1167), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n749), .B1(new_n1177), .B2(new_n789), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(G50), .B2(new_n838), .C1(new_n1128), .C2(new_n839), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1157), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1156), .A2(new_n1181), .ZN(G375));
  AOI22_X1  g0982(.A1(new_n830), .A2(G294), .B1(new_n768), .B2(G303), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n771), .A2(G116), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n297), .B1(new_n944), .B2(G97), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n933), .A4(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1018), .B1(new_n755), .B2(new_n503), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT121), .Z(new_n1188));
  AOI211_X1 g0988(.A(new_n1186), .B(new_n1188), .C1(G107), .C2(new_n766), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n815), .A2(G137), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1158), .B1(new_n272), .B2(new_n783), .C1(new_n819), .C2(new_n262), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n297), .B1(new_n818), .B2(new_n760), .C1(new_n772), .C2(new_n1089), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n941), .A2(new_n1092), .B1(new_n758), .B2(new_n1168), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1189), .B1(new_n1190), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1195), .A2(new_n800), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n748), .B1(G68), .B2(new_n838), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT120), .Z(new_n1198));
  AOI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(new_n909), .C2(new_n797), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1064), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n1200), .B2(new_n964), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n978), .B1(new_n1200), .B2(new_n1138), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1201), .B1(new_n1202), .B2(new_n1067), .ZN(G381));
  OR4_X1    g1003(.A1(G384), .A2(G375), .A3(G378), .A4(G381), .ZN(new_n1204));
  OR2_X1    g1004(.A1(G387), .A2(G390), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1204), .A2(G396), .A3(G393), .A4(new_n1205), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT122), .Z(G407));
  AND3_X1   g1007(.A1(new_n1140), .A2(new_n1154), .A3(new_n1141), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1154), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1139), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1150), .B(new_n1148), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n1147), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n710), .B1(new_n1213), .B2(KEYINPUT57), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1180), .B1(new_n1210), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(new_n691), .A3(new_n1101), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(G407), .A2(G213), .A3(new_n1216), .ZN(G409));
  XNOR2_X1  g1017(.A(G393), .B(G396), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G387), .A2(G390), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT124), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(G387), .B2(G390), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1219), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1205), .A2(new_n1220), .A3(new_n1222), .A4(new_n1218), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT62), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1200), .A2(new_n1138), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT60), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(new_n709), .A3(new_n1078), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1228), .A2(KEYINPUT60), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1201), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(G384), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(G213), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(G343), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(G2897), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n978), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1140), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n964), .B2(new_n1152), .ZN(new_n1246));
  AOI21_X1  g1046(.A(G378), .B1(new_n1246), .B2(new_n1179), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT123), .B1(new_n1215), .B2(G378), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1156), .A2(KEYINPUT123), .A3(G378), .A4(new_n1181), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1248), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1238), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1243), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1156), .A2(G378), .A3(new_n1181), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT123), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1247), .B1(new_n1257), .B2(new_n1250), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1236), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n1238), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1227), .B1(new_n1254), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1252), .A2(new_n1236), .A3(new_n1253), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT61), .B1(new_n1262), .B2(KEYINPUT62), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1226), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1242), .B1(new_n1258), .B2(new_n1238), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1257), .A2(new_n1250), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1238), .B1(new_n1266), .B2(new_n1248), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1265), .A2(KEYINPUT63), .B1(new_n1267), .B2(new_n1236), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1252), .A2(KEYINPUT63), .A3(new_n1236), .A4(new_n1253), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1226), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1268), .A2(new_n1270), .A3(KEYINPUT61), .ZN(new_n1271));
  OAI21_X1  g1071(.A(KEYINPUT125), .B1(new_n1264), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1226), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1260), .B2(new_n1227), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT62), .B1(new_n1262), .B2(new_n1265), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1273), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1262), .B1(new_n1254), .B2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1279), .A2(new_n1274), .A3(new_n1226), .A4(new_n1269), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT125), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1277), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1272), .A2(new_n1282), .ZN(G405));
  INV_X1    g1083(.A(KEYINPUT126), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1215), .B2(G378), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(G375), .A2(KEYINPUT126), .A3(new_n1101), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1266), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1287), .B(new_n1236), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1288), .B(new_n1273), .ZN(G402));
endmodule


