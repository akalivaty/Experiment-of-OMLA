

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U558 ( .A1(n773), .A2(n772), .ZN(n775) );
  XOR2_X1 U559 ( .A(n542), .B(KEYINPUT87), .Z(n523) );
  OR2_X1 U560 ( .A1(KEYINPUT103), .A2(n755), .ZN(n524) );
  NOR2_X1 U561 ( .A1(n734), .A2(n687), .ZN(n689) );
  NOR2_X1 U562 ( .A1(n973), .A2(n692), .ZN(n694) );
  INV_X1 U563 ( .A(KEYINPUT28), .ZN(n709) );
  INV_X1 U564 ( .A(n982), .ZN(n752) );
  OR2_X1 U565 ( .A1(n771), .A2(n752), .ZN(n753) );
  OR2_X1 U566 ( .A1(n732), .A2(n731), .ZN(n749) );
  NAND2_X1 U567 ( .A1(n686), .A2(n797), .ZN(n734) );
  INV_X1 U568 ( .A(KEYINPUT104), .ZN(n774) );
  INV_X1 U569 ( .A(G2105), .ZN(n536) );
  AND2_X1 U570 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U571 ( .A(n537), .B(KEYINPUT64), .ZN(n895) );
  NOR2_X1 U572 ( .A1(G651), .A2(n627), .ZN(n653) );
  NAND2_X1 U573 ( .A1(n523), .A2(n544), .ZN(n545) );
  XOR2_X1 U574 ( .A(G543), .B(KEYINPUT0), .Z(n627) );
  INV_X1 U575 ( .A(G651), .ZN(n531) );
  NOR2_X1 U576 ( .A1(n627), .A2(n531), .ZN(n649) );
  NAND2_X1 U577 ( .A1(n649), .A2(G77), .ZN(n525) );
  XNOR2_X1 U578 ( .A(n525), .B(KEYINPUT68), .ZN(n527) );
  NOR2_X1 U579 ( .A1(G543), .A2(G651), .ZN(n645) );
  NAND2_X1 U580 ( .A1(G90), .A2(n645), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U582 ( .A(n528), .B(KEYINPUT9), .ZN(n530) );
  NAND2_X1 U583 ( .A1(G52), .A2(n653), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n535) );
  NOR2_X1 U585 ( .A1(G543), .A2(n531), .ZN(n532) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n532), .Z(n646) );
  NAND2_X1 U587 ( .A1(G64), .A2(n646), .ZN(n533) );
  XNOR2_X1 U588 ( .A(KEYINPUT67), .B(n533), .ZN(n534) );
  NOR2_X1 U589 ( .A1(n535), .A2(n534), .ZN(G171) );
  AND2_X1 U590 ( .A1(G452), .A2(G94), .ZN(G173) );
  AND2_X1 U591 ( .A1(n536), .A2(G2104), .ZN(n898) );
  NAND2_X1 U592 ( .A1(G102), .A2(n898), .ZN(n539) );
  NOR2_X1 U593 ( .A1(n536), .A2(G2104), .ZN(n537) );
  NAND2_X1 U594 ( .A1(G126), .A2(n895), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n546) );
  XNOR2_X1 U596 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n541) );
  NOR2_X1 U597 ( .A1(G2104), .A2(G2105), .ZN(n540) );
  XNOR2_X2 U598 ( .A(n541), .B(n540), .ZN(n899) );
  NAND2_X1 U599 ( .A1(G138), .A2(n899), .ZN(n542) );
  AND2_X1 U600 ( .A1(G2104), .A2(G2105), .ZN(n894) );
  NAND2_X1 U601 ( .A1(G114), .A2(n894), .ZN(n543) );
  XNOR2_X1 U602 ( .A(n543), .B(KEYINPUT86), .ZN(n544) );
  NOR2_X1 U603 ( .A1(n546), .A2(n545), .ZN(G164) );
  INV_X1 U604 ( .A(G57), .ZN(G237) );
  INV_X1 U605 ( .A(G82), .ZN(G220) );
  NAND2_X1 U606 ( .A1(n894), .A2(G113), .ZN(n549) );
  NAND2_X1 U607 ( .A1(G101), .A2(n898), .ZN(n547) );
  XOR2_X1 U608 ( .A(KEYINPUT23), .B(n547), .Z(n548) );
  NAND2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G137), .A2(n899), .ZN(n551) );
  NAND2_X1 U611 ( .A1(G125), .A2(n895), .ZN(n550) );
  NAND2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U613 ( .A1(n553), .A2(n552), .ZN(G160) );
  NAND2_X1 U614 ( .A1(G51), .A2(n653), .ZN(n555) );
  NAND2_X1 U615 ( .A1(G63), .A2(n646), .ZN(n554) );
  NAND2_X1 U616 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U617 ( .A(KEYINPUT6), .B(n556), .ZN(n563) );
  NAND2_X1 U618 ( .A1(n645), .A2(G89), .ZN(n557) );
  XNOR2_X1 U619 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U620 ( .A1(G76), .A2(n649), .ZN(n558) );
  NAND2_X1 U621 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT74), .B(n560), .Z(n561) );
  XNOR2_X1 U623 ( .A(KEYINPUT5), .B(n561), .ZN(n562) );
  NOR2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U625 ( .A(KEYINPUT7), .B(n564), .Z(G168) );
  XOR2_X1 U626 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U627 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U629 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n567) );
  INV_X1 U630 ( .A(G223), .ZN(n831) );
  NAND2_X1 U631 ( .A1(G567), .A2(n831), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G234) );
  NAND2_X1 U633 ( .A1(n645), .A2(G81), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G68), .A2(n649), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U637 ( .A(KEYINPUT13), .B(n571), .Z(n574) );
  NAND2_X1 U638 ( .A1(n646), .A2(G56), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT14), .B(n572), .Z(n573) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n653), .A2(G43), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n973) );
  INV_X1 U643 ( .A(G860), .ZN(n599) );
  OR2_X1 U644 ( .A1(n973), .A2(n599), .ZN(G153) );
  INV_X1 U645 ( .A(G868), .ZN(n667) );
  NOR2_X1 U646 ( .A1(n667), .A2(G171), .ZN(n577) );
  XNOR2_X1 U647 ( .A(n577), .B(KEYINPUT71), .ZN(n588) );
  NAND2_X1 U648 ( .A1(G79), .A2(n649), .ZN(n579) );
  NAND2_X1 U649 ( .A1(G54), .A2(n653), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U651 ( .A(KEYINPUT73), .B(n580), .Z(n583) );
  NAND2_X1 U652 ( .A1(G92), .A2(n645), .ZN(n581) );
  XOR2_X1 U653 ( .A(KEYINPUT72), .B(n581), .Z(n582) );
  NOR2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n646), .A2(G66), .ZN(n584) );
  NAND2_X1 U656 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U657 ( .A(KEYINPUT15), .B(n586), .ZN(n975) );
  OR2_X1 U658 ( .A1(G868), .A2(n975), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n588), .A2(n587), .ZN(G284) );
  NAND2_X1 U660 ( .A1(G53), .A2(n653), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G65), .A2(n646), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G78), .A2(n649), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G91), .A2(n645), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n981) );
  INV_X1 U667 ( .A(n981), .ZN(G299) );
  NOR2_X1 U668 ( .A1(G286), .A2(n667), .ZN(n595) );
  XOR2_X1 U669 ( .A(KEYINPUT75), .B(n595), .Z(n597) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U672 ( .A(KEYINPUT76), .B(n598), .ZN(G297) );
  NAND2_X1 U673 ( .A1(n599), .A2(G559), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n600), .A2(n975), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n601), .B(KEYINPUT16), .ZN(n602) );
  XOR2_X1 U676 ( .A(KEYINPUT77), .B(n602), .Z(G148) );
  NOR2_X1 U677 ( .A1(G868), .A2(n973), .ZN(n605) );
  NAND2_X1 U678 ( .A1(G868), .A2(n975), .ZN(n603) );
  NOR2_X1 U679 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U680 ( .A1(n605), .A2(n604), .ZN(G282) );
  XNOR2_X1 U681 ( .A(G2100), .B(KEYINPUT79), .ZN(n615) );
  NAND2_X1 U682 ( .A1(G99), .A2(n898), .ZN(n607) );
  NAND2_X1 U683 ( .A1(G111), .A2(n894), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n895), .A2(G123), .ZN(n608) );
  XNOR2_X1 U686 ( .A(n608), .B(KEYINPUT18), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n899), .A2(G135), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n922) );
  XNOR2_X1 U690 ( .A(n922), .B(G2096), .ZN(n613) );
  XNOR2_X1 U691 ( .A(n613), .B(KEYINPUT78), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U693 ( .A1(n975), .A2(G559), .ZN(n664) );
  XNOR2_X1 U694 ( .A(n973), .B(n664), .ZN(n616) );
  NOR2_X1 U695 ( .A1(n616), .A2(G860), .ZN(n623) );
  NAND2_X1 U696 ( .A1(G93), .A2(n645), .ZN(n618) );
  NAND2_X1 U697 ( .A1(G67), .A2(n646), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U699 ( .A1(G80), .A2(n649), .ZN(n620) );
  NAND2_X1 U700 ( .A1(G55), .A2(n653), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n621) );
  OR2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n666) );
  XOR2_X1 U703 ( .A(n623), .B(n666), .Z(G145) );
  NAND2_X1 U704 ( .A1(G49), .A2(n653), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U707 ( .A1(n646), .A2(n626), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n627), .A2(G87), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U710 ( .A1(G62), .A2(n646), .ZN(n630) );
  XOR2_X1 U711 ( .A(KEYINPUT80), .B(n630), .Z(n635) );
  NAND2_X1 U712 ( .A1(G75), .A2(n649), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G88), .A2(n645), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U715 ( .A(KEYINPUT81), .B(n633), .Z(n634) );
  NOR2_X1 U716 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n653), .A2(G50), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n637), .A2(n636), .ZN(G303) );
  INV_X1 U719 ( .A(G303), .ZN(G166) );
  NAND2_X1 U720 ( .A1(G86), .A2(n645), .ZN(n639) );
  NAND2_X1 U721 ( .A1(G61), .A2(n646), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n649), .A2(G73), .ZN(n640) );
  XOR2_X1 U724 ( .A(KEYINPUT2), .B(n640), .Z(n641) );
  NOR2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n653), .A2(G48), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n644), .A2(n643), .ZN(G305) );
  NAND2_X1 U728 ( .A1(G85), .A2(n645), .ZN(n648) );
  NAND2_X1 U729 ( .A1(G60), .A2(n646), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U731 ( .A1(n649), .A2(G72), .ZN(n650) );
  XOR2_X1 U732 ( .A(KEYINPUT66), .B(n650), .Z(n651) );
  NOR2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n653), .A2(G47), .ZN(n654) );
  NAND2_X1 U735 ( .A1(n655), .A2(n654), .ZN(G290) );
  XNOR2_X1 U736 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n657) );
  XNOR2_X1 U737 ( .A(G288), .B(KEYINPUT19), .ZN(n656) );
  XNOR2_X1 U738 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n658), .B(n666), .ZN(n660) );
  XNOR2_X1 U740 ( .A(n981), .B(G166), .ZN(n659) );
  XNOR2_X1 U741 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n661), .B(G305), .ZN(n662) );
  XNOR2_X1 U743 ( .A(n662), .B(G290), .ZN(n663) );
  XNOR2_X1 U744 ( .A(n663), .B(n973), .ZN(n848) );
  XNOR2_X1 U745 ( .A(n664), .B(n848), .ZN(n665) );
  NAND2_X1 U746 ( .A1(n665), .A2(G868), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U748 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U753 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U755 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U756 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U757 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U758 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U759 ( .A1(G96), .A2(n676), .ZN(n835) );
  AND2_X1 U760 ( .A1(G2106), .A2(n835), .ZN(n681) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n677) );
  NOR2_X1 U762 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U763 ( .A1(G108), .A2(n678), .ZN(n836) );
  NAND2_X1 U764 ( .A1(G567), .A2(n836), .ZN(n679) );
  XOR2_X1 U765 ( .A(KEYINPUT84), .B(n679), .Z(n680) );
  NOR2_X1 U766 ( .A1(n681), .A2(n680), .ZN(G319) );
  INV_X1 U767 ( .A(G319), .ZN(n914) );
  NAND2_X1 U768 ( .A1(G483), .A2(G661), .ZN(n682) );
  NOR2_X1 U769 ( .A1(n914), .A2(n682), .ZN(n834) );
  NAND2_X1 U770 ( .A1(G36), .A2(n834), .ZN(n683) );
  XOR2_X1 U771 ( .A(KEYINPUT85), .B(n683), .Z(G176) );
  NOR2_X1 U772 ( .A1(G1971), .A2(G303), .ZN(n751) );
  NOR2_X1 U773 ( .A1(G1976), .A2(G288), .ZN(n684) );
  XOR2_X1 U774 ( .A(KEYINPUT102), .B(n684), .Z(n988) );
  NAND2_X1 U775 ( .A1(G160), .A2(G40), .ZN(n796) );
  INV_X1 U776 ( .A(n796), .ZN(n686) );
  NOR2_X1 U777 ( .A1(G164), .A2(G1384), .ZN(n797) );
  INV_X1 U778 ( .A(G1996), .ZN(n687) );
  INV_X1 U779 ( .A(KEYINPUT26), .ZN(n688) );
  XNOR2_X1 U780 ( .A(n689), .B(n688), .ZN(n691) );
  NAND2_X1 U781 ( .A1(n734), .A2(G1341), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U783 ( .A1(n975), .A2(n694), .ZN(n693) );
  XOR2_X1 U784 ( .A(n693), .B(KEYINPUT98), .Z(n700) );
  NAND2_X1 U785 ( .A1(n975), .A2(n694), .ZN(n698) );
  XNOR2_X1 U786 ( .A(n734), .B(KEYINPUT96), .ZN(n701) );
  INV_X1 U787 ( .A(n701), .ZN(n715) );
  NAND2_X1 U788 ( .A1(G2067), .A2(n715), .ZN(n696) );
  NAND2_X1 U789 ( .A1(G1348), .A2(n734), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n707) );
  NAND2_X1 U793 ( .A1(n701), .A2(G1956), .ZN(n702) );
  XNOR2_X1 U794 ( .A(KEYINPUT97), .B(n702), .ZN(n705) );
  NAND2_X1 U795 ( .A1(G2072), .A2(n715), .ZN(n703) );
  XNOR2_X1 U796 ( .A(n703), .B(KEYINPUT27), .ZN(n704) );
  NOR2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n981), .A2(n708), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n712) );
  NOR2_X1 U800 ( .A1(n981), .A2(n708), .ZN(n710) );
  XNOR2_X1 U801 ( .A(n710), .B(n709), .ZN(n711) );
  NAND2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n714) );
  XNOR2_X1 U803 ( .A(KEYINPUT29), .B(KEYINPUT99), .ZN(n713) );
  XNOR2_X1 U804 ( .A(n714), .B(n713), .ZN(n719) );
  XNOR2_X1 U805 ( .A(KEYINPUT25), .B(G2078), .ZN(n950) );
  NAND2_X1 U806 ( .A1(n950), .A2(n715), .ZN(n717) );
  XNOR2_X1 U807 ( .A(G1961), .B(KEYINPUT95), .ZN(n1017) );
  NAND2_X1 U808 ( .A1(n1017), .A2(n734), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n724) );
  NAND2_X1 U810 ( .A1(n724), .A2(G171), .ZN(n718) );
  NAND2_X1 U811 ( .A1(n719), .A2(n718), .ZN(n742) );
  NAND2_X1 U812 ( .A1(G8), .A2(n734), .ZN(n771) );
  NOR2_X1 U813 ( .A1(G1966), .A2(n771), .ZN(n729) );
  NOR2_X1 U814 ( .A1(G2084), .A2(n734), .ZN(n728) );
  NOR2_X1 U815 ( .A1(n729), .A2(n728), .ZN(n720) );
  NAND2_X1 U816 ( .A1(G8), .A2(n720), .ZN(n722) );
  XNOR2_X1 U817 ( .A(KEYINPUT100), .B(KEYINPUT30), .ZN(n721) );
  XNOR2_X1 U818 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U819 ( .A1(G168), .A2(n723), .ZN(n726) );
  NOR2_X1 U820 ( .A1(G171), .A2(n724), .ZN(n725) );
  NOR2_X1 U821 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U822 ( .A(KEYINPUT31), .B(n727), .Z(n740) );
  AND2_X1 U823 ( .A1(n742), .A2(n740), .ZN(n732) );
  AND2_X1 U824 ( .A1(G8), .A2(n728), .ZN(n730) );
  OR2_X1 U825 ( .A1(n730), .A2(n729), .ZN(n731) );
  INV_X1 U826 ( .A(G8), .ZN(n739) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n771), .ZN(n733) );
  XNOR2_X1 U828 ( .A(KEYINPUT101), .B(n733), .ZN(n737) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n734), .ZN(n735) );
  NOR2_X1 U830 ( .A1(G166), .A2(n735), .ZN(n736) );
  NAND2_X1 U831 ( .A1(n737), .A2(n736), .ZN(n738) );
  OR2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n743) );
  AND2_X1 U833 ( .A1(n740), .A2(n743), .ZN(n741) );
  NAND2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n746) );
  INV_X1 U835 ( .A(n743), .ZN(n744) );
  OR2_X1 U836 ( .A1(n744), .A2(G286), .ZN(n745) );
  NAND2_X1 U837 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U838 ( .A(n747), .B(KEYINPUT32), .ZN(n748) );
  NAND2_X1 U839 ( .A1(n749), .A2(n748), .ZN(n765) );
  NAND2_X1 U840 ( .A1(n988), .A2(n765), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n751), .A2(n750), .ZN(n754) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n982) );
  OR2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n755) );
  INV_X1 U844 ( .A(KEYINPUT33), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n524), .A2(n756), .ZN(n762) );
  XNOR2_X1 U846 ( .A(n988), .B(KEYINPUT103), .ZN(n757) );
  NAND2_X1 U847 ( .A1(n757), .A2(KEYINPUT33), .ZN(n758) );
  NOR2_X1 U848 ( .A1(n771), .A2(n758), .ZN(n760) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n969) );
  INV_X1 U850 ( .A(n969), .ZN(n759) );
  NOR2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n768) );
  NOR2_X1 U853 ( .A1(G2090), .A2(G303), .ZN(n763) );
  NAND2_X1 U854 ( .A1(G8), .A2(n763), .ZN(n764) );
  NAND2_X1 U855 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n766), .A2(n771), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n773) );
  NOR2_X1 U858 ( .A1(G1981), .A2(G305), .ZN(n769) );
  XOR2_X1 U859 ( .A(n769), .B(KEYINPUT24), .Z(n770) );
  NOR2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U861 ( .A(n775), .B(n774), .ZN(n814) );
  NAND2_X1 U862 ( .A1(G95), .A2(n898), .ZN(n777) );
  NAND2_X1 U863 ( .A1(G131), .A2(n899), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n782) );
  NAND2_X1 U865 ( .A1(G107), .A2(n894), .ZN(n779) );
  NAND2_X1 U866 ( .A1(G119), .A2(n895), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U868 ( .A(KEYINPUT89), .B(n780), .Z(n781) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U870 ( .A(KEYINPUT90), .B(n783), .Z(n910) );
  NAND2_X1 U871 ( .A1(G1991), .A2(n910), .ZN(n784) );
  XNOR2_X1 U872 ( .A(n784), .B(KEYINPUT91), .ZN(n795) );
  XOR2_X1 U873 ( .A(KEYINPUT92), .B(KEYINPUT38), .Z(n786) );
  NAND2_X1 U874 ( .A1(G105), .A2(n898), .ZN(n785) );
  XNOR2_X1 U875 ( .A(n786), .B(n785), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G117), .A2(n894), .ZN(n788) );
  NAND2_X1 U877 ( .A1(G129), .A2(n895), .ZN(n787) );
  NAND2_X1 U878 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U880 ( .A(KEYINPUT93), .B(n791), .Z(n793) );
  NAND2_X1 U881 ( .A1(n899), .A2(G141), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n905) );
  AND2_X1 U883 ( .A1(G1996), .A2(n905), .ZN(n794) );
  NOR2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n928) );
  NOR2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n826) );
  XOR2_X1 U886 ( .A(KEYINPUT94), .B(n826), .Z(n798) );
  NOR2_X1 U887 ( .A1(n928), .A2(n798), .ZN(n817) );
  INV_X1 U888 ( .A(n817), .ZN(n812) );
  XNOR2_X1 U889 ( .A(G1986), .B(G290), .ZN(n990) );
  AND2_X1 U890 ( .A1(n826), .A2(n990), .ZN(n810) );
  XOR2_X1 U891 ( .A(G2067), .B(KEYINPUT37), .Z(n822) );
  XNOR2_X1 U892 ( .A(KEYINPUT34), .B(KEYINPUT88), .ZN(n802) );
  NAND2_X1 U893 ( .A1(G104), .A2(n898), .ZN(n800) );
  NAND2_X1 U894 ( .A1(G140), .A2(n899), .ZN(n799) );
  NAND2_X1 U895 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U896 ( .A(n802), .B(n801), .ZN(n807) );
  NAND2_X1 U897 ( .A1(G116), .A2(n894), .ZN(n804) );
  NAND2_X1 U898 ( .A1(G128), .A2(n895), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U900 ( .A(KEYINPUT35), .B(n805), .Z(n806) );
  NOR2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U902 ( .A(KEYINPUT36), .B(n808), .Z(n909) );
  AND2_X1 U903 ( .A1(n822), .A2(n909), .ZN(n924) );
  NAND2_X1 U904 ( .A1(n826), .A2(n924), .ZN(n820) );
  INV_X1 U905 ( .A(n820), .ZN(n809) );
  NOR2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n829) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n905), .ZN(n931) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n815) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n910), .ZN(n923) );
  NOR2_X1 U911 ( .A1(n815), .A2(n923), .ZN(n816) );
  NOR2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U913 ( .A1(n931), .A2(n818), .ZN(n819) );
  XNOR2_X1 U914 ( .A(n819), .B(KEYINPUT39), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n824) );
  NOR2_X1 U916 ( .A1(n909), .A2(n822), .ZN(n823) );
  XNOR2_X1 U917 ( .A(n823), .B(KEYINPUT105), .ZN(n936) );
  NAND2_X1 U918 ( .A1(n824), .A2(n936), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U920 ( .A(n827), .B(KEYINPUT106), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U922 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U925 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n834), .A2(n833), .ZN(G188) );
  NOR2_X1 U929 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U930 ( .A(n837), .B(KEYINPUT108), .ZN(G325) );
  XNOR2_X1 U931 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U935 ( .A(G1348), .B(G2454), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n838), .B(G2430), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n839), .B(G1341), .ZN(n845) );
  XOR2_X1 U938 ( .A(G2443), .B(G2427), .Z(n841) );
  XNOR2_X1 U939 ( .A(G2438), .B(G2446), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n843) );
  XOR2_X1 U941 ( .A(G2451), .B(G2435), .Z(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  NAND2_X1 U944 ( .A1(n846), .A2(G14), .ZN(n847) );
  XNOR2_X1 U945 ( .A(KEYINPUT107), .B(n847), .ZN(G401) );
  XOR2_X1 U946 ( .A(n848), .B(G286), .Z(n850) );
  XNOR2_X1 U947 ( .A(n975), .B(G171), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  NOR2_X1 U949 ( .A1(G37), .A2(n851), .ZN(G397) );
  XOR2_X1 U950 ( .A(KEYINPUT112), .B(G2678), .Z(n853) );
  XNOR2_X1 U951 ( .A(KEYINPUT43), .B(G2100), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U953 ( .A(n854), .B(KEYINPUT42), .Z(n856) );
  XNOR2_X1 U954 ( .A(G2072), .B(G2078), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U956 ( .A(G2096), .B(G2090), .Z(n858) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2084), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U959 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U960 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(G227) );
  XOR2_X1 U962 ( .A(G1986), .B(G1976), .Z(n864) );
  XNOR2_X1 U963 ( .A(G1961), .B(G1971), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U965 ( .A(G1991), .B(G1981), .Z(n866) );
  XNOR2_X1 U966 ( .A(G1966), .B(G1996), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U968 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U969 ( .A(G2474), .B(KEYINPUT41), .ZN(n869) );
  XNOR2_X1 U970 ( .A(n870), .B(n869), .ZN(n872) );
  XOR2_X1 U971 ( .A(G1956), .B(KEYINPUT113), .Z(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(G229) );
  NAND2_X1 U973 ( .A1(G100), .A2(n898), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G112), .A2(n894), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n880) );
  NAND2_X1 U976 ( .A1(n895), .A2(G124), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n875), .B(KEYINPUT114), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n876), .B(KEYINPUT44), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G136), .A2(n899), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U981 ( .A1(n880), .A2(n879), .ZN(G162) );
  XOR2_X1 U982 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n882) );
  XNOR2_X1 U983 ( .A(G164), .B(n922), .ZN(n881) );
  XNOR2_X1 U984 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U985 ( .A(n883), .B(G162), .Z(n893) );
  NAND2_X1 U986 ( .A1(G103), .A2(n898), .ZN(n885) );
  NAND2_X1 U987 ( .A1(G139), .A2(n899), .ZN(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U989 ( .A(KEYINPUT115), .B(n886), .Z(n891) );
  NAND2_X1 U990 ( .A1(G115), .A2(n894), .ZN(n888) );
  NAND2_X1 U991 ( .A1(G127), .A2(n895), .ZN(n887) );
  NAND2_X1 U992 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U994 ( .A1(n891), .A2(n890), .ZN(n938) );
  XNOR2_X1 U995 ( .A(G160), .B(n938), .ZN(n892) );
  XNOR2_X1 U996 ( .A(n893), .B(n892), .ZN(n908) );
  NAND2_X1 U997 ( .A1(G118), .A2(n894), .ZN(n897) );
  NAND2_X1 U998 ( .A1(G130), .A2(n895), .ZN(n896) );
  NAND2_X1 U999 ( .A1(n897), .A2(n896), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(G106), .A2(n898), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(G142), .A2(n899), .ZN(n900) );
  NAND2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U1003 ( .A(n902), .B(KEYINPUT45), .Z(n903) );
  NOR2_X1 U1004 ( .A1(n904), .A2(n903), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1006 ( .A(n908), .B(n907), .Z(n912) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n913), .ZN(G395) );
  NOR2_X1 U1010 ( .A1(G401), .A2(n914), .ZN(n918) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(G397), .A2(n916), .ZN(n917) );
  NAND2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1015 ( .A1(n919), .A2(G395), .ZN(n920) );
  XNOR2_X1 U1016 ( .A(n920), .B(KEYINPUT116), .ZN(G308) );
  INV_X1 U1017 ( .A(G308), .ZN(G225) );
  INV_X1 U1018 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1019 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1030) );
  INV_X1 U1020 ( .A(KEYINPUT55), .ZN(n965) );
  XOR2_X1 U1021 ( .A(G2084), .B(G160), .Z(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(KEYINPUT117), .B(n927), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n934) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n932), .B(KEYINPUT51), .ZN(n933) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(n935), .B(KEYINPUT118), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n943) );
  XOR2_X1 U1033 ( .A(G2072), .B(n938), .Z(n940) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1036 ( .A(KEYINPUT50), .B(n941), .Z(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(KEYINPUT52), .B(n944), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n965), .A2(n945), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n946), .A2(G29), .ZN(n1028) );
  XNOR2_X1 U1041 ( .A(G2090), .B(G35), .ZN(n960) );
  XNOR2_X1 U1042 ( .A(G1996), .B(G32), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(G26), .B(G2067), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n955) );
  XOR2_X1 U1045 ( .A(G2072), .B(G33), .Z(n949) );
  NAND2_X1 U1046 ( .A1(n949), .A2(G28), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(G27), .B(n950), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(KEYINPUT119), .B(n951), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(G25), .B(G1991), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(KEYINPUT53), .B(n958), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1055 ( .A(G2084), .B(G34), .Z(n961) );
  XNOR2_X1 U1056 ( .A(KEYINPUT54), .B(n961), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(n965), .B(n964), .ZN(n967) );
  INV_X1 U1059 ( .A(G29), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(G11), .A2(n968), .ZN(n1026) );
  XNOR2_X1 U1062 ( .A(G16), .B(KEYINPUT56), .ZN(n997) );
  XNOR2_X1 U1063 ( .A(G1966), .B(G168), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(n971), .B(KEYINPUT57), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(KEYINPUT120), .B(n972), .ZN(n995) );
  XOR2_X1 U1067 ( .A(n973), .B(G1341), .Z(n980) );
  XNOR2_X1 U1068 ( .A(G171), .B(G1961), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(n974), .B(KEYINPUT121), .ZN(n977) );
  XOR2_X1 U1070 ( .A(G1348), .B(n975), .Z(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(KEYINPUT122), .B(n978), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n993) );
  XNOR2_X1 U1074 ( .A(n981), .B(G1956), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n986) );
  XOR2_X1 U1076 ( .A(G1971), .B(G303), .Z(n984) );
  XNOR2_X1 U1077 ( .A(KEYINPUT123), .B(n984), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1081 ( .A(KEYINPUT124), .B(n991), .Z(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n1024) );
  INV_X1 U1085 ( .A(G16), .ZN(n1022) );
  XNOR2_X1 U1086 ( .A(G1971), .B(G22), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(G24), .B(G1986), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(G1976), .B(G23), .Z(n1000) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XOR2_X1 U1091 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n1002) );
  XNOR2_X1 U1092 ( .A(n1003), .B(n1002), .ZN(n1016) );
  XOR2_X1 U1093 ( .A(G1348), .B(KEYINPUT59), .Z(n1004) );
  XNOR2_X1 U1094 ( .A(G4), .B(n1004), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(G19), .B(G1341), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G1956), .B(G20), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(G1981), .B(G6), .ZN(n1007) );
  NOR2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(n1011), .B(KEYINPUT60), .ZN(n1012) );
  XOR2_X1 U1102 ( .A(KEYINPUT125), .B(n1012), .Z(n1014) );
  XNOR2_X1 U1103 ( .A(G1966), .B(G21), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1019) );
  XOR2_X1 U1106 ( .A(G5), .B(n1017), .Z(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1020), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(n1030), .B(n1029), .ZN(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
  INV_X1 U1115 ( .A(G171), .ZN(G301) );
endmodule

