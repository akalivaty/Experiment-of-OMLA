//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT75), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G137), .ZN(new_n191));
  INV_X1    g005(.A(G221), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n192), .A2(new_n187), .A3(G953), .ZN(new_n193));
  XOR2_X1   g007(.A(new_n191), .B(new_n193), .Z(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT77), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G125), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(KEYINPUT77), .ZN(new_n200));
  OAI21_X1  g014(.A(G140), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(G125), .A2(G140), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n196), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT77), .B(G125), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n206));
  OAI211_X1 g020(.A(KEYINPUT78), .B(G146), .C1(new_n204), .C2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G140), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n203), .B1(new_n205), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT16), .ZN(new_n210));
  OR2_X1    g024(.A1(KEYINPUT78), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(new_n205), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n196), .A3(new_n208), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT78), .A2(G146), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n211), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G119), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT76), .B1(new_n216), .B2(G128), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT76), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G119), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(G128), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT24), .B(G110), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n219), .A2(KEYINPUT23), .A3(G119), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n216), .A2(G128), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n221), .B(new_n225), .C1(new_n226), .C2(KEYINPUT23), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n224), .B1(G110), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n207), .A2(new_n215), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT79), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT79), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n207), .A2(new_n215), .A3(new_n231), .A4(new_n228), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(G125), .B(G140), .Z(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(G146), .ZN(new_n235));
  OR2_X1    g049(.A1(new_n227), .A2(G110), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n222), .A2(new_n223), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n210), .A2(G146), .A3(new_n213), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT80), .B1(new_n233), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT80), .ZN(new_n243));
  AOI211_X1 g057(.A(new_n243), .B(new_n240), .C1(new_n230), .C2(new_n232), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n195), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n233), .A2(new_n241), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n194), .ZN(new_n247));
  AOI21_X1  g061(.A(G902), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n253), .B1(new_n248), .B2(new_n250), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n190), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n245), .A2(new_n247), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n190), .A2(G902), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(G214), .B1(G237), .B2(G902), .ZN(new_n261));
  XOR2_X1   g075(.A(G116), .B(G119), .Z(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT2), .B(G113), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n262), .A2(KEYINPUT67), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n265));
  XOR2_X1   g079(.A(KEYINPUT2), .B(G113), .Z(new_n266));
  XNOR2_X1  g080(.A(G116), .B(G119), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI22_X1  g082(.A1(new_n264), .A2(new_n268), .B1(new_n267), .B2(new_n266), .ZN(new_n269));
  INV_X1    g083(.A(G104), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT3), .B1(new_n270), .B2(G107), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT3), .ZN(new_n272));
  INV_X1    g086(.A(G107), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(G104), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n270), .A2(G107), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n271), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G101), .ZN(new_n277));
  OR2_X1    g091(.A1(new_n277), .A2(KEYINPUT4), .ZN(new_n278));
  INV_X1    g092(.A(G101), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n271), .A2(new_n274), .A3(new_n279), .A4(new_n275), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(KEYINPUT4), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n269), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n275), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n270), .A2(G107), .ZN(new_n284));
  OAI21_X1  g098(.A(G101), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n280), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT5), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n216), .A3(G116), .ZN(new_n289));
  OAI211_X1 g103(.A(G113), .B(new_n289), .C1(new_n262), .C2(new_n288), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n287), .B(new_n290), .C1(new_n264), .C2(new_n268), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n282), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G110), .B(G122), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n282), .A2(new_n293), .A3(new_n291), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT6), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n297), .A2(KEYINPUT83), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n295), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(G143), .B(G146), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT0), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n300), .B1(new_n301), .B2(new_n219), .ZN(new_n302));
  XOR2_X1   g116(.A(KEYINPUT0), .B(G128), .Z(new_n303));
  OAI21_X1  g117(.A(new_n302), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n212), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n300), .A2(new_n306), .A3(G128), .ZN(new_n307));
  INV_X1    g121(.A(G146), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G143), .ZN(new_n309));
  INV_X1    g123(.A(G143), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G146), .ZN(new_n311));
  AOI21_X1  g125(.A(G128), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n306), .A2(new_n308), .A3(G143), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT65), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n308), .A2(G143), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT1), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT65), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n316), .B(new_n317), .C1(new_n300), .C2(G128), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n307), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n305), .B1(new_n319), .B2(new_n212), .ZN(new_n320));
  INV_X1    g134(.A(G224), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(G953), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT84), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n320), .B(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n292), .B(new_n294), .C1(KEYINPUT83), .C2(new_n297), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n299), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(KEYINPUT7), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n305), .B(new_n327), .C1(new_n319), .C2(new_n212), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n296), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n290), .B1(new_n264), .B2(new_n268), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n286), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n291), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n293), .B(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n327), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n332), .A2(new_n334), .B1(new_n320), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(G902), .B1(new_n329), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(G210), .B1(G237), .B2(G902), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n326), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n326), .B2(new_n337), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n261), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT86), .ZN(new_n342));
  XNOR2_X1  g156(.A(G113), .B(G122), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(new_n270), .ZN(new_n344));
  INV_X1    g158(.A(G237), .ZN(new_n345));
  INV_X1    g159(.A(G953), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(G214), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n310), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n345), .A2(new_n346), .A3(G143), .A4(G214), .ZN(new_n349));
  NAND2_X1  g163(.A1(KEYINPUT18), .A2(G131), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n209), .A2(new_n308), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n349), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(KEYINPUT18), .A3(G131), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT87), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n354), .A2(new_n355), .ZN(new_n357));
  OAI221_X1 g171(.A(new_n351), .B1(new_n235), .B2(new_n352), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G131), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n353), .B(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT17), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI211_X1 g176(.A(new_n361), .B(new_n359), .C1(new_n348), .C2(new_n349), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n207), .B2(new_n215), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT90), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI211_X1 g180(.A(KEYINPUT90), .B(new_n363), .C1(new_n207), .C2(new_n215), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n344), .B(new_n358), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n353), .B(G131), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT88), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n360), .A2(KEYINPUT88), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n234), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n209), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n374), .B1(new_n375), .B2(KEYINPUT19), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n308), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n371), .A2(new_n372), .A3(new_n239), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n358), .ZN(new_n379));
  INV_X1    g193(.A(new_n344), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n368), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT91), .ZN(new_n383));
  NOR2_X1   g197(.A1(G475), .A2(G902), .ZN(new_n384));
  XOR2_X1   g198(.A(new_n384), .B(KEYINPUT92), .Z(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT91), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n368), .A2(new_n387), .A3(new_n381), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n383), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n385), .A2(KEYINPUT20), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n389), .A2(KEYINPUT20), .B1(new_n382), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n358), .B1(new_n366), .B2(new_n367), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n380), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n368), .ZN(new_n394));
  INV_X1    g208(.A(G902), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n396), .A2(G475), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G116), .B(G122), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n273), .ZN(new_n400));
  INV_X1    g214(.A(G116), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT14), .A3(G122), .ZN(new_n402));
  XOR2_X1   g216(.A(G116), .B(G122), .Z(new_n403));
  OAI211_X1 g217(.A(G107), .B(new_n402), .C1(new_n403), .C2(KEYINPUT14), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n310), .A2(G128), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n310), .A2(G128), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G134), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n406), .A2(new_n407), .A3(G134), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n400), .B(new_n404), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n400), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n399), .A2(new_n273), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT93), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n403), .A2(G107), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT93), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n400), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n411), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT13), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n405), .B1(new_n407), .B2(new_n420), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n421), .A2(KEYINPUT94), .B1(KEYINPUT13), .B2(new_n406), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(KEYINPUT94), .B2(new_n421), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G134), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n419), .A2(new_n424), .A3(KEYINPUT95), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT95), .B1(new_n419), .B2(new_n424), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n412), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT9), .B(G234), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(G217), .A3(new_n346), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n430), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n412), .B(new_n432), .C1(new_n425), .C2(new_n426), .ZN(new_n433));
  AOI21_X1  g247(.A(G902), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G478), .ZN(new_n435));
  NOR2_X1   g249(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n435), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n434), .B(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(G902), .B(G953), .C1(new_n187), .C2(new_n345), .ZN(new_n441));
  XOR2_X1   g255(.A(new_n441), .B(KEYINPUT97), .Z(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(G898), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n346), .A2(G952), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n187), .B2(new_n345), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G469), .ZN(new_n449));
  XNOR2_X1  g263(.A(G110), .B(G140), .ZN(new_n450));
  INV_X1    g264(.A(G227), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(G953), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n450), .B(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n300), .A2(new_n306), .A3(G128), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n310), .A2(G146), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n219), .B1(new_n456), .B2(new_n315), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n457), .A3(new_n316), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n287), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT10), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n278), .A2(new_n304), .A3(new_n281), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n287), .A2(KEYINPUT10), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n461), .B(new_n462), .C1(new_n319), .C2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT11), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n409), .B2(G137), .ZN(new_n466));
  INV_X1    g280(.A(G137), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(KEYINPUT11), .A3(G134), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n409), .A2(G137), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G131), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n466), .A2(new_n468), .A3(new_n359), .A4(new_n469), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(KEYINPUT64), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT64), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n474), .A3(G131), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n454), .B1(new_n464), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n317), .B1(new_n457), .B2(new_n316), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n312), .A2(KEYINPUT65), .A3(new_n313), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n455), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT82), .B1(new_n481), .B2(new_n287), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT82), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n319), .A2(new_n483), .A3(new_n286), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n459), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n477), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT12), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n485), .A2(KEYINPUT12), .A3(new_n477), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n478), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n464), .A2(new_n477), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n464), .A2(new_n477), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n454), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n449), .B(new_n395), .C1(new_n490), .C2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(new_n454), .A3(new_n493), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n491), .B1(new_n488), .B2(new_n489), .ZN(new_n497));
  OAI211_X1 g311(.A(G469), .B(new_n496), .C1(new_n497), .C2(new_n454), .ZN(new_n498));
  NAND2_X1  g312(.A1(G469), .A2(G902), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n495), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n192), .B1(new_n429), .B2(new_n395), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n342), .A2(new_n398), .A3(new_n448), .A4(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n269), .ZN(new_n506));
  INV_X1    g320(.A(new_n469), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n409), .A2(G137), .ZN(new_n508));
  OAI21_X1  g322(.A(G131), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n472), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n481), .A2(KEYINPUT66), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT66), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n319), .B2(new_n510), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n473), .A2(new_n475), .A3(new_n304), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT30), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n506), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT68), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n481), .A2(new_n519), .A3(new_n511), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT68), .B1(new_n319), .B2(new_n510), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT30), .A4(new_n515), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT69), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n522), .A2(new_n523), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n518), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT31), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n520), .A2(new_n521), .A3(new_n506), .A4(new_n515), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT26), .B(G101), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n345), .A2(new_n346), .A3(G210), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n532), .B(new_n533), .Z(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n526), .A2(new_n527), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT72), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n526), .A2(KEYINPUT72), .A3(new_n527), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n516), .A2(new_n517), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n269), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n522), .A2(new_n523), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n522), .A2(new_n523), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n536), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT71), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT71), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n526), .A2(new_n549), .A3(new_n536), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(KEYINPUT31), .A3(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n516), .A2(new_n269), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT28), .B1(new_n552), .B2(new_n529), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT73), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n515), .B(new_n506), .C1(new_n319), .C2(new_n510), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT28), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n554), .B1(new_n553), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n535), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n541), .A2(new_n551), .A3(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(G472), .A2(G902), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n561), .A2(KEYINPUT74), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT74), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT32), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n520), .A2(new_n521), .A3(new_n515), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n269), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n557), .B1(new_n567), .B2(new_n528), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n557), .B2(new_n556), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT29), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n535), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(G902), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n555), .A2(new_n559), .A3(new_n535), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n546), .A2(new_n529), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n570), .B1(new_n574), .B2(new_n534), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n572), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G472), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n561), .A2(KEYINPUT32), .A3(new_n562), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n260), .B(new_n505), .C1(new_n565), .C2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(G101), .ZN(G3));
  AND3_X1   g395(.A1(new_n255), .A2(new_n258), .A3(new_n503), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n561), .A2(new_n562), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT74), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n561), .A2(KEYINPUT74), .A3(new_n562), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n561), .A2(new_n395), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G472), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n582), .A2(new_n585), .A3(new_n586), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n431), .A2(new_n433), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT33), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n431), .A2(new_n592), .A3(new_n433), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(G478), .A3(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n435), .A2(new_n395), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n434), .B2(new_n435), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n389), .A2(KEYINPUT20), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n382), .A2(new_n390), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n397), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n341), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n447), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n589), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT34), .B(G104), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G6));
  INV_X1    g421(.A(new_n589), .ZN(new_n608));
  INV_X1    g422(.A(new_n440), .ZN(new_n609));
  XOR2_X1   g423(.A(new_n447), .B(KEYINPUT99), .Z(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n603), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT20), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n383), .A2(new_n612), .A3(new_n386), .A4(new_n388), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n598), .A2(KEYINPUT98), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n598), .A2(new_n613), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI211_X1 g431(.A(new_n397), .B(new_n611), .C1(new_n614), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n608), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT35), .B(G107), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G9));
  NAND3_X1  g435(.A1(new_n585), .A2(new_n588), .A3(new_n586), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n504), .ZN(new_n623));
  INV_X1    g437(.A(new_n253), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n256), .A2(new_n395), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(new_n249), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n189), .B1(new_n626), .B2(new_n251), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n242), .A2(new_n244), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n195), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n257), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(KEYINPUT100), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n255), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n623), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT37), .B(G110), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  INV_X1    g453(.A(KEYINPUT32), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n585), .A2(new_n640), .A3(new_n586), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n577), .A2(new_n578), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n500), .A2(new_n502), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n341), .ZN(new_n645));
  INV_X1    g459(.A(new_n446), .ZN(new_n646));
  INV_X1    g460(.A(G900), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n646), .B1(new_n442), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n440), .A2(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n598), .A2(KEYINPUT98), .A3(new_n613), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT98), .B1(new_n598), .B2(new_n613), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n601), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n633), .B2(new_n635), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n643), .A2(new_n645), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT101), .B(G128), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G30));
  XOR2_X1   g470(.A(new_n648), .B(KEYINPUT39), .Z(new_n657));
  NAND2_X1  g471(.A1(new_n503), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n659));
  INV_X1    g473(.A(new_n261), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n339), .A2(new_n340), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT38), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n550), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n549), .B1(new_n526), .B2(new_n536), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n534), .B1(new_n567), .B2(new_n528), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(KEYINPUT102), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n666), .A2(KEYINPUT102), .ZN(new_n668));
  NOR4_X1   g482(.A1(new_n664), .A2(new_n665), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n669), .B2(G902), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n578), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n641), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n636), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n600), .A2(new_n601), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n609), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(KEYINPUT40), .B2(new_n658), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n663), .A2(new_n672), .A3(new_n673), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G143), .ZN(G45));
  AND2_X1   g492(.A1(new_n594), .A2(new_n596), .ZN(new_n679));
  INV_X1    g493(.A(new_n648), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n679), .B(new_n680), .C1(new_n391), .C2(new_n397), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n633), .B2(new_n635), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n643), .A2(new_n645), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  AOI21_X1  g498(.A(new_n259), .B1(new_n641), .B2(new_n642), .ZN(new_n685));
  INV_X1    g499(.A(new_n604), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n490), .A2(new_n494), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n395), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(G469), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n502), .A3(new_n495), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT103), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n685), .A2(new_n686), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND3_X1  g508(.A1(new_n685), .A2(new_n618), .A3(new_n691), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  AND2_X1   g510(.A1(new_n398), .A2(new_n448), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n690), .A2(new_n341), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n643), .A2(new_n697), .A3(new_n636), .A4(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT104), .B(G119), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G21));
  NAND2_X1  g515(.A1(new_n569), .A2(KEYINPUT105), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n535), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n569), .A2(KEYINPUT105), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n541), .B(new_n551), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n562), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n588), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n259), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n674), .A2(new_n609), .A3(new_n603), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n708), .A2(new_n610), .A3(new_n691), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  INV_X1    g526(.A(new_n707), .ZN(new_n713));
  INV_X1    g527(.A(new_n681), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n636), .A3(new_n714), .A4(new_n698), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  INV_X1    g530(.A(KEYINPUT42), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n644), .A2(KEYINPUT106), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n661), .A2(new_n261), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n644), .B2(KEYINPUT106), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n714), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n643), .A2(new_n260), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT107), .B1(new_n583), .B2(new_n640), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n579), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n583), .A2(KEYINPUT107), .A3(new_n640), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n259), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n714), .A2(new_n718), .A3(KEYINPUT42), .A4(new_n720), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n717), .A2(new_n723), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n359), .ZN(G33));
  NAND2_X1  g546(.A1(new_n718), .A2(new_n720), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n652), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n685), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G134), .ZN(G36));
  NAND3_X1  g550(.A1(new_n600), .A2(new_n601), .A3(new_n679), .ZN(new_n737));
  XOR2_X1   g551(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n398), .A2(KEYINPUT43), .A3(new_n679), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n737), .A2(KEYINPUT109), .A3(new_n738), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n622), .A3(new_n636), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n496), .B1(new_n497), .B2(new_n454), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(G469), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n748), .A2(new_n749), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n499), .ZN(new_n754));
  INV_X1    g568(.A(new_n495), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n499), .B1(new_n751), .B2(new_n752), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n501), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(new_n261), .A3(new_n661), .A4(new_n657), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n744), .A2(KEYINPUT44), .A3(new_n622), .A4(new_n636), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n762), .A2(new_n763), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n747), .B(new_n761), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G137), .ZN(G39));
  XNOR2_X1  g582(.A(new_n759), .B(KEYINPUT47), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n260), .A2(new_n681), .A3(new_n719), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n641), .A3(new_n642), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  AOI211_X1 g586(.A(new_n259), .B(new_n504), .C1(new_n641), .C2(new_n642), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n602), .A2(new_n342), .A3(new_n610), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n589), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT111), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n563), .A2(new_n564), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n774), .A3(new_n588), .A4(new_n582), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n580), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n342), .A2(new_n610), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n674), .A2(new_n440), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  AOI22_X1  g599(.A1(new_n608), .A2(new_n785), .B1(new_n623), .B2(new_n636), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n777), .A2(new_n781), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n617), .A2(new_n614), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n500), .A2(new_n502), .A3(new_n680), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n440), .A2(new_n261), .A3(new_n661), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n788), .A2(new_n791), .A3(new_n601), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n641), .B2(new_n642), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n721), .A2(new_n707), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n636), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT42), .B1(new_n685), .B2(new_n722), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT32), .B1(new_n561), .B2(new_n562), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n578), .B(new_n577), .C1(new_n797), .C2(KEYINPUT107), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n260), .B1(new_n798), .B2(new_n726), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n729), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n735), .B(new_n795), .C1(new_n796), .C2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n692), .A2(new_n695), .A3(new_n699), .A4(new_n711), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n787), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n654), .A2(new_n715), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n654), .A2(KEYINPUT112), .A3(new_n715), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n709), .A2(new_n627), .A3(new_n632), .A4(new_n789), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n808), .B1(new_n672), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n806), .A2(new_n683), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n672), .A2(new_n809), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n654), .A2(new_n683), .A3(new_n812), .A4(new_n715), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n808), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n803), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n645), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n641), .B2(new_n642), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n820), .A2(new_n682), .B1(new_n672), .B2(new_n809), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(KEYINPUT52), .A3(new_n654), .A4(new_n715), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n814), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n803), .A2(KEYINPUT53), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n818), .A2(new_n824), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n787), .A2(new_n801), .A3(new_n802), .A4(new_n817), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n801), .A2(new_n802), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n580), .A2(new_n778), .A3(new_n780), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n778), .B1(new_n580), .B2(new_n780), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n505), .A2(new_n779), .A3(new_n588), .ZN(new_n830));
  OAI22_X1  g644(.A1(new_n830), .A2(new_n673), .B1(new_n589), .B2(new_n784), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n828), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n827), .A2(new_n823), .A3(new_n832), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n815), .A2(new_n826), .B1(new_n833), .B2(new_n817), .ZN(new_n834));
  XOR2_X1   g648(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n835));
  AOI22_X1  g649(.A1(new_n825), .A2(KEYINPUT54), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n672), .A2(new_n259), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n690), .A2(new_n446), .A3(new_n719), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n674), .A3(new_n679), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT114), .Z(new_n841));
  NAND3_X1  g655(.A1(new_n708), .A2(new_n744), .A3(new_n646), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n662), .A2(new_n660), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n842), .A2(new_n690), .A3(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT50), .ZN(new_n845));
  INV_X1    g659(.A(new_n769), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n689), .A2(new_n495), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n846), .B1(new_n502), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n842), .A2(new_n719), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n673), .A2(new_n707), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n744), .A2(new_n838), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n849), .A2(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n841), .A2(new_n845), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n852), .A2(new_n728), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT48), .Z(new_n858));
  INV_X1    g672(.A(new_n698), .ZN(new_n859));
  INV_X1    g673(.A(new_n602), .ZN(new_n860));
  OAI221_X1 g674(.A(new_n445), .B1(new_n859), .B2(new_n842), .C1(new_n839), .C2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT115), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n854), .A2(new_n855), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n836), .A2(new_n856), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n865), .B1(G952), .B2(G953), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n848), .A2(KEYINPUT49), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n848), .A2(KEYINPUT49), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n662), .A2(new_n261), .A3(new_n502), .ZN(new_n869));
  NOR4_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n737), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n837), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n866), .A2(new_n871), .ZN(G75));
  NOR2_X1   g686(.A1(new_n834), .A2(new_n395), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(G210), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n299), .A2(new_n325), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(new_n324), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT55), .ZN(new_n877));
  NOR2_X1   g691(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n874), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n877), .B1(new_n874), .B2(new_n878), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n346), .A2(G952), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(G51));
  AOI21_X1  g696(.A(KEYINPUT118), .B1(new_n834), .B2(new_n835), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n833), .A2(new_n817), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n803), .A2(new_n815), .A3(KEYINPUT53), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n835), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n886), .A2(KEYINPUT118), .A3(new_n887), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n499), .B(KEYINPUT117), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT57), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n687), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n753), .B(KEYINPUT119), .Z(new_n895));
  NAND2_X1  g709(.A1(new_n873), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n881), .B1(new_n894), .B2(new_n896), .ZN(G54));
  NAND3_X1  g711(.A1(new_n873), .A2(KEYINPUT58), .A3(G475), .ZN(new_n898));
  INV_X1    g712(.A(new_n388), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n387), .B1(new_n368), .B2(new_n381), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n898), .A2(new_n902), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n903), .A2(new_n904), .A3(new_n881), .ZN(G60));
  XNOR2_X1  g719(.A(new_n595), .B(KEYINPUT59), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n591), .B(new_n593), .C1(new_n836), .C2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n906), .B1(new_n591), .B2(new_n593), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n889), .A2(new_n890), .A3(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n881), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n907), .A2(new_n909), .A3(new_n910), .ZN(G63));
  NAND2_X1  g725(.A1(G217), .A2(G902), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT60), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n813), .A2(new_n808), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n654), .A2(KEYINPUT112), .A3(new_n715), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT112), .B1(new_n654), .B2(new_n715), .ZN(new_n917));
  INV_X1    g731(.A(new_n683), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n915), .B1(new_n919), .B2(new_n810), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n795), .A2(new_n735), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n731), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n802), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n832), .A2(new_n922), .A3(KEYINPUT53), .A4(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT53), .B1(new_n803), .B2(new_n823), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n630), .B(new_n914), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n886), .A2(KEYINPUT121), .A3(new_n630), .A4(new_n914), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n256), .B(KEYINPUT122), .Z(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n834), .B2(new_n913), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n929), .A2(new_n910), .A3(new_n930), .A4(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n933), .A2(KEYINPUT120), .A3(KEYINPUT61), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT61), .B1(new_n933), .B2(KEYINPUT120), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(G66));
  OAI21_X1  g750(.A(G953), .B1(new_n443), .B2(new_n321), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n832), .A2(new_n923), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n939), .B2(G953), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n875), .B1(G898), .B2(new_n346), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT123), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n940), .B(new_n942), .ZN(G69));
  OAI21_X1  g757(.A(new_n542), .B1(new_n524), .B2(new_n525), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(new_n376), .Z(new_n945));
  NAND2_X1  g759(.A1(new_n919), .A2(new_n677), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT62), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n658), .A2(new_n719), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n685), .B(new_n948), .C1(new_n602), .C2(new_n783), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n767), .A2(new_n771), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n919), .A2(new_n951), .A3(new_n677), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n947), .A2(new_n950), .A3(new_n346), .A4(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n945), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n451), .A2(G900), .A3(G953), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n759), .A2(new_n657), .A3(new_n710), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n958));
  OR3_X1    g772(.A1(new_n957), .A2(new_n799), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n957), .B2(new_n799), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n731), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n961), .A2(new_n962), .A3(new_n735), .A4(new_n771), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n747), .A2(new_n761), .ZN(new_n964));
  INV_X1    g778(.A(new_n766), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(new_n764), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n918), .B1(new_n804), .B2(new_n805), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n807), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT124), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n767), .A2(new_n919), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n963), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n956), .B1(new_n972), .B2(G953), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n955), .B1(new_n973), .B2(new_n945), .ZN(G72));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n975));
  AOI211_X1 g789(.A(new_n938), .B(new_n963), .C1(new_n969), .C2(new_n971), .ZN(new_n976));
  NAND2_X1  g790(.A1(G472), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT63), .Z(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n975), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n972), .A2(new_n939), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n981), .A2(KEYINPUT126), .A3(new_n978), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n546), .A2(new_n534), .A3(new_n529), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n534), .B1(new_n546), .B2(new_n529), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n947), .A2(new_n950), .A3(new_n939), .A4(new_n952), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(new_n978), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n548), .B(new_n550), .C1(new_n574), .C2(new_n534), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n978), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n818), .B2(new_n824), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n987), .A2(new_n990), .A3(new_n881), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n984), .A2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n984), .A2(new_n991), .A3(KEYINPUT127), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(G57));
endmodule


