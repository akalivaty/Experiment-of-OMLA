

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U550 ( .A1(G2105), .A2(G2104), .ZN(n558) );
  INV_X1 U551 ( .A(n734), .ZN(n751) );
  XNOR2_X1 U552 ( .A(n524), .B(n523), .ZN(n774) );
  OR2_X1 U553 ( .A1(n760), .A2(n750), .ZN(n758) );
  AND2_X1 U554 ( .A1(n529), .A2(n528), .ZN(G160) );
  NAND2_X1 U555 ( .A1(n774), .A2(n522), .ZN(n521) );
  AND2_X1 U556 ( .A1(n775), .A2(n968), .ZN(n522) );
  XNOR2_X1 U557 ( .A(n713), .B(n712), .ZN(n715) );
  AND2_X1 U558 ( .A1(n521), .A2(n766), .ZN(n767) );
  INV_X1 U559 ( .A(G2104), .ZN(n564) );
  INV_X1 U560 ( .A(KEYINPUT89), .ZN(n711) );
  NOR2_X1 U561 ( .A1(n717), .A2(G299), .ZN(n535) );
  XNOR2_X1 U562 ( .A(KEYINPUT92), .B(KEYINPUT30), .ZN(n740) );
  INV_X1 U563 ( .A(KEYINPUT32), .ZN(n523) );
  NAND2_X1 U564 ( .A1(n526), .A2(n517), .ZN(n525) );
  INV_X1 U565 ( .A(KEYINPUT17), .ZN(n557) );
  NOR2_X1 U566 ( .A1(n603), .A2(n602), .ZN(n905) );
  NOR2_X1 U567 ( .A1(G651), .A2(n676), .ZN(n671) );
  AND2_X1 U568 ( .A1(n568), .A2(n565), .ZN(n529) );
  XNOR2_X1 U569 ( .A(n563), .B(n562), .ZN(n528) );
  AND2_X1 U570 ( .A1(n525), .A2(n520), .ZN(n516) );
  AND2_X1 U571 ( .A1(n785), .A2(n519), .ZN(n517) );
  XOR2_X1 U572 ( .A(n746), .B(KEYINPUT93), .Z(n518) );
  XNOR2_X1 U573 ( .A(n734), .B(n711), .ZN(n723) );
  NOR2_X1 U574 ( .A1(G164), .A2(G1384), .ZN(n786) );
  XOR2_X1 U575 ( .A(n784), .B(KEYINPUT88), .Z(n519) );
  AND2_X1 U576 ( .A1(n818), .A2(n822), .ZN(n520) );
  NAND2_X1 U577 ( .A1(n762), .A2(n763), .ZN(n775) );
  NAND2_X1 U578 ( .A1(n758), .A2(n757), .ZN(n524) );
  NAND2_X1 U579 ( .A1(n527), .A2(n773), .ZN(n526) );
  XNOR2_X1 U580 ( .A(n769), .B(KEYINPUT95), .ZN(n527) );
  NAND2_X1 U581 ( .A1(n731), .A2(n530), .ZN(n732) );
  NAND2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n530) );
  XNOR2_X1 U583 ( .A(n535), .B(KEYINPUT91), .ZN(n531) );
  NAND2_X1 U584 ( .A1(n533), .A2(n534), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n727), .A2(n726), .ZN(n533) );
  NAND2_X1 U586 ( .A1(n730), .A2(n729), .ZN(n534) );
  XNOR2_X2 U587 ( .A(n558), .B(n557), .ZN(n896) );
  XNOR2_X1 U588 ( .A(n599), .B(KEYINPUT13), .ZN(n536) );
  INV_X1 U589 ( .A(KEYINPUT27), .ZN(n712) );
  XNOR2_X1 U590 ( .A(n741), .B(n740), .ZN(n742) );
  INV_X1 U591 ( .A(G2105), .ZN(n566) );
  AND2_X2 U592 ( .A1(n566), .A2(G2104), .ZN(n893) );
  NOR2_X1 U593 ( .A1(G651), .A2(G543), .ZN(n662) );
  NAND2_X1 U594 ( .A1(G91), .A2(n662), .ZN(n539) );
  INV_X1 U595 ( .A(G651), .ZN(n540) );
  NOR2_X1 U596 ( .A1(G543), .A2(n540), .ZN(n537) );
  XOR2_X1 U597 ( .A(KEYINPUT1), .B(n537), .Z(n675) );
  NAND2_X1 U598 ( .A1(G65), .A2(n675), .ZN(n538) );
  NAND2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n545) );
  XOR2_X1 U600 ( .A(G543), .B(KEYINPUT0), .Z(n676) );
  NAND2_X1 U601 ( .A1(G53), .A2(n671), .ZN(n543) );
  OR2_X1 U602 ( .A1(n540), .A2(n676), .ZN(n541) );
  XOR2_X2 U603 ( .A(KEYINPUT68), .B(n541), .Z(n660) );
  NAND2_X1 U604 ( .A1(G78), .A2(n660), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n544) );
  OR2_X1 U606 ( .A1(n545), .A2(n544), .ZN(G299) );
  NAND2_X1 U607 ( .A1(n662), .A2(G89), .ZN(n546) );
  XNOR2_X1 U608 ( .A(n546), .B(KEYINPUT4), .ZN(n548) );
  NAND2_X1 U609 ( .A1(G76), .A2(n660), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U611 ( .A(n549), .B(KEYINPUT5), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n671), .A2(G51), .ZN(n550) );
  XNOR2_X1 U613 ( .A(n550), .B(KEYINPUT72), .ZN(n552) );
  NAND2_X1 U614 ( .A1(G63), .A2(n675), .ZN(n551) );
  NAND2_X1 U615 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U616 ( .A(KEYINPUT6), .B(n553), .Z(n554) );
  NAND2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U618 ( .A(n556), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U619 ( .A1(G137), .A2(n896), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G2105), .A2(G2104), .ZN(n559) );
  XNOR2_X2 U621 ( .A(n559), .B(KEYINPUT65), .ZN(n627) );
  NAND2_X1 U622 ( .A1(G113), .A2(n627), .ZN(n560) );
  NAND2_X1 U623 ( .A1(n561), .A2(n560), .ZN(n563) );
  INV_X1 U624 ( .A(KEYINPUT66), .ZN(n562) );
  AND2_X1 U625 ( .A1(n564), .A2(G2105), .ZN(n889) );
  NAND2_X1 U626 ( .A1(n889), .A2(G125), .ZN(n565) );
  NAND2_X1 U627 ( .A1(G101), .A2(n893), .ZN(n567) );
  XOR2_X1 U628 ( .A(KEYINPUT23), .B(n567), .Z(n568) );
  XOR2_X1 U629 ( .A(G2438), .B(G2454), .Z(n570) );
  XNOR2_X1 U630 ( .A(G2435), .B(G2430), .ZN(n569) );
  XNOR2_X1 U631 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U632 ( .A(n571), .B(G2427), .Z(n573) );
  XNOR2_X1 U633 ( .A(G1341), .B(G1348), .ZN(n572) );
  XNOR2_X1 U634 ( .A(n573), .B(n572), .ZN(n577) );
  XOR2_X1 U635 ( .A(G2443), .B(G2446), .Z(n575) );
  XNOR2_X1 U636 ( .A(KEYINPUT102), .B(G2451), .ZN(n574) );
  XNOR2_X1 U637 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U638 ( .A(n577), .B(n576), .Z(n578) );
  AND2_X1 U639 ( .A1(G14), .A2(n578), .ZN(G401) );
  AND2_X1 U640 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U641 ( .A(G132), .ZN(G219) );
  INV_X1 U642 ( .A(G82), .ZN(G220) );
  INV_X1 U643 ( .A(G57), .ZN(G237) );
  INV_X1 U644 ( .A(G120), .ZN(G236) );
  NAND2_X1 U645 ( .A1(n893), .A2(G102), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n579), .B(KEYINPUT86), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G138), .A2(n896), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G114), .A2(n627), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G126), .A2(n889), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U652 ( .A1(n585), .A2(n584), .ZN(G164) );
  NAND2_X1 U653 ( .A1(G52), .A2(n671), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G64), .A2(n675), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n592) );
  NAND2_X1 U656 ( .A1(G90), .A2(n662), .ZN(n589) );
  NAND2_X1 U657 ( .A1(G77), .A2(n660), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U659 ( .A(KEYINPUT9), .B(n590), .Z(n591) );
  NOR2_X1 U660 ( .A1(n592), .A2(n591), .ZN(G171) );
  XOR2_X1 U661 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U662 ( .A1(G7), .A2(G661), .ZN(n593) );
  XOR2_X1 U663 ( .A(n593), .B(KEYINPUT10), .Z(n915) );
  NAND2_X1 U664 ( .A1(n915), .A2(G567), .ZN(n594) );
  XOR2_X1 U665 ( .A(KEYINPUT11), .B(n594), .Z(G234) );
  NAND2_X1 U666 ( .A1(G81), .A2(n662), .ZN(n595) );
  XNOR2_X1 U667 ( .A(n595), .B(KEYINPUT70), .ZN(n596) );
  XNOR2_X1 U668 ( .A(n596), .B(KEYINPUT12), .ZN(n598) );
  NAND2_X1 U669 ( .A1(G68), .A2(n660), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U671 ( .A1(G43), .A2(n671), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n536), .A2(n600), .ZN(n603) );
  NAND2_X1 U673 ( .A1(n675), .A2(G56), .ZN(n601) );
  XOR2_X1 U674 ( .A(KEYINPUT14), .B(n601), .Z(n602) );
  NAND2_X1 U675 ( .A1(n905), .A2(G860), .ZN(G153) );
  INV_X1 U676 ( .A(G171), .ZN(G301) );
  NAND2_X1 U677 ( .A1(G868), .A2(G301), .ZN(n613) );
  NAND2_X1 U678 ( .A1(n671), .A2(G54), .ZN(n610) );
  NAND2_X1 U679 ( .A1(G92), .A2(n662), .ZN(n605) );
  NAND2_X1 U680 ( .A1(G66), .A2(n675), .ZN(n604) );
  NAND2_X1 U681 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U682 ( .A1(G79), .A2(n660), .ZN(n606) );
  XNOR2_X1 U683 ( .A(KEYINPUT71), .B(n606), .ZN(n607) );
  NOR2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n609) );
  AND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U686 ( .A(KEYINPUT15), .B(n611), .ZN(n729) );
  INV_X1 U687 ( .A(G868), .ZN(n687) );
  NAND2_X1 U688 ( .A1(n729), .A2(n687), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(G284) );
  XOR2_X1 U690 ( .A(KEYINPUT73), .B(n687), .Z(n614) );
  NOR2_X1 U691 ( .A1(G286), .A2(n614), .ZN(n616) );
  NOR2_X1 U692 ( .A1(G868), .A2(G299), .ZN(n615) );
  NOR2_X1 U693 ( .A1(n616), .A2(n615), .ZN(G297) );
  INV_X1 U694 ( .A(G860), .ZN(n617) );
  NAND2_X1 U695 ( .A1(G559), .A2(n617), .ZN(n618) );
  XNOR2_X1 U696 ( .A(KEYINPUT74), .B(n618), .ZN(n619) );
  INV_X1 U697 ( .A(n729), .ZN(n976) );
  NAND2_X1 U698 ( .A1(n619), .A2(n976), .ZN(n620) );
  XNOR2_X1 U699 ( .A(KEYINPUT16), .B(n620), .ZN(G148) );
  INV_X1 U700 ( .A(n905), .ZN(n983) );
  NOR2_X1 U701 ( .A1(G868), .A2(n983), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G868), .A2(n976), .ZN(n621) );
  NOR2_X1 U703 ( .A1(G559), .A2(n621), .ZN(n622) );
  NOR2_X1 U704 ( .A1(n623), .A2(n622), .ZN(G282) );
  NAND2_X1 U705 ( .A1(G99), .A2(n893), .ZN(n625) );
  NAND2_X1 U706 ( .A1(G135), .A2(n896), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n625), .A2(n624), .ZN(n632) );
  NAND2_X1 U708 ( .A1(G123), .A2(n889), .ZN(n626) );
  XNOR2_X1 U709 ( .A(n626), .B(KEYINPUT18), .ZN(n630) );
  NAND2_X1 U710 ( .A1(G111), .A2(n627), .ZN(n628) );
  XOR2_X1 U711 ( .A(KEYINPUT75), .B(n628), .Z(n629) );
  NAND2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n928) );
  XNOR2_X1 U714 ( .A(n928), .B(G2096), .ZN(n633) );
  INV_X1 U715 ( .A(G2100), .ZN(n850) );
  NAND2_X1 U716 ( .A1(n633), .A2(n850), .ZN(G156) );
  NAND2_X1 U717 ( .A1(G67), .A2(n675), .ZN(n635) );
  NAND2_X1 U718 ( .A1(G80), .A2(n660), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U720 ( .A1(G93), .A2(n662), .ZN(n636) );
  XNOR2_X1 U721 ( .A(KEYINPUT77), .B(n636), .ZN(n637) );
  NOR2_X1 U722 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n671), .A2(G55), .ZN(n639) );
  NAND2_X1 U724 ( .A1(n640), .A2(n639), .ZN(n688) );
  XNOR2_X1 U725 ( .A(n983), .B(KEYINPUT76), .ZN(n642) );
  NAND2_X1 U726 ( .A1(G559), .A2(n976), .ZN(n641) );
  XNOR2_X1 U727 ( .A(n642), .B(n641), .ZN(n685) );
  NOR2_X1 U728 ( .A1(n685), .A2(G860), .ZN(n643) );
  XOR2_X1 U729 ( .A(n688), .B(n643), .Z(G145) );
  NAND2_X1 U730 ( .A1(G50), .A2(n671), .ZN(n645) );
  NAND2_X1 U731 ( .A1(G75), .A2(n660), .ZN(n644) );
  NAND2_X1 U732 ( .A1(n645), .A2(n644), .ZN(n651) );
  NAND2_X1 U733 ( .A1(G62), .A2(n675), .ZN(n646) );
  XNOR2_X1 U734 ( .A(n646), .B(KEYINPUT80), .ZN(n649) );
  NAND2_X1 U735 ( .A1(G88), .A2(n662), .ZN(n647) );
  XOR2_X1 U736 ( .A(KEYINPUT81), .B(n647), .Z(n648) );
  NAND2_X1 U737 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U738 ( .A1(n651), .A2(n650), .ZN(G166) );
  INV_X1 U739 ( .A(G166), .ZN(G303) );
  NAND2_X1 U740 ( .A1(n675), .A2(G60), .ZN(n654) );
  NAND2_X1 U741 ( .A1(G47), .A2(n671), .ZN(n652) );
  XOR2_X1 U742 ( .A(KEYINPUT69), .B(n652), .Z(n653) );
  NAND2_X1 U743 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U744 ( .A1(G85), .A2(n662), .ZN(n655) );
  XNOR2_X1 U745 ( .A(KEYINPUT67), .B(n655), .ZN(n656) );
  NOR2_X1 U746 ( .A1(n657), .A2(n656), .ZN(n659) );
  NAND2_X1 U747 ( .A1(G72), .A2(n660), .ZN(n658) );
  NAND2_X1 U748 ( .A1(n659), .A2(n658), .ZN(G290) );
  NAND2_X1 U749 ( .A1(n660), .A2(G73), .ZN(n661) );
  XOR2_X1 U750 ( .A(KEYINPUT2), .B(n661), .Z(n668) );
  NAND2_X1 U751 ( .A1(n662), .A2(G86), .ZN(n663) );
  XNOR2_X1 U752 ( .A(n663), .B(KEYINPUT78), .ZN(n665) );
  NAND2_X1 U753 ( .A1(G61), .A2(n675), .ZN(n664) );
  NAND2_X1 U754 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U755 ( .A(KEYINPUT79), .B(n666), .Z(n667) );
  NOR2_X1 U756 ( .A1(n668), .A2(n667), .ZN(n670) );
  NAND2_X1 U757 ( .A1(n671), .A2(G48), .ZN(n669) );
  NAND2_X1 U758 ( .A1(n670), .A2(n669), .ZN(G305) );
  NAND2_X1 U759 ( .A1(G49), .A2(n671), .ZN(n673) );
  NAND2_X1 U760 ( .A1(G74), .A2(G651), .ZN(n672) );
  NAND2_X1 U761 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U762 ( .A1(n675), .A2(n674), .ZN(n678) );
  NAND2_X1 U763 ( .A1(n676), .A2(G87), .ZN(n677) );
  NAND2_X1 U764 ( .A1(n678), .A2(n677), .ZN(G288) );
  XOR2_X1 U765 ( .A(G303), .B(G290), .Z(n679) );
  XNOR2_X1 U766 ( .A(n679), .B(G305), .ZN(n680) );
  XNOR2_X1 U767 ( .A(KEYINPUT19), .B(n680), .ZN(n682) );
  XNOR2_X1 U768 ( .A(G288), .B(KEYINPUT82), .ZN(n681) );
  XNOR2_X1 U769 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U770 ( .A(n683), .B(G299), .ZN(n684) );
  XNOR2_X1 U771 ( .A(n684), .B(n688), .ZN(n904) );
  XNOR2_X1 U772 ( .A(n685), .B(n904), .ZN(n686) );
  NAND2_X1 U773 ( .A1(n686), .A2(G868), .ZN(n690) );
  NAND2_X1 U774 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U775 ( .A1(n690), .A2(n689), .ZN(G295) );
  NAND2_X1 U776 ( .A1(G2078), .A2(G2084), .ZN(n691) );
  XOR2_X1 U777 ( .A(KEYINPUT20), .B(n691), .Z(n692) );
  NAND2_X1 U778 ( .A1(G2090), .A2(n692), .ZN(n693) );
  XNOR2_X1 U779 ( .A(KEYINPUT21), .B(n693), .ZN(n694) );
  NAND2_X1 U780 ( .A1(n694), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U781 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U782 ( .A1(G236), .A2(G237), .ZN(n695) );
  NAND2_X1 U783 ( .A1(G69), .A2(n695), .ZN(n696) );
  XNOR2_X1 U784 ( .A(KEYINPUT83), .B(n696), .ZN(n697) );
  NAND2_X1 U785 ( .A1(n697), .A2(G108), .ZN(n837) );
  NAND2_X1 U786 ( .A1(G567), .A2(n837), .ZN(n698) );
  XNOR2_X1 U787 ( .A(n698), .B(KEYINPUT84), .ZN(n703) );
  NOR2_X1 U788 ( .A1(G220), .A2(G219), .ZN(n699) );
  XOR2_X1 U789 ( .A(KEYINPUT22), .B(n699), .Z(n700) );
  NOR2_X1 U790 ( .A1(G218), .A2(n700), .ZN(n701) );
  NAND2_X1 U791 ( .A1(G96), .A2(n701), .ZN(n838) );
  NAND2_X1 U792 ( .A1(G2106), .A2(n838), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U794 ( .A(KEYINPUT85), .B(n704), .Z(n839) );
  NAND2_X1 U795 ( .A1(G661), .A2(G483), .ZN(n705) );
  NOR2_X1 U796 ( .A1(n839), .A2(n705), .ZN(n836) );
  NAND2_X1 U797 ( .A1(n836), .A2(G36), .ZN(G176) );
  AND2_X1 U798 ( .A1(n786), .A2(G40), .ZN(n707) );
  NAND2_X1 U799 ( .A1(G160), .A2(n707), .ZN(n709) );
  INV_X1 U800 ( .A(KEYINPUT64), .ZN(n708) );
  XNOR2_X2 U801 ( .A(n709), .B(n708), .ZN(n734) );
  INV_X1 U802 ( .A(n734), .ZN(n710) );
  NAND2_X2 U803 ( .A1(n710), .A2(G8), .ZN(n783) );
  NAND2_X1 U804 ( .A1(G2072), .A2(n723), .ZN(n713) );
  INV_X1 U805 ( .A(n723), .ZN(n733) );
  NAND2_X1 U806 ( .A1(n733), .A2(G1956), .ZN(n714) );
  NAND2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n717) );
  NAND2_X1 U808 ( .A1(G299), .A2(n717), .ZN(n716) );
  XNOR2_X1 U809 ( .A(n716), .B(KEYINPUT28), .ZN(n731) );
  NOR2_X1 U810 ( .A1(n729), .A2(n983), .ZN(n722) );
  NAND2_X1 U811 ( .A1(G1996), .A2(n734), .ZN(n718) );
  XNOR2_X1 U812 ( .A(n718), .B(KEYINPUT26), .ZN(n720) );
  NAND2_X1 U813 ( .A1(G1341), .A2(n751), .ZN(n719) );
  NAND2_X1 U814 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U815 ( .A(KEYINPUT90), .B(n721), .Z(n728) );
  NAND2_X1 U816 ( .A1(n722), .A2(n728), .ZN(n727) );
  NAND2_X1 U817 ( .A1(G1348), .A2(n751), .ZN(n725) );
  NAND2_X1 U818 ( .A1(G2067), .A2(n723), .ZN(n724) );
  NAND2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n728), .A2(n905), .ZN(n730) );
  XNOR2_X1 U821 ( .A(n732), .B(KEYINPUT29), .ZN(n738) );
  XOR2_X1 U822 ( .A(G2078), .B(KEYINPUT25), .Z(n944) );
  NOR2_X1 U823 ( .A1(n944), .A2(n733), .ZN(n736) );
  NOR2_X1 U824 ( .A1(G1961), .A2(n734), .ZN(n735) );
  NOR2_X1 U825 ( .A1(n736), .A2(n735), .ZN(n743) );
  NOR2_X1 U826 ( .A1(G301), .A2(n743), .ZN(n737) );
  NOR2_X1 U827 ( .A1(n738), .A2(n737), .ZN(n748) );
  NOR2_X1 U828 ( .A1(G1966), .A2(n783), .ZN(n761) );
  NOR2_X1 U829 ( .A1(n751), .A2(G2084), .ZN(n759) );
  NOR2_X1 U830 ( .A1(n761), .A2(n759), .ZN(n739) );
  NAND2_X1 U831 ( .A1(G8), .A2(n739), .ZN(n741) );
  NOR2_X1 U832 ( .A1(n742), .A2(G168), .ZN(n745) );
  AND2_X1 U833 ( .A1(G301), .A2(n743), .ZN(n744) );
  NOR2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U835 ( .A(n518), .B(KEYINPUT31), .ZN(n747) );
  NOR2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U837 ( .A(n749), .B(KEYINPUT94), .ZN(n760) );
  INV_X1 U838 ( .A(G286), .ZN(n750) );
  INV_X1 U839 ( .A(G8), .ZN(n756) );
  NOR2_X1 U840 ( .A1(n751), .A2(G2090), .ZN(n753) );
  NOR2_X1 U841 ( .A1(G1971), .A2(n783), .ZN(n752) );
  NOR2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n754), .A2(G303), .ZN(n755) );
  OR2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U845 ( .A1(G8), .A2(n759), .ZN(n763) );
  NOR2_X1 U846 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n968) );
  INV_X1 U848 ( .A(n968), .ZN(n765) );
  NOR2_X1 U849 ( .A1(G1976), .A2(G288), .ZN(n770) );
  NOR2_X1 U850 ( .A1(G1971), .A2(G303), .ZN(n764) );
  NOR2_X1 U851 ( .A1(n770), .A2(n764), .ZN(n969) );
  OR2_X1 U852 ( .A1(n765), .A2(n969), .ZN(n766) );
  NOR2_X1 U853 ( .A1(n783), .A2(n767), .ZN(n768) );
  NOR2_X1 U854 ( .A1(KEYINPUT33), .A2(n768), .ZN(n769) );
  XNOR2_X1 U855 ( .A(G1981), .B(G305), .ZN(n989) );
  NAND2_X1 U856 ( .A1(n770), .A2(KEYINPUT33), .ZN(n771) );
  NOR2_X1 U857 ( .A1(n783), .A2(n771), .ZN(n772) );
  NOR2_X1 U858 ( .A1(n989), .A2(n772), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n775), .A2(n774), .ZN(n778) );
  NOR2_X1 U860 ( .A1(G2090), .A2(G303), .ZN(n776) );
  NAND2_X1 U861 ( .A1(G8), .A2(n776), .ZN(n777) );
  NAND2_X1 U862 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U863 ( .A1(n779), .A2(n783), .ZN(n785) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n780) );
  XNOR2_X1 U865 ( .A(KEYINPUT87), .B(n780), .ZN(n781) );
  XNOR2_X1 U866 ( .A(KEYINPUT24), .B(n781), .ZN(n782) );
  NOR2_X1 U867 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U868 ( .A1(G160), .A2(G40), .ZN(n787) );
  NOR2_X1 U869 ( .A1(n786), .A2(n787), .ZN(n826) );
  NAND2_X1 U870 ( .A1(G95), .A2(n893), .ZN(n789) );
  NAND2_X1 U871 ( .A1(G131), .A2(n896), .ZN(n788) );
  NAND2_X1 U872 ( .A1(n789), .A2(n788), .ZN(n793) );
  NAND2_X1 U873 ( .A1(G107), .A2(n627), .ZN(n791) );
  NAND2_X1 U874 ( .A1(G119), .A2(n889), .ZN(n790) );
  NAND2_X1 U875 ( .A1(n791), .A2(n790), .ZN(n792) );
  OR2_X1 U876 ( .A1(n793), .A2(n792), .ZN(n886) );
  NAND2_X1 U877 ( .A1(G1991), .A2(n886), .ZN(n802) );
  NAND2_X1 U878 ( .A1(G141), .A2(n896), .ZN(n795) );
  NAND2_X1 U879 ( .A1(G129), .A2(n889), .ZN(n794) );
  NAND2_X1 U880 ( .A1(n795), .A2(n794), .ZN(n798) );
  NAND2_X1 U881 ( .A1(n893), .A2(G105), .ZN(n796) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n796), .Z(n797) );
  NOR2_X1 U883 ( .A1(n798), .A2(n797), .ZN(n800) );
  NAND2_X1 U884 ( .A1(n627), .A2(G117), .ZN(n799) );
  NAND2_X1 U885 ( .A1(n800), .A2(n799), .ZN(n880) );
  NAND2_X1 U886 ( .A1(G1996), .A2(n880), .ZN(n801) );
  NAND2_X1 U887 ( .A1(n802), .A2(n801), .ZN(n924) );
  NAND2_X1 U888 ( .A1(n826), .A2(n924), .ZN(n818) );
  NAND2_X1 U889 ( .A1(G104), .A2(n893), .ZN(n804) );
  NAND2_X1 U890 ( .A1(G140), .A2(n896), .ZN(n803) );
  NAND2_X1 U891 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U892 ( .A(KEYINPUT34), .B(n805), .ZN(n810) );
  NAND2_X1 U893 ( .A1(G116), .A2(n627), .ZN(n807) );
  NAND2_X1 U894 ( .A1(G128), .A2(n889), .ZN(n806) );
  NAND2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U896 ( .A(KEYINPUT35), .B(n808), .Z(n809) );
  NOR2_X1 U897 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U898 ( .A(KEYINPUT36), .B(n811), .ZN(n881) );
  XNOR2_X1 U899 ( .A(KEYINPUT37), .B(G2067), .ZN(n824) );
  NOR2_X1 U900 ( .A1(n881), .A2(n824), .ZN(n925) );
  NAND2_X1 U901 ( .A1(n826), .A2(n925), .ZN(n822) );
  XNOR2_X1 U902 ( .A(G1986), .B(G290), .ZN(n973) );
  NAND2_X1 U903 ( .A1(n973), .A2(n826), .ZN(n812) );
  NAND2_X1 U904 ( .A1(n516), .A2(n812), .ZN(n829) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n886), .ZN(n813) );
  XOR2_X1 U906 ( .A(KEYINPUT97), .B(n813), .Z(n929) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n814) );
  XNOR2_X1 U908 ( .A(KEYINPUT96), .B(n814), .ZN(n815) );
  NOR2_X1 U909 ( .A1(n929), .A2(n815), .ZN(n816) );
  XOR2_X1 U910 ( .A(KEYINPUT98), .B(n816), .Z(n817) );
  NAND2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n819) );
  OR2_X1 U912 ( .A1(n880), .A2(G1996), .ZN(n921) );
  NAND2_X1 U913 ( .A1(n819), .A2(n921), .ZN(n820) );
  XNOR2_X1 U914 ( .A(n820), .B(KEYINPUT99), .ZN(n821) );
  XNOR2_X1 U915 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n881), .A2(n824), .ZN(n926) );
  NAND2_X1 U918 ( .A1(n825), .A2(n926), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n829), .A2(n828), .ZN(n832) );
  XOR2_X1 U921 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n830) );
  XNOR2_X1 U922 ( .A(KEYINPUT40), .B(n830), .ZN(n831) );
  XNOR2_X1 U923 ( .A(n832), .B(n831), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n915), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U926 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n834) );
  XOR2_X1 U928 ( .A(KEYINPUT103), .B(n834), .Z(n835) );
  NAND2_X1 U929 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U931 ( .A(G108), .ZN(G238) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  INV_X1 U935 ( .A(n839), .ZN(G319) );
  XNOR2_X1 U936 ( .A(G1996), .B(KEYINPUT106), .ZN(n849) );
  XOR2_X1 U937 ( .A(G1956), .B(G1961), .Z(n841) );
  XNOR2_X1 U938 ( .A(G1991), .B(G1976), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U940 ( .A(G1966), .B(G1971), .Z(n843) );
  XNOR2_X1 U941 ( .A(G1986), .B(G1981), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U943 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U944 ( .A(G2474), .B(KEYINPUT41), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(G229) );
  XNOR2_X1 U947 ( .A(n850), .B(KEYINPUT105), .ZN(n852) );
  XNOR2_X1 U948 ( .A(KEYINPUT104), .B(KEYINPUT43), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U950 ( .A(KEYINPUT42), .B(G2090), .Z(n854) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2072), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U953 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U954 ( .A(G2678), .B(G2096), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(n860) );
  XOR2_X1 U956 ( .A(G2078), .B(G2084), .Z(n859) );
  XNOR2_X1 U957 ( .A(n860), .B(n859), .ZN(G227) );
  NAND2_X1 U958 ( .A1(G100), .A2(n893), .ZN(n862) );
  NAND2_X1 U959 ( .A1(G112), .A2(n627), .ZN(n861) );
  NAND2_X1 U960 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n863), .B(KEYINPUT107), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G136), .A2(n896), .ZN(n864) );
  NAND2_X1 U963 ( .A1(n865), .A2(n864), .ZN(n868) );
  NAND2_X1 U964 ( .A1(n889), .A2(G124), .ZN(n866) );
  XOR2_X1 U965 ( .A(KEYINPUT44), .B(n866), .Z(n867) );
  NOR2_X1 U966 ( .A1(n868), .A2(n867), .ZN(G162) );
  XOR2_X1 U967 ( .A(KEYINPUT48), .B(KEYINPUT110), .Z(n870) );
  XNOR2_X1 U968 ( .A(KEYINPUT46), .B(KEYINPUT109), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(n879) );
  NAND2_X1 U970 ( .A1(G118), .A2(n627), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G130), .A2(n889), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U973 ( .A1(G106), .A2(n893), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G142), .A2(n896), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U976 ( .A(n875), .B(KEYINPUT45), .Z(n876) );
  NOR2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U978 ( .A(n879), .B(n878), .Z(n885) );
  XOR2_X1 U979 ( .A(n881), .B(n880), .Z(n883) );
  XNOR2_X1 U980 ( .A(G164), .B(G160), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n888) );
  XNOR2_X1 U983 ( .A(n886), .B(n928), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n901) );
  NAND2_X1 U985 ( .A1(G115), .A2(n627), .ZN(n891) );
  NAND2_X1 U986 ( .A1(G127), .A2(n889), .ZN(n890) );
  NAND2_X1 U987 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n892), .B(KEYINPUT47), .ZN(n895) );
  NAND2_X1 U989 ( .A1(G103), .A2(n893), .ZN(n894) );
  NAND2_X1 U990 ( .A1(n895), .A2(n894), .ZN(n899) );
  NAND2_X1 U991 ( .A1(n896), .A2(G139), .ZN(n897) );
  XOR2_X1 U992 ( .A(KEYINPUT108), .B(n897), .Z(n898) );
  NOR2_X1 U993 ( .A1(n899), .A2(n898), .ZN(n916) );
  XNOR2_X1 U994 ( .A(G162), .B(n916), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(n903) );
  XOR2_X1 U997 ( .A(KEYINPUT111), .B(n903), .Z(G395) );
  XNOR2_X1 U998 ( .A(G286), .B(n904), .ZN(n907) );
  XOR2_X1 U999 ( .A(n976), .B(n905), .Z(n906) );
  XNOR2_X1 U1000 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1001 ( .A(n908), .B(G171), .Z(n909) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n909), .ZN(G397) );
  NOR2_X1 U1003 ( .A1(G229), .A2(G227), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1005 ( .A1(G401), .A2(n911), .ZN(n912) );
  AND2_X1 U1006 ( .A1(G319), .A2(n912), .ZN(n914) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1008 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(G69), .ZN(G235) );
  INV_X1 U1011 ( .A(n915), .ZN(G223) );
  XNOR2_X1 U1012 ( .A(G2072), .B(n916), .ZN(n919) );
  XNOR2_X1 U1013 ( .A(G164), .B(G2078), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(n917), .B(KEYINPUT114), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1016 ( .A(n920), .B(KEYINPUT50), .ZN(n939) );
  XNOR2_X1 U1017 ( .A(G2090), .B(G162), .ZN(n922) );
  NAND2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(n923), .B(KEYINPUT51), .ZN(n937) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n927) );
  NAND2_X1 U1021 ( .A1(n927), .A2(n926), .ZN(n935) );
  NOR2_X1 U1022 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1023 ( .A(KEYINPUT112), .B(n930), .Z(n932) );
  XOR2_X1 U1024 ( .A(G160), .B(G2084), .Z(n931) );
  NOR2_X1 U1025 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1026 ( .A(n933), .B(KEYINPUT113), .ZN(n934) );
  NOR2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1028 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1029 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1030 ( .A(n940), .B(KEYINPUT52), .ZN(n941) );
  XNOR2_X1 U1031 ( .A(KEYINPUT55), .B(KEYINPUT115), .ZN(n962) );
  NAND2_X1 U1032 ( .A1(n941), .A2(n962), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(KEYINPUT116), .B(n942), .ZN(n943) );
  NAND2_X1 U1034 ( .A1(n943), .A2(G29), .ZN(n1025) );
  XOR2_X1 U1035 ( .A(G1996), .B(G32), .Z(n947) );
  XNOR2_X1 U1036 ( .A(n944), .B(KEYINPUT117), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(n945), .B(G27), .ZN(n946) );
  NAND2_X1 U1038 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1039 ( .A(n948), .B(KEYINPUT118), .ZN(n951) );
  XOR2_X1 U1040 ( .A(G1991), .B(G25), .Z(n949) );
  NAND2_X1 U1041 ( .A1(n949), .A2(G28), .ZN(n950) );
  NOR2_X1 U1042 ( .A1(n951), .A2(n950), .ZN(n955) );
  XNOR2_X1 U1043 ( .A(G2067), .B(G26), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(G33), .B(G2072), .ZN(n952) );
  NOR2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(n956), .B(KEYINPUT53), .ZN(n959) );
  XOR2_X1 U1048 ( .A(G2084), .B(G34), .Z(n957) );
  XNOR2_X1 U1049 ( .A(KEYINPUT54), .B(n957), .ZN(n958) );
  NAND2_X1 U1050 ( .A1(n959), .A2(n958), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(G35), .B(G2090), .ZN(n960) );
  NOR2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(n963), .B(n962), .ZN(n964) );
  NOR2_X1 U1054 ( .A1(G29), .A2(n964), .ZN(n965) );
  XNOR2_X1 U1055 ( .A(KEYINPUT119), .B(n965), .ZN(n966) );
  NAND2_X1 U1056 ( .A1(n966), .A2(G11), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(n967), .B(KEYINPUT120), .ZN(n1023) );
  INV_X1 U1058 ( .A(G16), .ZN(n1019) );
  XOR2_X1 U1059 ( .A(n1019), .B(KEYINPUT56), .Z(n995) );
  AND2_X1 U1060 ( .A1(G303), .A2(G1971), .ZN(n971) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n981) );
  XOR2_X1 U1063 ( .A(G301), .B(G1961), .Z(n975) );
  XNOR2_X1 U1064 ( .A(G1956), .B(G299), .ZN(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n979) );
  XOR2_X1 U1067 ( .A(G1348), .B(n976), .Z(n977) );
  XNOR2_X1 U1068 ( .A(KEYINPUT122), .B(n977), .ZN(n978) );
  NOR2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(KEYINPUT123), .B(n982), .ZN(n986) );
  XOR2_X1 U1072 ( .A(n983), .B(G1341), .Z(n984) );
  XNOR2_X1 U1073 ( .A(n984), .B(KEYINPUT124), .ZN(n985) );
  NAND2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(KEYINPUT125), .B(n987), .ZN(n993) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G168), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(n988), .B(KEYINPUT121), .ZN(n990) );
  NOR2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n991), .Z(n992) );
  NAND2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n1021) );
  XOR2_X1 U1082 ( .A(G1976), .B(G23), .Z(n997) );
  XOR2_X1 U1083 ( .A(G1971), .B(G22), .Z(n996) );
  NAND2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(G24), .B(G1986), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1087 ( .A(KEYINPUT58), .B(n1000), .Z(n1016) );
  XOR2_X1 U1088 ( .A(G1961), .B(G5), .Z(n1011) );
  XNOR2_X1 U1089 ( .A(G1348), .B(KEYINPUT59), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(n1001), .B(G4), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(G1981), .B(G6), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G1341), .B(G19), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(KEYINPUT126), .B(G1956), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(G20), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(KEYINPUT60), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(G21), .B(G1966), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1026), .ZN(G150) );
  INV_X1 U1110 ( .A(G150), .ZN(G311) );
endmodule

