//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT65), .Z(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n209), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT67), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g0026(.A1(new_n224), .A2(new_n225), .ZN(new_n227));
  AND2_X1   g0027(.A1(KEYINPUT66), .A2(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(KEYINPUT66), .A2(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NOR4_X1   g0033(.A1(new_n213), .A2(new_n226), .A3(new_n227), .A4(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G150), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n230), .A2(G33), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n252), .B1(new_n207), .B2(new_n201), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n231), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n257), .ZN(new_n261));
  INV_X1    g0061(.A(G50), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n262), .B1(new_n206), .B2(G20), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n261), .A2(new_n263), .B1(new_n262), .B2(new_n260), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT9), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G222), .A2(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G223), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n267), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n271), .B(new_n272), .C1(G77), .C2(new_n267), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT69), .B(G41), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n275), .B(new_n206), .C1(G45), .C2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  INV_X1    g0079(.A(G45), .ZN(new_n280));
  AOI21_X1  g0080(.A(G1), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n272), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G226), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n273), .A2(new_n278), .A3(new_n283), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n265), .A2(new_n266), .B1(G200), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G190), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n285), .B1(new_n266), .B2(new_n265), .C1(new_n286), .C2(new_n284), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n287), .B(KEYINPUT10), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n284), .A2(G179), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT70), .ZN(new_n290));
  INV_X1    g0090(.A(new_n265), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(new_n284), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n282), .A2(G244), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n278), .A2(new_n296), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n297), .A2(KEYINPUT71), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n267), .A2(G232), .ZN(new_n299));
  INV_X1    g0099(.A(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT3), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT3), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G33), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n299), .A2(new_n269), .B1(G107), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n267), .A2(G1698), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(new_n216), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n272), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n297), .A2(KEYINPUT71), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n298), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G200), .ZN(new_n311));
  INV_X1    g0111(.A(new_n254), .ZN(new_n312));
  OR2_X1    g0112(.A1(KEYINPUT66), .A2(G20), .ZN(new_n313));
  NAND2_X1  g0113(.A1(KEYINPUT66), .A2(G20), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n312), .A2(new_n251), .B1(new_n315), .B2(G77), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT72), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT15), .B(G87), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n317), .B1(new_n253), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n316), .A2(KEYINPUT72), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n257), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n261), .A2(new_n322), .B1(new_n202), .B2(new_n260), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n311), .B(new_n325), .C1(new_n286), .C2(new_n310), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n310), .A2(G179), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n310), .A2(new_n292), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n295), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n254), .B1(new_n206), .B2(G20), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n331), .A2(new_n261), .B1(new_n260), .B2(new_n254), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT78), .ZN(new_n334));
  INV_X1    g0134(.A(G58), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(new_n215), .ZN(new_n336));
  NOR2_X1   g0136(.A1(G58), .A2(G68), .ZN(new_n337));
  OAI21_X1  g0137(.A(G20), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n251), .A2(G159), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT16), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(G20), .B1(new_n301), .B2(new_n303), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT7), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT7), .B1(new_n304), .B2(new_n230), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT74), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n347), .B(new_n349), .C1(new_n315), .C2(new_n267), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(G68), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT75), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n349), .B1(new_n315), .B2(new_n267), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT74), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(new_n350), .A3(new_n345), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(KEYINPUT75), .A3(G68), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n343), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT76), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n344), .B2(KEYINPUT7), .ZN(new_n361));
  OAI211_X1 g0161(.A(KEYINPUT76), .B(new_n349), .C1(new_n267), .C2(G20), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n315), .A2(new_n349), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT77), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n301), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n300), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n303), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n340), .B1(new_n370), .B2(G68), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n257), .B1(new_n371), .B2(KEYINPUT16), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n334), .B1(new_n359), .B2(new_n372), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n355), .A2(KEYINPUT74), .B1(KEYINPUT7), .B2(new_n344), .ZN(new_n374));
  AOI211_X1 g0174(.A(new_n353), .B(new_n215), .C1(new_n374), .C2(new_n350), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT75), .B1(new_n357), .B2(G68), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n342), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n257), .ZN(new_n378));
  INV_X1    g0178(.A(new_n340), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n361), .A2(new_n362), .B1(new_n368), .B2(new_n364), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(new_n215), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n378), .B1(new_n381), .B2(new_n341), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n377), .A2(KEYINPUT78), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n333), .B1(new_n373), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n282), .A2(G232), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n278), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n386), .B(KEYINPUT79), .ZN(new_n387));
  INV_X1    g0187(.A(G226), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G1698), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(G223), .B2(G1698), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n390), .A2(new_n304), .B1(new_n300), .B2(new_n217), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n272), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n393), .A2(G179), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n278), .A2(new_n392), .A3(new_n385), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n387), .A2(new_n394), .B1(new_n292), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT18), .B1(new_n384), .B2(new_n397), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n377), .A2(KEYINPUT78), .A3(new_n382), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT78), .B1(new_n377), .B2(new_n382), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n332), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT18), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n402), .A3(new_n396), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n387), .A2(new_n286), .A3(new_n392), .ZN(new_n404));
  INV_X1    g0204(.A(G200), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n395), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n332), .B(new_n407), .C1(new_n399), .C2(new_n400), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT17), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n384), .A2(KEYINPUT17), .A3(new_n407), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n398), .A2(new_n403), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n251), .A2(G50), .B1(G20), .B2(new_n215), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n253), .B2(new_n202), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n414), .A2(new_n257), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n415), .A2(KEYINPUT11), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(KEYINPUT11), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT12), .B1(new_n259), .B2(G68), .ZN(new_n418));
  OR3_X1    g0218(.A1(new_n259), .A2(KEYINPUT12), .A3(G68), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n215), .B1(new_n206), .B2(G20), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n418), .A2(new_n419), .B1(new_n261), .B2(new_n420), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n416), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n272), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n267), .A2(new_n269), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT73), .B1(new_n425), .B2(new_n388), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT73), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n267), .A2(new_n427), .A3(G226), .A4(new_n269), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n299), .A2(G1698), .B1(G33), .B2(G97), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n424), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n282), .A2(G238), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n278), .A2(new_n432), .ZN(new_n433));
  OR3_X1    g0233(.A1(new_n431), .A2(KEYINPUT13), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT13), .B1(new_n431), .B2(new_n433), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT14), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(G169), .ZN(new_n438));
  INV_X1    g0238(.A(G179), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(new_n436), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n437), .B1(new_n436), .B2(G169), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n423), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n436), .A2(G200), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(new_n422), .C1(new_n286), .C2(new_n436), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n330), .A2(new_n412), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT80), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n279), .A2(KEYINPUT69), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT69), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G41), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT5), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n280), .A2(G1), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n447), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(KEYINPUT80), .B(new_n452), .C1(new_n276), .C2(KEYINPUT5), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n279), .A2(KEYINPUT5), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n454), .A2(new_n275), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n218), .A2(new_n269), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(G257), .B2(new_n269), .ZN(new_n459));
  INV_X1    g0259(.A(G294), .ZN(new_n460));
  OAI22_X1  g0260(.A1(new_n459), .A2(new_n304), .B1(new_n300), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n272), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(G264), .A3(new_n424), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT88), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT88), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n464), .A2(new_n467), .A3(G264), .A4(new_n424), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n463), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n463), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n465), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n469), .A2(G179), .B1(new_n471), .B2(G169), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  OR2_X1    g0273(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n475));
  INV_X1    g0275(.A(G107), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n260), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n474), .B(new_n475), .C1(new_n477), .C2(KEYINPUT87), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(KEYINPUT87), .ZN(new_n479));
  XNOR2_X1  g0279(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n206), .A2(G33), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n259), .A2(new_n481), .A3(new_n231), .A4(new_n256), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G107), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT84), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(KEYINPUT24), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n230), .A2(new_n267), .A3(G87), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT22), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT22), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n230), .A2(new_n267), .A3(new_n491), .A4(G87), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G116), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(G20), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT82), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(KEYINPUT82), .B(KEYINPUT23), .C1(new_n207), .C2(G107), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT83), .ZN(new_n501));
  NOR2_X1   g0301(.A1(KEYINPUT23), .A2(G107), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n501), .B1(new_n315), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n501), .B(new_n502), .C1(new_n228), .C2(new_n229), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n500), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n488), .B1(new_n493), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n490), .A2(new_n492), .ZN(new_n508));
  OR2_X1    g0308(.A1(new_n503), .A2(new_n505), .ZN(new_n509));
  XNOR2_X1  g0309(.A(KEYINPUT84), .B(KEYINPUT24), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n500), .A4(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(new_n257), .A3(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(KEYINPUT85), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT85), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n508), .A2(new_n509), .A3(new_n500), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n378), .B1(new_n515), .B2(new_n488), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n516), .B2(new_n511), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n486), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n473), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n512), .A2(KEYINPUT85), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n516), .A2(new_n514), .A3(new_n511), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI22_X1  g0322(.A1(new_n469), .A2(G200), .B1(G190), .B2(new_n471), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n523), .A3(new_n486), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G283), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n300), .A2(G97), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n230), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G116), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n256), .A2(new_n231), .B1(G20), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT20), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n528), .A2(KEYINPUT20), .A3(new_n530), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n259), .A2(G116), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n483), .B2(G116), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n464), .A2(G270), .A3(new_n424), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n267), .A2(G257), .A3(new_n269), .ZN(new_n540));
  INV_X1    g0340(.A(G303), .ZN(new_n541));
  INV_X1    g0341(.A(G264), .ZN(new_n542));
  OAI221_X1 g0342(.A(new_n540), .B1(new_n541), .B2(new_n267), .C1(new_n306), .C2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n439), .B1(new_n543), .B2(new_n272), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n538), .A2(new_n457), .A3(new_n539), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n272), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n539), .A2(new_n546), .A3(new_n457), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n292), .B1(new_n535), .B2(new_n537), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT21), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n549), .B1(new_n547), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OR2_X1    g0352(.A1(new_n547), .A2(new_n286), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n538), .B1(new_n547), .B2(G200), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n318), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(new_n259), .ZN(new_n557));
  NOR2_X1   g0357(.A1(G97), .A2(G107), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n217), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  INV_X1    g0360(.A(G97), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n560), .A2(new_n300), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n559), .B1(new_n562), .B2(new_n315), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n313), .A2(G33), .A3(G97), .A4(new_n314), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n560), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n230), .A2(new_n267), .A3(G68), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n557), .B1(new_n567), .B2(new_n257), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n483), .A2(new_n556), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n453), .A2(new_n218), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n452), .A2(new_n274), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n424), .A3(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n301), .A2(new_n303), .A3(G238), .A4(new_n269), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n494), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n301), .A2(new_n303), .A3(G244), .A4(G1698), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT81), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n267), .A2(KEYINPUT81), .A3(G244), .A4(G1698), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n439), .B(new_n573), .C1(new_n580), .C2(new_n424), .ZN(new_n581));
  INV_X1    g0381(.A(new_n573), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n579), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(new_n494), .A3(new_n574), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n582), .B1(new_n584), .B2(new_n272), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n570), .B(new_n581), .C1(new_n585), .C2(G169), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n482), .A2(new_n217), .ZN(new_n587));
  AOI211_X1 g0387(.A(new_n557), .B(new_n587), .C1(new_n567), .C2(new_n257), .ZN(new_n588));
  OAI211_X1 g0388(.A(G190), .B(new_n573), .C1(new_n580), .C2(new_n424), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n588), .B(new_n589), .C1(new_n585), .C2(new_n405), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n260), .A2(new_n561), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n482), .B2(new_n561), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n251), .A2(G77), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT6), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n596), .A2(new_n561), .A3(G107), .ZN(new_n597));
  XNOR2_X1  g0397(.A(G97), .B(G107), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n597), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n595), .B1(new_n599), .B2(new_n230), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n370), .B2(G107), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n594), .B1(new_n601), .B2(new_n378), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n464), .A2(G257), .A3(new_n424), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n301), .A2(new_n303), .A3(G250), .A4(G1698), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n301), .A2(new_n303), .A3(G244), .A4(new_n269), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT4), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n526), .B(new_n605), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n272), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n457), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n292), .B1(new_n604), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n603), .A2(new_n439), .A3(new_n457), .A4(new_n610), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n602), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(G200), .B1(new_n604), .B2(new_n611), .ZN(new_n615));
  INV_X1    g0415(.A(new_n600), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n380), .B2(new_n476), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n593), .B1(new_n617), .B2(new_n257), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n603), .A2(G190), .A3(new_n457), .A4(new_n610), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n615), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n591), .A2(new_n614), .A3(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n446), .A2(new_n525), .A3(new_n555), .A4(new_n621), .ZN(G372));
  NAND2_X1  g0422(.A1(new_n442), .A2(new_n329), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n444), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n410), .A2(new_n411), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n398), .B(new_n403), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n626), .A2(new_n288), .B1(new_n290), .B2(new_n293), .ZN(new_n627));
  INV_X1    g0427(.A(new_n586), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n602), .A2(new_n613), .A3(new_n612), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(new_n591), .A3(KEYINPUT26), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n586), .A2(new_n590), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n631), .B1(new_n614), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n628), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT90), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT89), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n614), .A2(new_n620), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n524), .A2(new_n638), .A3(new_n591), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n552), .B1(new_n473), .B2(new_n518), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n552), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n485), .B1(new_n520), .B2(new_n521), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(new_n472), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n644), .A2(new_n621), .A3(KEYINPUT89), .A4(new_n524), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n636), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n446), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n627), .A2(new_n648), .ZN(G369));
  NAND3_X1  g0449(.A1(new_n230), .A2(new_n206), .A3(G13), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G343), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n538), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n555), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n642), .B2(new_n657), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  INV_X1    g0460(.A(new_n656), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n525), .B1(new_n643), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n519), .B2(new_n661), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n642), .A2(new_n656), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n525), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n473), .A2(new_n518), .A3(new_n661), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n664), .A2(new_n668), .ZN(G399));
  NOR2_X1   g0469(.A1(new_n559), .A2(G116), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT91), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n210), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(new_n277), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n672), .A2(new_n675), .A3(G1), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n232), .B2(new_n675), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n656), .B1(new_n636), .B2(new_n646), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g0480(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n644), .A2(new_n621), .A3(new_n524), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n656), .B1(new_n682), .B2(new_n634), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n680), .A2(new_n681), .B1(KEYINPUT29), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n585), .A2(new_n462), .A3(new_n544), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n539), .A2(new_n457), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n466), .A2(new_n468), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n604), .A2(new_n611), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n689), .A2(G179), .A3(new_n585), .ZN(new_n693));
  INV_X1    g0493(.A(new_n469), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(new_n694), .A3(new_n547), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n690), .A2(new_n691), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n692), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n656), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT31), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n525), .A2(new_n555), .A3(new_n621), .A4(new_n661), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n697), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n684), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n678), .B1(new_n705), .B2(G1), .ZN(G364));
  INV_X1    g0506(.A(G13), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n315), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n206), .B1(new_n708), .B2(G45), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n674), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n660), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(G330), .B2(new_n659), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n210), .A2(new_n267), .ZN(new_n714));
  INV_X1    g0514(.A(G355), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n714), .A2(new_n715), .B1(G116), .B2(new_n210), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n210), .A2(new_n304), .ZN(new_n717));
  INV_X1    g0517(.A(new_n232), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n717), .B1(new_n280), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n249), .A2(G45), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n716), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n207), .B1(KEYINPUT93), .B2(new_n292), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n292), .A2(KEYINPUT93), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n231), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n711), .B1(new_n721), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n230), .A2(G190), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n405), .A2(G179), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G283), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n230), .A2(new_n439), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G190), .A2(G200), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G311), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G179), .A2(G200), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n230), .B1(G190), .B2(new_n740), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n738), .A2(new_n739), .B1(new_n741), .B2(new_n460), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n731), .A2(G179), .A3(G200), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  XNOR2_X1  g0544(.A(KEYINPUT33), .B(G317), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n735), .B(new_n742), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n731), .A2(new_n740), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n747), .A2(KEYINPUT94), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(KEYINPUT94), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G329), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n736), .A2(G190), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n405), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G326), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n732), .A2(G20), .A3(G190), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n756), .A2(KEYINPUT96), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(KEYINPUT96), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n304), .B1(new_n759), .B2(new_n541), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n753), .A2(G200), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n760), .B1(G322), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n746), .A2(new_n752), .A3(new_n755), .A4(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G159), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n750), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT95), .B(KEYINPUT32), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n765), .B(new_n766), .Z(new_n767));
  INV_X1    g0567(.A(new_n754), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n267), .B1(new_n561), .B2(new_n741), .C1(new_n768), .C2(new_n262), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(G58), .B2(new_n761), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n202), .A2(new_n738), .B1(new_n733), .B2(new_n476), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n759), .A2(new_n217), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n771), .B(new_n772), .C1(G68), .C2(new_n744), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n763), .B1(new_n767), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n730), .B1(new_n775), .B2(new_n724), .ZN(new_n776));
  INV_X1    g0576(.A(new_n727), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n659), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n713), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(G396));
  NOR2_X1   g0580(.A1(new_n329), .A2(new_n656), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n326), .B1(new_n325), .B2(new_n661), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(new_n782), .B2(new_n329), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n680), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n641), .A2(new_n645), .ZN(new_n786));
  AOI21_X1  g0586(.A(KEYINPUT26), .B1(new_n629), .B2(new_n591), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n614), .A2(new_n632), .A3(new_n631), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n586), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n635), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n634), .A2(KEYINPUT90), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n661), .B(new_n783), .C1(new_n786), .C2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n704), .B1(new_n785), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n711), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n785), .A2(new_n704), .A3(new_n793), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n711), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n724), .A2(new_n725), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(new_n202), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n724), .ZN(new_n801));
  INV_X1    g0601(.A(new_n738), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n744), .A2(G150), .B1(new_n802), .B2(G159), .ZN(new_n803));
  INV_X1    g0603(.A(new_n761), .ZN(new_n804));
  INV_X1    g0604(.A(G143), .ZN(new_n805));
  INV_X1    g0605(.A(G137), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n803), .B1(new_n804), .B2(new_n805), .C1(new_n806), .C2(new_n768), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT34), .ZN(new_n808));
  INV_X1    g0608(.A(new_n759), .ZN(new_n809));
  INV_X1    g0609(.A(new_n741), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n809), .A2(G50), .B1(G58), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n733), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G68), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n811), .A2(new_n267), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G132), .B2(new_n751), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n761), .A2(G294), .B1(G97), .B2(new_n810), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n817), .A2(KEYINPUT99), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(KEYINPUT99), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n750), .A2(new_n739), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n304), .B1(new_n217), .B2(new_n733), .C1(new_n759), .C2(new_n476), .ZN(new_n821));
  NOR4_X1   g0621(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n754), .A2(G303), .B1(new_n802), .B2(G116), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n743), .A2(KEYINPUT97), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n743), .A2(KEYINPUT97), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n823), .B1(new_n826), .B2(new_n734), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT98), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n808), .A2(new_n815), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n800), .B1(new_n801), .B2(new_n829), .C1(new_n783), .C2(new_n726), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n797), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G384));
  NOR2_X1   g0632(.A1(new_n708), .A2(new_n206), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n422), .A2(new_n661), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n445), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n442), .B(new_n444), .C1(new_n422), .C2(new_n661), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n784), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n703), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n340), .B1(new_n354), .B2(new_n358), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n257), .B1(new_n840), .B2(KEYINPUT16), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n359), .B1(new_n841), .B2(KEYINPUT103), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n379), .B1(new_n375), .B2(new_n376), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n378), .B1(new_n843), .B2(new_n341), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT103), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n333), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(new_n654), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n412), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n377), .B1(new_n844), .B2(new_n845), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n841), .A2(KEYINPUT103), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n332), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n853), .A2(new_n396), .B1(new_n384), .B2(new_n407), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n653), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n850), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n408), .B1(new_n384), .B2(new_n397), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n850), .B1(new_n384), .B2(new_n654), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(KEYINPUT38), .B(new_n849), .C1(new_n856), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n408), .B1(new_n847), .B2(new_n397), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT37), .B1(new_n862), .B2(new_n848), .ZN(new_n863));
  INV_X1    g0663(.A(new_n859), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT38), .B1(new_n865), .B2(new_n849), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n839), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT107), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT40), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n853), .A2(new_n396), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n855), .A2(new_n872), .A3(new_n408), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n859), .B1(new_n873), .B2(KEYINPUT37), .ZN(new_n874));
  INV_X1    g0674(.A(new_n849), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n838), .B1(new_n876), .B2(new_n860), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT107), .B1(new_n877), .B2(KEYINPUT40), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT105), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n384), .A2(new_n654), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT37), .B1(new_n857), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT104), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n857), .B2(new_n858), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT37), .B1(new_n401), .B2(new_n653), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n401), .A2(new_n396), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n884), .A2(KEYINPUT104), .A3(new_n885), .A4(new_n408), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n881), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n412), .A2(new_n880), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n879), .B1(new_n889), .B2(new_n871), .ZN(new_n890));
  AOI211_X1 g0690(.A(KEYINPUT105), .B(KEYINPUT38), .C1(new_n887), .C2(new_n888), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n860), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n838), .A2(new_n869), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n870), .A2(new_n878), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n446), .A2(new_n703), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  INV_X1    g0697(.A(G330), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT108), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n781), .B1(new_n679), .B2(new_n783), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n835), .A2(new_n836), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT102), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n781), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n903), .B1(new_n793), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT102), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n904), .B(new_n908), .C1(new_n866), .C2(new_n861), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n398), .A2(new_n403), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n654), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n860), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n889), .A2(new_n871), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT105), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n889), .A2(new_n879), .A3(new_n871), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n913), .B1(new_n876), .B2(new_n860), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT106), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n863), .A2(new_n864), .B1(new_n412), .B2(new_n848), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT39), .B1(new_n921), .B2(KEYINPUT38), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n890), .B2(new_n891), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT39), .B1(new_n861), .B2(new_n866), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT106), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n920), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n442), .A2(new_n656), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n912), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n684), .A2(new_n446), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n931), .A2(new_n627), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n930), .B(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n833), .B1(new_n901), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n901), .B2(new_n933), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n315), .A2(G1), .A3(G13), .A4(G116), .ZN(new_n936));
  INV_X1    g0736(.A(new_n599), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n937), .B2(KEYINPUT35), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(KEYINPUT35), .B2(new_n937), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT100), .Z(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(KEYINPUT36), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(KEYINPUT36), .ZN(new_n943));
  OAI21_X1  g0743(.A(G77), .B1(new_n335), .B2(new_n215), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n944), .A2(new_n232), .B1(G50), .B2(new_n215), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(G1), .A3(new_n707), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT101), .Z(new_n947));
  NAND4_X1  g0747(.A1(new_n935), .A2(new_n942), .A3(new_n943), .A4(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT109), .Z(G367));
  OAI221_X1 g0749(.A(new_n728), .B1(new_n210), .B2(new_n318), .C1(new_n241), .C2(new_n717), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT111), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n952), .A2(new_n953), .A3(new_n798), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n661), .A2(new_n588), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(new_n586), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n591), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n541), .A2(new_n804), .B1(new_n768), .B2(new_n739), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n733), .A2(new_n561), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n738), .A2(new_n734), .B1(new_n741), .B2(new_n476), .ZN(new_n961));
  NOR4_X1   g0761(.A1(new_n959), .A2(new_n267), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n826), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT46), .B1(new_n759), .B2(new_n529), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n759), .A2(KEYINPUT46), .A3(new_n529), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n963), .A2(G294), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(G317), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n962), .B(new_n966), .C1(new_n967), .C2(new_n750), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n267), .B1(new_n202), .B2(new_n733), .C1(new_n768), .C2(new_n805), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G150), .B2(new_n761), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n963), .A2(G159), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n751), .A2(G137), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n741), .A2(new_n215), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n335), .B2(new_n759), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G50), .B2(new_n802), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n970), .A2(new_n971), .A3(new_n972), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n968), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT47), .Z(new_n979));
  OAI221_X1 g0779(.A(new_n954), .B1(new_n777), .B2(new_n958), .C1(new_n979), .C2(new_n801), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n638), .B1(new_n618), .B2(new_n661), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n629), .A2(new_n656), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n668), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT44), .Z(new_n986));
  NOR2_X1   g0786(.A1(new_n668), .A2(new_n984), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n664), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(KEYINPUT110), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n989), .B(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n666), .B1(new_n663), .B2(new_n665), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(new_n660), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n705), .A2(new_n994), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n705), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n674), .B(KEYINPUT41), .Z(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n710), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n983), .A2(new_n525), .A3(new_n665), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n614), .B1(new_n981), .B2(new_n519), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n1001), .A2(KEYINPUT42), .B1(new_n661), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(KEYINPUT42), .B2(new_n1001), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT43), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n958), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1005), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n664), .A2(new_n983), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n980), .B1(new_n1000), .B2(new_n1012), .ZN(G387));
  OR2_X1    g0813(.A1(new_n663), .A2(new_n777), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n238), .A2(new_n280), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1015), .A2(new_n717), .B1(new_n672), .B2(new_n714), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n254), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT50), .B1(new_n254), .B2(G50), .ZN(new_n1018));
  AOI21_X1  g0818(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n672), .A2(new_n1017), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1016), .A2(new_n1020), .B1(new_n476), .B2(new_n673), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n711), .B1(new_n1021), .B2(new_n729), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n741), .A2(new_n318), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n809), .A2(G77), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n215), .B2(new_n738), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1023), .B(new_n1025), .C1(new_n312), .C2(new_n744), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n754), .A2(G159), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n304), .B(new_n960), .C1(G50), .C2(new_n761), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n751), .A2(G150), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n751), .A2(G326), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n267), .B1(new_n812), .B2(G116), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n759), .A2(new_n460), .B1(new_n734), .B2(new_n741), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n754), .A2(G322), .B1(new_n802), .B2(G303), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n967), .B2(new_n804), .C1(new_n826), .C2(new_n739), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n1036), .B2(new_n1035), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1031), .B(new_n1032), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1030), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1022), .B1(new_n1042), .B2(new_n724), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n994), .A2(new_n710), .B1(new_n1014), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n995), .A2(new_n674), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n705), .A2(new_n994), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(G393));
  AND3_X1   g0847(.A1(new_n246), .A2(new_n210), .A3(new_n304), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n728), .B1(new_n561), .B2(new_n210), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n711), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G311), .A2(new_n761), .B1(new_n754), .B2(G317), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT52), .Z(new_n1052));
  OAI21_X1  g0852(.A(new_n304), .B1(new_n733), .B2(new_n476), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n759), .A2(new_n734), .B1(new_n529), .B2(new_n741), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(G294), .C2(new_n802), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n963), .A2(G303), .B1(new_n751), .B2(G322), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1052), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n826), .A2(new_n262), .B1(new_n254), .B2(new_n738), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT113), .Z(new_n1059));
  INV_X1    g0859(.A(G150), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1060), .A2(new_n768), .B1(new_n804), .B2(new_n764), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT51), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1061), .A2(new_n1062), .B1(G77), .B2(new_n810), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1059), .B(new_n1063), .C1(new_n1062), .C2(new_n1061), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n267), .B1(new_n217), .B2(new_n733), .C1(new_n759), .C2(new_n215), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n751), .B2(G143), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT112), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1057), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1050), .B1(new_n1068), .B2(new_n724), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n777), .B2(new_n983), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n989), .B(new_n664), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n996), .A2(new_n674), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1071), .A2(new_n995), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1070), .B1(new_n709), .B2(new_n1071), .C1(new_n1072), .C2(new_n1073), .ZN(G390));
  OAI21_X1  g0874(.A(KEYINPUT114), .B1(new_n906), .B2(new_n929), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT114), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1076), .B(new_n928), .C1(new_n902), .C2(new_n903), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n920), .A2(new_n926), .A3(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n704), .A2(new_n783), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n903), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n892), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n781), .B1(new_n683), .B2(new_n326), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n928), .B1(new_n903), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1079), .A2(new_n1082), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1082), .B1(new_n1079), .B2(new_n1087), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n710), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n798), .B1(new_n254), .B2(new_n799), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G128), .A2(new_n754), .B1(new_n761), .B2(G132), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT54), .B(G143), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT116), .Z(new_n1095));
  AOI21_X1  g0895(.A(new_n304), .B1(new_n1095), .B2(new_n802), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n812), .A2(G50), .B1(new_n810), .B2(G159), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1093), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n759), .A2(new_n1060), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT53), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n806), .B2(new_n826), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1098), .B(new_n1101), .C1(G125), .C2(new_n751), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT117), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n768), .A2(new_n734), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n804), .A2(new_n529), .ZN(new_n1105));
  NOR4_X1   g0905(.A1(new_n1104), .A2(new_n1105), .A3(new_n267), .A4(new_n772), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n813), .B1(new_n202), .B2(new_n741), .C1(new_n561), .C2(new_n738), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n963), .B2(G107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1106), .B(new_n1108), .C1(new_n460), .C2(new_n750), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1111), .A2(KEYINPUT118), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n724), .B1(new_n1111), .B2(KEYINPUT118), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1092), .B1(new_n1112), .B2(new_n1113), .C1(new_n927), .C2(new_n726), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1091), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1082), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n923), .A2(new_n925), .A3(new_n924), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n925), .B1(new_n923), .B2(new_n924), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1116), .B1(new_n1120), .B2(new_n1086), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1079), .A2(new_n1082), .A3(new_n1087), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n704), .A2(new_n446), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n932), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n704), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n903), .B1(new_n1125), .B2(new_n784), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1082), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n902), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1082), .A2(new_n1084), .A3(new_n1126), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1124), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1121), .A2(new_n1122), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT115), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1121), .A2(KEYINPUT115), .A3(new_n1131), .A4(new_n1122), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n932), .A2(new_n1123), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n675), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1115), .B1(new_n1136), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(G378));
  NOR2_X1   g0943(.A1(new_n277), .A2(new_n267), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1024), .A2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT119), .Z(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n335), .B2(new_n733), .C1(new_n734), .C2(new_n750), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT120), .Z(new_n1148));
  OAI221_X1 g0948(.A(new_n974), .B1(new_n738), .B2(new_n318), .C1(new_n561), .C2(new_n743), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n476), .A2(new_n804), .B1(new_n768), .B2(new_n529), .ZN(new_n1150));
  OR3_X1    g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT58), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(G33), .A2(G41), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1144), .A2(G50), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(G124), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1155), .B1(new_n764), .B2(new_n733), .C1(new_n750), .C2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n809), .A2(new_n1095), .B1(G132), .B2(new_n744), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G125), .A2(new_n754), .B1(new_n761), .B2(G128), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n802), .A2(G137), .B1(new_n810), .B2(G150), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1158), .B1(KEYINPUT59), .B2(new_n1162), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1156), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1153), .A2(new_n1154), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT121), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n801), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n1167), .B2(new_n1166), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n798), .B1(new_n262), .B2(new_n799), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n291), .A2(new_n654), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n295), .B(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1169), .B(new_n1170), .C1(new_n726), .C2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n930), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n898), .B1(new_n892), .B2(new_n893), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT122), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n868), .B1(new_n867), .B2(new_n869), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n877), .A2(KEYINPUT107), .A3(KEYINPUT40), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1178), .B(new_n1179), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n870), .A2(new_n878), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1179), .B1(new_n1184), .B2(new_n1178), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1174), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1183), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n1179), .A3(new_n1178), .A4(new_n1186), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1177), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1178), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(KEYINPUT122), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1192), .A2(new_n1182), .A3(new_n1174), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1193), .A2(new_n930), .A3(new_n1188), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1190), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1176), .B1(new_n1196), .B2(new_n710), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT115), .B1(new_n1090), .B2(new_n1131), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1135), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1139), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1200), .B2(new_n1196), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1124), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1190), .A2(KEYINPUT57), .A3(new_n1194), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n674), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1197), .B1(new_n1201), .B2(new_n1204), .ZN(G375));
  NAND3_X1  g1005(.A1(new_n1124), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1140), .A2(new_n999), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n903), .A2(new_n725), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n724), .A2(G68), .A3(new_n725), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n304), .B1(new_n202), .B2(new_n733), .C1(new_n768), .C2(new_n460), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G283), .B2(new_n761), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n963), .A2(G116), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n751), .A2(G303), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n738), .A2(new_n476), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1023), .B(new_n1214), .C1(new_n809), .C2(G97), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n751), .A2(G128), .B1(G159), .B2(new_n809), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT123), .Z(new_n1218));
  NAND2_X1  g1018(.A1(new_n963), .A2(new_n1095), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n738), .A2(new_n1060), .B1(new_n741), .B2(new_n262), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n304), .B(new_n1220), .C1(G58), .C2(new_n812), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G132), .A2(new_n754), .B1(new_n761), .B2(G137), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1219), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1216), .B1(new_n1218), .B2(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n798), .B(new_n1209), .C1(new_n1224), .C2(new_n724), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1138), .A2(new_n710), .B1(new_n1208), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1207), .A2(new_n1226), .ZN(G381));
  NOR4_X1   g1027(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1228));
  INV_X1    g1028(.A(G387), .ZN(new_n1229));
  INV_X1    g1029(.A(G381), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1228), .A2(new_n1142), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  OR2_X1    g1031(.A1(G375), .A2(new_n1231), .ZN(G407));
  NAND3_X1  g1032(.A1(new_n1142), .A2(G213), .A3(new_n655), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G407), .B(G213), .C1(G375), .C2(new_n1233), .ZN(G409));
  OAI211_X1 g1034(.A(G378), .B(new_n1197), .C1(new_n1201), .C2(new_n1204), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1193), .A2(new_n930), .A3(new_n1188), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n930), .B1(new_n1193), .B2(new_n1188), .ZN(new_n1237));
  OAI21_X1  g1037(.A(KEYINPUT124), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT124), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1190), .A2(new_n1239), .A3(new_n1194), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1240), .A3(new_n710), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1175), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1202), .A2(new_n998), .A3(new_n1195), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1142), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1235), .A2(new_n1244), .B1(G213), .B2(new_n655), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT126), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1140), .A2(KEYINPUT60), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1247), .A2(new_n1206), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1206), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n674), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1226), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n831), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(G384), .A3(new_n1226), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n655), .A2(G213), .A3(G2897), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1245), .A2(new_n1246), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1246), .B2(new_n1245), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(G393), .B(new_n779), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(G390), .B(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(new_n1229), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT61), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1235), .A2(new_n1244), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n655), .A2(G213), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n1255), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1266), .B1(new_n1270), .B2(KEYINPUT63), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT63), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1269), .A2(KEYINPUT125), .A3(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT125), .B1(new_n1269), .B2(new_n1272), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1261), .B(new_n1271), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT61), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  AND4_X1   g1078(.A1(KEYINPUT62), .A2(new_n1267), .A3(new_n1255), .A4(new_n1268), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT62), .B1(new_n1245), .B2(new_n1255), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1278), .B(KEYINPUT127), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1264), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1269), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1245), .A2(KEYINPUT62), .A3(new_n1255), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT127), .B1(new_n1287), .B2(new_n1278), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1275), .B1(new_n1283), .B2(new_n1288), .ZN(G405));
  NAND2_X1  g1089(.A1(G375), .A2(new_n1142), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1235), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(new_n1255), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(new_n1282), .ZN(G402));
endmodule


