

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737;

  XNOR2_X1 U368 ( .A(n367), .B(n366), .ZN(n570) );
  NOR2_X1 U369 ( .A1(n589), .A2(n512), .ZN(n375) );
  INV_X1 U370 ( .A(n650), .ZN(n589) );
  NOR2_X1 U371 ( .A1(n696), .A2(G902), .ZN(n440) );
  XOR2_X1 U372 ( .A(n690), .B(n689), .Z(n346) );
  NAND2_X2 U373 ( .A1(n520), .A2(n661), .ZN(n553) );
  NOR2_X1 U374 ( .A1(n413), .A2(n411), .ZN(n594) );
  XNOR2_X2 U375 ( .A(n531), .B(KEYINPUT1), .ZN(n653) );
  OR2_X2 U376 ( .A1(n690), .A2(n597), .ZN(n370) );
  XNOR2_X2 U377 ( .A(n422), .B(n421), .ZN(n716) );
  AND2_X1 U378 ( .A1(n580), .A2(n734), .ZN(n582) );
  AND2_X1 U379 ( .A1(n563), .A2(n564), .ZN(n367) );
  XOR2_X1 U380 ( .A(G143), .B(G128), .Z(n457) );
  NOR2_X1 U381 ( .A1(n547), .A2(KEYINPUT104), .ZN(n415) );
  NOR2_X1 U382 ( .A1(n403), .A2(n476), .ZN(n402) );
  INV_X1 U383 ( .A(n404), .ZN(n403) );
  XOR2_X1 U384 ( .A(G137), .B(G140), .Z(n487) );
  INV_X1 U385 ( .A(G472), .ZN(n504) );
  AND2_X1 U386 ( .A1(n610), .A2(n503), .ZN(n505) );
  XNOR2_X1 U387 ( .A(n393), .B(KEYINPUT5), .ZN(n392) );
  NAND2_X1 U388 ( .A1(n499), .A2(G210), .ZN(n393) );
  XNOR2_X1 U389 ( .A(n500), .B(n391), .ZN(n390) );
  XNOR2_X1 U390 ( .A(G137), .B(G113), .ZN(n500) );
  XNOR2_X1 U391 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n391) );
  INV_X1 U392 ( .A(n677), .ZN(n401) );
  INV_X1 U393 ( .A(n555), .ZN(n406) );
  INV_X1 U394 ( .A(KEYINPUT44), .ZN(n581) );
  AND2_X1 U395 ( .A1(n359), .A2(n412), .ZN(n411) );
  AND2_X1 U396 ( .A1(n547), .A2(KEYINPUT104), .ZN(n412) );
  INV_X1 U397 ( .A(KEYINPUT106), .ZN(n593) );
  NOR2_X1 U398 ( .A1(G953), .A2(G237), .ZN(n499) );
  XNOR2_X1 U399 ( .A(n433), .B(n432), .ZN(n725) );
  XOR2_X1 U400 ( .A(G134), .B(G131), .Z(n432) );
  XNOR2_X1 U401 ( .A(n457), .B(n427), .ZN(n433) );
  INV_X1 U402 ( .A(KEYINPUT4), .ZN(n427) );
  XOR2_X1 U403 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n424) );
  XNOR2_X1 U404 ( .A(n438), .B(G469), .ZN(n439) );
  XNOR2_X1 U405 ( .A(n725), .B(n394), .ZN(n502) );
  INV_X1 U406 ( .A(G146), .ZN(n394) );
  XOR2_X1 U407 ( .A(G104), .B(G107), .Z(n435) );
  NAND2_X1 U408 ( .A1(n383), .A2(n382), .ZN(n556) );
  NOR2_X1 U409 ( .A1(n507), .A2(n633), .ZN(n551) );
  INV_X1 U410 ( .A(KEYINPUT112), .ZN(n360) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n576) );
  INV_X1 U412 ( .A(KEYINPUT22), .ZN(n366) );
  XNOR2_X1 U413 ( .A(n493), .B(n416), .ZN(n494) );
  XNOR2_X1 U414 ( .A(n650), .B(KEYINPUT6), .ZN(n583) );
  XNOR2_X1 U415 ( .A(n613), .B(n354), .ZN(n369) );
  NAND2_X1 U416 ( .A1(n608), .A2(n609), .ZN(n613) );
  XNOR2_X1 U417 ( .A(KEYINPUT85), .B(G110), .ZN(n718) );
  INV_X1 U418 ( .A(KEYINPUT71), .ZN(n373) );
  XNOR2_X1 U419 ( .A(G146), .B(G125), .ZN(n447) );
  XNOR2_X1 U420 ( .A(n544), .B(n521), .ZN(n662) );
  OR2_X2 U421 ( .A1(n646), .A2(n562), .ZN(n652) );
  XOR2_X1 U422 ( .A(KEYINPUT89), .B(KEYINPUT20), .Z(n478) );
  INV_X1 U423 ( .A(G902), .ZN(n503) );
  XNOR2_X1 U424 ( .A(n347), .B(n502), .ZN(n610) );
  XNOR2_X1 U425 ( .A(n392), .B(n390), .ZN(n501) );
  NOR2_X1 U426 ( .A1(n644), .A2(n405), .ZN(n404) );
  INV_X1 U427 ( .A(n643), .ZN(n405) );
  XNOR2_X1 U428 ( .A(KEYINPUT10), .B(n447), .ZN(n486) );
  OR2_X1 U429 ( .A1(G237), .A2(G902), .ZN(n508) );
  NAND2_X1 U430 ( .A1(n534), .A2(n388), .ZN(n387) );
  INV_X1 U431 ( .A(n534), .ZN(n386) );
  INV_X1 U432 ( .A(n669), .ZN(n355) );
  AND2_X1 U433 ( .A1(n401), .A2(n559), .ZN(n400) );
  NAND2_X1 U434 ( .A1(n600), .A2(n599), .ZN(n608) );
  AND2_X1 U435 ( .A1(n607), .A2(G472), .ZN(n609) );
  XNOR2_X1 U436 ( .A(n582), .B(n581), .ZN(n596) );
  XNOR2_X1 U437 ( .A(KEYINPUT8), .B(KEYINPUT66), .ZN(n462) );
  XNOR2_X1 U438 ( .A(G128), .B(G110), .ZN(n484) );
  XNOR2_X1 U439 ( .A(n364), .B(G134), .ZN(n460) );
  XNOR2_X1 U440 ( .A(G143), .B(G122), .ZN(n449) );
  XOR2_X1 U441 ( .A(G131), .B(G140), .Z(n444) );
  XNOR2_X1 U442 ( .A(n361), .B(n430), .ZN(n690) );
  XNOR2_X1 U443 ( .A(n716), .B(n425), .ZN(n361) );
  NAND2_X1 U444 ( .A1(G234), .A2(G237), .ZN(n470) );
  NOR2_X1 U445 ( .A1(n531), .A2(n514), .ZN(n519) );
  XNOR2_X1 U446 ( .A(n375), .B(n513), .ZN(n514) );
  BUF_X1 U447 ( .A(n693), .Z(n704) );
  XNOR2_X1 U448 ( .A(n395), .B(n502), .ZN(n696) );
  XNOR2_X1 U449 ( .A(n434), .B(n350), .ZN(n396) );
  INV_X1 U450 ( .A(G953), .ZN(n687) );
  XNOR2_X1 U451 ( .A(n389), .B(n536), .ZN(n736) );
  NAND2_X1 U452 ( .A1(n556), .A2(n635), .ZN(n389) );
  NAND2_X1 U453 ( .A1(n379), .A2(n569), .ZN(n380) );
  XNOR2_X1 U454 ( .A(n554), .B(KEYINPUT36), .ZN(n379) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n734) );
  XNOR2_X1 U456 ( .A(KEYINPUT35), .B(KEYINPUT75), .ZN(n397) );
  BUF_X1 U457 ( .A(G116), .Z(n364) );
  INV_X1 U458 ( .A(KEYINPUT96), .ZN(n362) );
  NOR2_X1 U459 ( .A1(n646), .A2(n585), .ZN(n618) );
  AND2_X1 U460 ( .A1(n369), .A2(n368), .ZN(n617) );
  INV_X1 U461 ( .A(KEYINPUT56), .ZN(n371) );
  XNOR2_X1 U462 ( .A(n505), .B(n504), .ZN(n650) );
  XOR2_X1 U463 ( .A(n498), .B(n501), .Z(n347) );
  XOR2_X1 U464 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n348) );
  AND2_X1 U465 ( .A1(n518), .A2(n517), .ZN(n349) );
  XOR2_X1 U466 ( .A(n487), .B(n435), .Z(n350) );
  XOR2_X1 U467 ( .A(n431), .B(KEYINPUT86), .Z(n351) );
  AND2_X1 U468 ( .A1(n406), .A2(n402), .ZN(n352) );
  AND2_X1 U469 ( .A1(n386), .A2(n535), .ZN(n353) );
  INV_X1 U470 ( .A(n708), .ZN(n368) );
  XOR2_X1 U471 ( .A(KEYINPUT15), .B(G902), .Z(n597) );
  XOR2_X1 U472 ( .A(n612), .B(n611), .Z(n354) );
  INV_X1 U473 ( .A(n356), .ZN(n670) );
  OR2_X2 U474 ( .A1(n588), .A2(n583), .ZN(n356) );
  XNOR2_X1 U475 ( .A(n577), .B(n578), .ZN(n399) );
  NAND2_X1 U476 ( .A1(n662), .A2(n661), .ZN(n523) );
  NOR2_X1 U477 ( .A1(n540), .A2(n378), .ZN(n377) );
  NAND2_X1 U478 ( .A1(n560), .A2(n400), .ZN(n358) );
  XNOR2_X1 U479 ( .A(n358), .B(KEYINPUT0), .ZN(n561) );
  NAND2_X1 U480 ( .A1(n357), .A2(n352), .ZN(n600) );
  INV_X1 U481 ( .A(n712), .ZN(n357) );
  XNOR2_X2 U482 ( .A(n407), .B(KEYINPUT45), .ZN(n712) );
  NAND2_X1 U483 ( .A1(n408), .A2(n409), .ZN(n359) );
  XNOR2_X1 U484 ( .A(n551), .B(n360), .ZN(n552) );
  XNOR2_X1 U485 ( .A(n381), .B(KEYINPUT48), .ZN(n555) );
  XNOR2_X2 U486 ( .A(n363), .B(n362), .ZN(n620) );
  NAND2_X1 U487 ( .A1(n365), .A2(n589), .ZN(n363) );
  XNOR2_X1 U488 ( .A(n587), .B(KEYINPUT93), .ZN(n365) );
  NAND2_X1 U489 ( .A1(n406), .A2(n404), .ZN(n726) );
  NAND2_X1 U490 ( .A1(n399), .A2(n579), .ZN(n398) );
  XNOR2_X2 U491 ( .A(n370), .B(n351), .ZN(n520) );
  XNOR2_X1 U492 ( .A(n372), .B(n371), .ZN(G51) );
  NAND2_X1 U493 ( .A1(n692), .A2(n368), .ZN(n372) );
  NOR2_X2 U494 ( .A1(n570), .A2(n569), .ZN(n584) );
  NOR2_X2 U495 ( .A1(n589), .A2(n588), .ZN(n658) );
  INV_X1 U496 ( .A(n639), .ZN(n409) );
  XNOR2_X1 U497 ( .A(n592), .B(KEYINPUT98), .ZN(n639) );
  XNOR2_X1 U498 ( .A(n437), .B(n396), .ZN(n395) );
  XNOR2_X1 U499 ( .A(n374), .B(n373), .ZN(n549) );
  AND2_X1 U500 ( .A1(n548), .A2(n547), .ZN(n374) );
  NAND2_X1 U501 ( .A1(n414), .A2(n376), .ZN(n413) );
  NAND2_X1 U502 ( .A1(n410), .A2(n409), .ZN(n376) );
  NAND2_X1 U503 ( .A1(n377), .A2(n380), .ZN(n381) );
  NAND2_X1 U504 ( .A1(n550), .A2(n349), .ZN(n378) );
  INV_X1 U505 ( .A(n380), .ZN(n641) );
  NAND2_X1 U506 ( .A1(n385), .A2(n353), .ZN(n382) );
  AND2_X1 U507 ( .A1(n384), .A2(n387), .ZN(n383) );
  NAND2_X1 U508 ( .A1(n543), .A2(n388), .ZN(n384) );
  INV_X1 U509 ( .A(n543), .ZN(n385) );
  INV_X1 U510 ( .A(n535), .ZN(n388) );
  NOR2_X2 U511 ( .A1(n712), .A2(n726), .ZN(n645) );
  XNOR2_X2 U512 ( .A(n553), .B(KEYINPUT19), .ZN(n560) );
  NOR2_X2 U513 ( .A1(n595), .A2(n596), .ZN(n407) );
  INV_X1 U514 ( .A(n620), .ZN(n408) );
  NOR2_X1 U515 ( .A1(n620), .A2(KEYINPUT104), .ZN(n410) );
  NOR2_X1 U516 ( .A1(n618), .A2(n415), .ZN(n414) );
  XNOR2_X1 U517 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X1 U518 ( .A1(n727), .A2(G952), .ZN(n708) );
  XOR2_X1 U519 ( .A(KEYINPUT90), .B(KEYINPUT25), .Z(n416) );
  XOR2_X1 U520 ( .A(n695), .B(n694), .Z(n417) );
  INV_X1 U521 ( .A(n736), .ZN(n537) );
  XNOR2_X1 U522 ( .A(n539), .B(KEYINPUT46), .ZN(n540) );
  XNOR2_X1 U523 ( .A(G101), .B(G116), .ZN(n418) );
  XNOR2_X1 U524 ( .A(KEYINPUT38), .B(KEYINPUT72), .ZN(n521) );
  INV_X1 U525 ( .A(KEYINPUT62), .ZN(n611) );
  XNOR2_X1 U526 ( .A(n602), .B(n601), .ZN(n603) );
  INV_X1 U527 ( .A(KEYINPUT80), .ZN(n614) );
  XNOR2_X1 U528 ( .A(n696), .B(n417), .ZN(n697) );
  XNOR2_X1 U529 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U530 ( .A(n617), .B(n616), .ZN(G57) );
  INV_X1 U531 ( .A(n418), .ZN(n420) );
  XNOR2_X1 U532 ( .A(KEYINPUT3), .B(G119), .ZN(n419) );
  XNOR2_X1 U533 ( .A(n420), .B(n419), .ZN(n497) );
  XNOR2_X1 U534 ( .A(n497), .B(KEYINPUT16), .ZN(n422) );
  XOR2_X1 U535 ( .A(G113), .B(G104), .Z(n448) );
  XOR2_X1 U536 ( .A(G122), .B(G107), .Z(n456) );
  XOR2_X1 U537 ( .A(n448), .B(n456), .Z(n421) );
  XOR2_X2 U538 ( .A(KEYINPUT64), .B(G953), .Z(n727) );
  NAND2_X1 U539 ( .A1(G224), .A2(n727), .ZN(n423) );
  XNOR2_X1 U540 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U541 ( .A(KEYINPUT68), .B(n718), .ZN(n436) );
  INV_X1 U542 ( .A(n447), .ZN(n426) );
  XOR2_X1 U543 ( .A(n436), .B(n426), .Z(n429) );
  XNOR2_X1 U544 ( .A(n433), .B(KEYINPUT18), .ZN(n428) );
  XNOR2_X1 U545 ( .A(n429), .B(n428), .ZN(n430) );
  NAND2_X1 U546 ( .A1(G210), .A2(n508), .ZN(n431) );
  NAND2_X1 U547 ( .A1(G227), .A2(n727), .ZN(n434) );
  XOR2_X1 U548 ( .A(G101), .B(n436), .Z(n437) );
  INV_X1 U549 ( .A(KEYINPUT67), .ZN(n438) );
  XNOR2_X2 U550 ( .A(n440), .B(n439), .ZN(n531) );
  INV_X1 U551 ( .A(n653), .ZN(n569) );
  XNOR2_X1 U552 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n454) );
  XOR2_X1 U553 ( .A(KEYINPUT99), .B(KEYINPUT11), .Z(n442) );
  XNOR2_X1 U554 ( .A(KEYINPUT100), .B(KEYINPUT12), .ZN(n441) );
  XNOR2_X1 U555 ( .A(n442), .B(n441), .ZN(n446) );
  NAND2_X1 U556 ( .A1(G214), .A2(n499), .ZN(n443) );
  XNOR2_X1 U557 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U558 ( .A(n446), .B(n445), .ZN(n452) );
  XOR2_X1 U559 ( .A(n486), .B(n448), .Z(n450) );
  XNOR2_X1 U560 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U561 ( .A(n452), .B(n451), .ZN(n602) );
  NOR2_X1 U562 ( .A1(G902), .A2(n602), .ZN(n453) );
  XNOR2_X1 U563 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U564 ( .A(G475), .B(n455), .Z(n541) );
  INV_X1 U565 ( .A(n541), .ZN(n516) );
  XOR2_X1 U566 ( .A(KEYINPUT102), .B(KEYINPUT7), .Z(n459) );
  XNOR2_X1 U567 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U568 ( .A(n459), .B(n458), .ZN(n468) );
  XOR2_X1 U569 ( .A(KEYINPUT103), .B(KEYINPUT9), .Z(n461) );
  XNOR2_X1 U570 ( .A(n461), .B(n460), .ZN(n466) );
  NAND2_X1 U571 ( .A1(G234), .A2(n727), .ZN(n464) );
  XNOR2_X1 U572 ( .A(n462), .B(KEYINPUT79), .ZN(n463) );
  XNOR2_X1 U573 ( .A(n464), .B(n463), .ZN(n489) );
  NAND2_X1 U574 ( .A1(n489), .A2(G217), .ZN(n465) );
  XOR2_X1 U575 ( .A(n466), .B(n465), .Z(n467) );
  XNOR2_X1 U576 ( .A(n468), .B(n467), .ZN(n701) );
  NOR2_X1 U577 ( .A1(n701), .A2(G902), .ZN(n469) );
  XOR2_X1 U578 ( .A(n469), .B(G478), .Z(n542) );
  NOR2_X1 U579 ( .A1(n516), .A2(n542), .ZN(n635) );
  INV_X1 U580 ( .A(n635), .ZN(n633) );
  XOR2_X1 U581 ( .A(n470), .B(KEYINPUT14), .Z(n677) );
  OR2_X1 U582 ( .A1(n503), .A2(n677), .ZN(n471) );
  NOR2_X1 U583 ( .A1(n727), .A2(n471), .ZN(n472) );
  XNOR2_X1 U584 ( .A(n472), .B(KEYINPUT107), .ZN(n473) );
  NOR2_X1 U585 ( .A1(G900), .A2(n473), .ZN(n475) );
  NAND2_X1 U586 ( .A1(G952), .A2(n687), .ZN(n557) );
  NOR2_X1 U587 ( .A1(n677), .A2(n557), .ZN(n474) );
  NOR2_X1 U588 ( .A1(n475), .A2(n474), .ZN(n530) );
  INV_X1 U589 ( .A(n597), .ZN(n476) );
  NAND2_X1 U590 ( .A1(G234), .A2(n476), .ZN(n477) );
  XNOR2_X1 U591 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U592 ( .A(KEYINPUT88), .B(n479), .ZN(n492) );
  NAND2_X1 U593 ( .A1(G221), .A2(n492), .ZN(n480) );
  XNOR2_X1 U594 ( .A(KEYINPUT21), .B(n480), .ZN(n647) );
  NOR2_X1 U595 ( .A1(n530), .A2(n647), .ZN(n496) );
  XNOR2_X1 U596 ( .A(G119), .B(KEYINPUT87), .ZN(n481) );
  XNOR2_X1 U597 ( .A(n348), .B(n481), .ZN(n483) );
  INV_X1 U598 ( .A(KEYINPUT74), .ZN(n482) );
  XNOR2_X1 U599 ( .A(n483), .B(n482), .ZN(n485) );
  XNOR2_X1 U600 ( .A(n485), .B(n484), .ZN(n488) );
  XOR2_X1 U601 ( .A(n487), .B(n486), .Z(n723) );
  XOR2_X1 U602 ( .A(n723), .B(n488), .Z(n491) );
  NAND2_X1 U603 ( .A1(G221), .A2(n489), .ZN(n490) );
  XNOR2_X1 U604 ( .A(n491), .B(n490), .ZN(n703) );
  NOR2_X1 U605 ( .A1(G902), .A2(n703), .ZN(n495) );
  NAND2_X1 U606 ( .A1(G217), .A2(n492), .ZN(n493) );
  XNOR2_X2 U607 ( .A(n495), .B(n494), .ZN(n646) );
  NAND2_X1 U608 ( .A1(n496), .A2(n646), .ZN(n512) );
  BUF_X1 U609 ( .A(n497), .Z(n498) );
  NOR2_X1 U610 ( .A1(n512), .A2(n583), .ZN(n506) );
  XOR2_X1 U611 ( .A(KEYINPUT108), .B(n506), .Z(n507) );
  NAND2_X1 U612 ( .A1(G214), .A2(n508), .ZN(n661) );
  NAND2_X1 U613 ( .A1(n551), .A2(n661), .ZN(n509) );
  NOR2_X1 U614 ( .A1(n569), .A2(n509), .ZN(n510) );
  XNOR2_X1 U615 ( .A(n510), .B(KEYINPUT43), .ZN(n511) );
  NOR2_X1 U616 ( .A1(n520), .A2(n511), .ZN(n644) );
  XOR2_X1 U617 ( .A(KEYINPUT110), .B(KEYINPUT28), .Z(n513) );
  NAND2_X1 U618 ( .A1(n519), .A2(n560), .ZN(n632) );
  NAND2_X1 U619 ( .A1(n632), .A2(KEYINPUT47), .ZN(n515) );
  XNOR2_X1 U620 ( .A(n515), .B(KEYINPUT78), .ZN(n518) );
  NAND2_X1 U621 ( .A1(n542), .A2(n516), .ZN(n627) );
  NAND2_X1 U622 ( .A1(n633), .A2(n627), .ZN(n547) );
  INV_X1 U623 ( .A(n547), .ZN(n666) );
  NAND2_X1 U624 ( .A1(n666), .A2(KEYINPUT47), .ZN(n517) );
  INV_X1 U625 ( .A(n519), .ZN(n526) );
  INV_X1 U626 ( .A(n520), .ZN(n544) );
  INV_X1 U627 ( .A(KEYINPUT111), .ZN(n522) );
  XNOR2_X1 U628 ( .A(n523), .B(n522), .ZN(n665) );
  NOR2_X1 U629 ( .A1(n541), .A2(n542), .ZN(n524) );
  XNOR2_X1 U630 ( .A(n524), .B(KEYINPUT105), .ZN(n664) );
  NOR2_X1 U631 ( .A1(n665), .A2(n664), .ZN(n525) );
  XNOR2_X1 U632 ( .A(n525), .B(KEYINPUT41), .ZN(n681) );
  NOR2_X1 U633 ( .A1(n526), .A2(n681), .ZN(n527) );
  XNOR2_X1 U634 ( .A(n527), .B(KEYINPUT42), .ZN(n737) );
  INV_X1 U635 ( .A(n737), .ZN(n538) );
  NAND2_X1 U636 ( .A1(n650), .A2(n661), .ZN(n528) );
  XNOR2_X1 U637 ( .A(KEYINPUT30), .B(n528), .ZN(n529) );
  NOR2_X1 U638 ( .A1(n530), .A2(n529), .ZN(n533) );
  XOR2_X1 U639 ( .A(n647), .B(KEYINPUT91), .Z(n562) );
  NOR2_X2 U640 ( .A1(n531), .A2(n652), .ZN(n532) );
  XNOR2_X1 U641 ( .A(KEYINPUT92), .B(n532), .ZN(n586) );
  NAND2_X1 U642 ( .A1(n533), .A2(n586), .ZN(n543) );
  INV_X1 U643 ( .A(n662), .ZN(n534) );
  XNOR2_X1 U644 ( .A(KEYINPUT69), .B(KEYINPUT39), .ZN(n535) );
  INV_X1 U645 ( .A(KEYINPUT40), .ZN(n536) );
  NAND2_X1 U646 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U647 ( .A1(n542), .A2(n541), .ZN(n573) );
  NOR2_X1 U648 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U649 ( .A(n545), .B(KEYINPUT109), .ZN(n546) );
  NOR2_X1 U650 ( .A1(n573), .A2(n546), .ZN(n631) );
  NOR2_X1 U651 ( .A1(KEYINPUT47), .A2(n632), .ZN(n548) );
  NOR2_X1 U652 ( .A1(n631), .A2(n549), .ZN(n550) );
  NOR2_X1 U653 ( .A1(n553), .A2(n552), .ZN(n554) );
  INV_X1 U654 ( .A(n627), .ZN(n638) );
  NAND2_X1 U655 ( .A1(n556), .A2(n638), .ZN(n643) );
  INV_X1 U656 ( .A(n664), .ZN(n564) );
  NOR2_X1 U657 ( .A1(G898), .A2(n687), .ZN(n720) );
  NAND2_X1 U658 ( .A1(n720), .A2(G902), .ZN(n558) );
  NAND2_X1 U659 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U660 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U661 ( .A1(n646), .A2(n583), .ZN(n565) );
  NOR2_X1 U662 ( .A1(n653), .A2(n565), .ZN(n566) );
  XNOR2_X1 U663 ( .A(n566), .B(KEYINPUT77), .ZN(n567) );
  NOR2_X1 U664 ( .A1(n570), .A2(n567), .ZN(n568) );
  XNOR2_X1 U665 ( .A(KEYINPUT32), .B(n568), .ZN(n735) );
  AND2_X1 U666 ( .A1(n646), .A2(n589), .ZN(n571) );
  NAND2_X1 U667 ( .A1(n571), .A2(n584), .ZN(n625) );
  INV_X1 U668 ( .A(n625), .ZN(n572) );
  NOR2_X1 U669 ( .A1(n735), .A2(n572), .ZN(n580) );
  XOR2_X1 U670 ( .A(n573), .B(KEYINPUT76), .Z(n579) );
  XOR2_X1 U671 ( .A(KEYINPUT70), .B(KEYINPUT34), .Z(n578) );
  NOR2_X1 U672 ( .A1(n652), .A2(n653), .ZN(n574) );
  XNOR2_X1 U673 ( .A(n574), .B(KEYINPUT73), .ZN(n588) );
  XNOR2_X1 U674 ( .A(KEYINPUT81), .B(KEYINPUT33), .ZN(n669) );
  INV_X1 U675 ( .A(n561), .ZN(n575) );
  NAND2_X1 U676 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U677 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U678 ( .A1(n586), .A2(n575), .ZN(n587) );
  XOR2_X1 U679 ( .A(KEYINPUT31), .B(KEYINPUT97), .Z(n591) );
  NAND2_X1 U680 ( .A1(n658), .A2(n575), .ZN(n590) );
  XNOR2_X1 U681 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U682 ( .A(n594), .B(n593), .ZN(n595) );
  NAND2_X1 U683 ( .A1(n597), .A2(KEYINPUT2), .ZN(n598) );
  XOR2_X1 U684 ( .A(KEYINPUT65), .B(n598), .Z(n599) );
  NAND2_X1 U685 ( .A1(KEYINPUT2), .A2(n645), .ZN(n607) );
  AND2_X2 U686 ( .A1(n608), .A2(n607), .ZN(n693) );
  NAND2_X1 U687 ( .A1(n693), .A2(G475), .ZN(n604) );
  XOR2_X1 U688 ( .A(KEYINPUT59), .B(KEYINPUT122), .Z(n601) );
  XNOR2_X1 U689 ( .A(n604), .B(n603), .ZN(n605) );
  NOR2_X2 U690 ( .A1(n605), .A2(n708), .ZN(n606) );
  XNOR2_X1 U691 ( .A(n606), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U692 ( .A(n610), .B(KEYINPUT83), .Z(n612) );
  XNOR2_X1 U693 ( .A(KEYINPUT63), .B(KEYINPUT84), .ZN(n615) );
  XOR2_X1 U694 ( .A(n618), .B(G101), .Z(G3) );
  NAND2_X1 U695 ( .A1(n620), .A2(n635), .ZN(n619) );
  XNOR2_X1 U696 ( .A(n619), .B(G104), .ZN(G6) );
  XOR2_X1 U697 ( .A(KEYINPUT113), .B(KEYINPUT27), .Z(n622) );
  NAND2_X1 U698 ( .A1(n638), .A2(n620), .ZN(n621) );
  XNOR2_X1 U699 ( .A(n622), .B(n621), .ZN(n624) );
  XOR2_X1 U700 ( .A(G107), .B(KEYINPUT26), .Z(n623) );
  XNOR2_X1 U701 ( .A(n624), .B(n623), .ZN(G9) );
  XNOR2_X1 U702 ( .A(G110), .B(KEYINPUT114), .ZN(n626) );
  XNOR2_X1 U703 ( .A(n626), .B(n625), .ZN(G12) );
  NOR2_X1 U704 ( .A1(n627), .A2(n632), .ZN(n629) );
  XNOR2_X1 U705 ( .A(KEYINPUT29), .B(KEYINPUT115), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n629), .B(n628), .ZN(n630) );
  XOR2_X1 U707 ( .A(G128), .B(n630), .Z(G30) );
  XOR2_X1 U708 ( .A(G143), .B(n631), .Z(G45) );
  NOR2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U710 ( .A(G146), .B(n634), .Z(G48) );
  NAND2_X1 U711 ( .A1(n639), .A2(n635), .ZN(n636) );
  XNOR2_X1 U712 ( .A(n636), .B(KEYINPUT116), .ZN(n637) );
  XNOR2_X1 U713 ( .A(G113), .B(n637), .ZN(G15) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n640), .B(n364), .ZN(G18) );
  XNOR2_X1 U716 ( .A(G125), .B(n641), .ZN(n642) );
  XNOR2_X1 U717 ( .A(n642), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U718 ( .A(G134), .B(n643), .ZN(G36) );
  XOR2_X1 U719 ( .A(G140), .B(n644), .Z(G42) );
  XNOR2_X1 U720 ( .A(KEYINPUT2), .B(n645), .ZN(n680) );
  NAND2_X1 U721 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U722 ( .A(KEYINPUT49), .B(n648), .ZN(n649) );
  NOR2_X1 U723 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U724 ( .A(KEYINPUT117), .B(n651), .ZN(n656) );
  NAND2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U726 ( .A(KEYINPUT50), .B(n654), .Z(n655) );
  NOR2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U729 ( .A(KEYINPUT51), .B(n659), .Z(n660) );
  NOR2_X1 U730 ( .A1(n681), .A2(n660), .ZN(n673) );
  NOR2_X1 U731 ( .A1(n386), .A2(n661), .ZN(n663) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n668) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n671) );
  XOR2_X1 U735 ( .A(n670), .B(n669), .Z(n682) );
  NOR2_X1 U736 ( .A1(n671), .A2(n682), .ZN(n672) );
  NOR2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U738 ( .A(n674), .B(KEYINPUT52), .ZN(n675) );
  XNOR2_X1 U739 ( .A(KEYINPUT118), .B(n675), .ZN(n676) );
  NOR2_X1 U740 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U741 ( .A1(n678), .A2(G952), .ZN(n679) );
  NAND2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n685) );
  NOR2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U744 ( .A(KEYINPUT119), .B(n683), .Z(n684) );
  NOR2_X1 U745 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U746 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U747 ( .A(KEYINPUT53), .B(n688), .Z(G75) );
  NAND2_X1 U748 ( .A1(n693), .A2(G210), .ZN(n691) );
  XOR2_X1 U749 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n689) );
  XNOR2_X1 U750 ( .A(n691), .B(n346), .ZN(n692) );
  NAND2_X1 U751 ( .A1(n704), .A2(G469), .ZN(n698) );
  XOR2_X1 U752 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n695) );
  XNOR2_X1 U753 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n694) );
  NOR2_X1 U754 ( .A1(n708), .A2(n699), .ZN(G54) );
  NAND2_X1 U755 ( .A1(G478), .A2(n704), .ZN(n700) );
  XNOR2_X1 U756 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U757 ( .A1(n708), .A2(n702), .ZN(G63) );
  XOR2_X1 U758 ( .A(n703), .B(KEYINPUT123), .Z(n706) );
  NAND2_X1 U759 ( .A1(n704), .A2(G217), .ZN(n705) );
  XNOR2_X1 U760 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U761 ( .A1(n708), .A2(n707), .ZN(G66) );
  NAND2_X1 U762 ( .A1(G224), .A2(G953), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n709), .B(KEYINPUT124), .ZN(n710) );
  XNOR2_X1 U764 ( .A(KEYINPUT61), .B(n710), .ZN(n711) );
  AND2_X1 U765 ( .A1(n711), .A2(G898), .ZN(n714) );
  NOR2_X1 U766 ( .A1(G953), .A2(n712), .ZN(n713) );
  NOR2_X1 U767 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n715), .B(KEYINPUT125), .ZN(n722) );
  XOR2_X1 U769 ( .A(n716), .B(KEYINPUT126), .Z(n717) );
  XNOR2_X1 U770 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n722), .B(n721), .ZN(G69) );
  XOR2_X1 U773 ( .A(n723), .B(KEYINPUT127), .Z(n724) );
  XNOR2_X1 U774 ( .A(n725), .B(n724), .ZN(n729) );
  XNOR2_X1 U775 ( .A(n726), .B(n729), .ZN(n728) );
  NAND2_X1 U776 ( .A1(n728), .A2(n727), .ZN(n733) );
  XNOR2_X1 U777 ( .A(G227), .B(n729), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n730), .A2(G900), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n731), .A2(G953), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n733), .A2(n732), .ZN(G72) );
  XNOR2_X1 U781 ( .A(n734), .B(G122), .ZN(G24) );
  XOR2_X1 U782 ( .A(G119), .B(n735), .Z(G21) );
  XOR2_X1 U783 ( .A(n736), .B(G131), .Z(G33) );
  XOR2_X1 U784 ( .A(n737), .B(G137), .Z(G39) );
endmodule

