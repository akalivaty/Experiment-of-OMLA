//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n450, new_n451, new_n453,
    new_n455, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g024(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n450));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(G223));
  INV_X1    g027(.A(new_n451), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n453), .A2(G567), .ZN(G234));
  NAND2_X1  g029(.A1(new_n453), .A2(G2106), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT69), .ZN(G217));
  NOR4_X1   g031(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT2), .ZN(new_n458));
  NOR4_X1   g033(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(G261));
  INV_X1    g035(.A(G261), .ZN(G325));
  INV_X1    g036(.A(G2106), .ZN(new_n462));
  INV_X1    g037(.A(G567), .ZN(new_n463));
  OAI22_X1  g038(.A1(new_n458), .A2(new_n462), .B1(new_n463), .B2(new_n459), .ZN(new_n464));
  XOR2_X1   g039(.A(new_n464), .B(KEYINPUT70), .Z(G319));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(KEYINPUT71), .A3(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT71), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n474), .B1(KEYINPUT72), .B2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT3), .B1(new_n476), .B2(KEYINPUT71), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n473), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(G137), .A3(new_n466), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n476), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G101), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT73), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n479), .A2(KEYINPUT73), .A3(new_n481), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n470), .B1(new_n484), .B2(new_n485), .ZN(G160));
  NAND2_X1  g061(.A1(new_n478), .A2(new_n466), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G112), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n471), .A2(KEYINPUT71), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n474), .A2(G2104), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n493), .A2(KEYINPUT3), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n466), .B1(new_n495), .B2(new_n473), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(new_n496), .B2(G124), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n489), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G2105), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n502), .B1(new_n496), .B2(G126), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n466), .A2(G138), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n467), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n504), .B1(new_n478), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(KEYINPUT74), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(new_n495), .B2(new_n473), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  NOR3_X1   g086(.A1(new_n510), .A2(new_n511), .A3(new_n504), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n503), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT75), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT75), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n515), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  XOR2_X1   g096(.A(KEYINPUT76), .B(G88), .Z(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n515), .A2(G62), .ZN(new_n524));
  INV_X1    g099(.A(G75), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT77), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OR3_X1    g102(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT77), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT6), .B(G651), .Z(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n526), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n529), .A2(G651), .B1(new_n531), .B2(G50), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n523), .A2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND3_X1  g109(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT78), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT79), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n530), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n516), .A2(KEYINPUT79), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n542), .A2(G543), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G51), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n521), .A2(G89), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n540), .A2(new_n546), .A3(new_n547), .ZN(G168));
  NAND2_X1  g123(.A1(new_n521), .A2(G90), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(G52), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G651), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  NAND2_X1  g130(.A1(new_n521), .A2(G81), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n545), .A2(G43), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(new_n552), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g138(.A(KEYINPUT80), .B(KEYINPUT8), .Z(new_n564));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n568));
  INV_X1    g143(.A(G78), .ZN(new_n569));
  INV_X1    g144(.A(new_n515), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI221_X1 g146(.A(new_n568), .B1(new_n569), .B2(new_n526), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n570), .A2(new_n571), .B1(new_n569), .B2(new_n526), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT81), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n573), .A2(new_n575), .B1(G91), .B2(new_n521), .ZN(new_n576));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OR3_X1    g152(.A1(new_n544), .A2(KEYINPUT9), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT9), .B1(new_n544), .B2(new_n577), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G299));
  NAND3_X1  g156(.A1(new_n540), .A2(new_n546), .A3(new_n547), .ZN(G286));
  NAND2_X1  g157(.A1(new_n521), .A2(G87), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT82), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n515), .A2(G74), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n545), .A2(G49), .B1(G651), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(G288));
  AOI22_X1  g163(.A1(new_n521), .A2(G86), .B1(G48), .B2(new_n531), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT84), .Z(new_n591));
  NAND2_X1  g166(.A1(new_n515), .A2(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(KEYINPUT83), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n592), .A2(KEYINPUT83), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT85), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g172(.A(KEYINPUT85), .B(G651), .C1(new_n593), .C2(new_n594), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n589), .B1(new_n597), .B2(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n518), .A2(new_n520), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  INV_X1    g177(.A(G47), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n601), .A2(new_n602), .B1(new_n544), .B2(new_n603), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n604), .A2(KEYINPUT86), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n604), .A2(KEYINPUT86), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n605), .A2(new_n606), .B1(new_n552), .B2(new_n607), .ZN(G290));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NOR2_X1   g184(.A1(G301), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G54), .ZN(new_n611));
  XOR2_X1   g186(.A(KEYINPUT89), .B(G66), .Z(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(new_n515), .B1(G79), .B2(G543), .ZN(new_n613));
  OAI22_X1  g188(.A1(new_n544), .A2(new_n611), .B1(new_n552), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n521), .A2(G92), .ZN(new_n615));
  XOR2_X1   g190(.A(KEYINPUT87), .B(KEYINPUT10), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT88), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n614), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G92), .ZN(new_n619));
  OR3_X1    g194(.A1(new_n601), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT90), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n610), .B1(new_n622), .B2(new_n609), .ZN(G284));
  AOI21_X1  g198(.A(new_n610), .B1(new_n622), .B2(new_n609), .ZN(G321));
  NAND2_X1  g199(.A1(G299), .A2(new_n609), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n609), .B2(G168), .ZN(G297));
  OAI21_X1  g201(.A(new_n625), .B1(new_n609), .B2(G168), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n622), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n622), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n467), .A2(new_n480), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT12), .Z(new_n635));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  OAI22_X1  g211(.A1(new_n635), .A2(KEYINPUT13), .B1(KEYINPUT91), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(KEYINPUT13), .B2(new_n635), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(KEYINPUT91), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n496), .A2(G123), .ZN(new_n641));
  INV_X1    g216(.A(G135), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n466), .A2(G111), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  OAI221_X1 g219(.A(new_n641), .B1(new_n487), .B2(new_n642), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n640), .A2(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT92), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n657), .A2(new_n660), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(G401));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  NOR2_X1   g239(.A1(G2072), .A2(G2078), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n444), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n664), .B1(new_n667), .B2(KEYINPUT93), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(KEYINPUT93), .B2(new_n667), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n666), .B(KEYINPUT17), .ZN(new_n672));
  INV_X1    g247(.A(new_n664), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n669), .B(new_n671), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n671), .A2(new_n666), .A3(new_n673), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT18), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n672), .A2(new_n673), .A3(new_n670), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2096), .B(G2100), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1971), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(new_n686), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT20), .Z(new_n690));
  AOI211_X1 g265(.A(new_n688), .B(new_n690), .C1(new_n683), .C2(new_n687), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n698), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(G1971), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(G23), .ZN(new_n702));
  INV_X1    g277(.A(G288), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n698), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT33), .B(G1976), .Z(new_n705));
  OAI21_X1  g280(.A(new_n701), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n704), .B2(new_n705), .ZN(new_n707));
  MUX2_X1   g282(.A(G6), .B(G305), .S(G16), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT95), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT32), .B(G1981), .Z(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n707), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(KEYINPUT34), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(KEYINPUT34), .ZN(new_n715));
  MUX2_X1   g290(.A(G24), .B(G290), .S(G16), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1986), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n718), .A2(G25), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n496), .A2(G119), .ZN(new_n720));
  OR2_X1    g295(.A1(G95), .A2(G2105), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n721), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n722));
  INV_X1    g297(.A(G131), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n720), .B(new_n722), .C1(new_n723), .C2(new_n487), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n719), .B1(new_n724), .B2(G29), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT94), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT96), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n725), .A2(new_n727), .B1(new_n728), .B2(KEYINPUT36), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n725), .B2(new_n727), .ZN(new_n730));
  OR4_X1    g305(.A1(new_n714), .A2(new_n715), .A3(new_n717), .A4(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n728), .A2(KEYINPUT36), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  INV_X1    g309(.A(G34), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n735), .A2(KEYINPUT24), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(KEYINPUT24), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n718), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G160), .B2(new_n718), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G2084), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n488), .A2(G141), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n496), .A2(G129), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT26), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n745), .A2(new_n746), .B1(G105), .B2(new_n480), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n741), .A2(new_n742), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(new_n718), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n718), .B2(G32), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT27), .B(G1996), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT31), .B(G11), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT30), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n755), .A2(G28), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n718), .B1(new_n755), .B2(G28), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n754), .B1(new_n756), .B2(new_n757), .C1(new_n645), .C2(new_n718), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n718), .A2(G33), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT25), .Z(new_n761));
  AOI22_X1  g336(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  INV_X1    g337(.A(G139), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n761), .B1(new_n762), .B2(new_n466), .C1(new_n487), .C2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n759), .B1(new_n764), .B2(G29), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n758), .B1(new_n766), .B2(G2072), .ZN(new_n767));
  NOR2_X1   g342(.A1(G16), .A2(G19), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n561), .B2(G16), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G1341), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n751), .A2(new_n752), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n753), .A2(new_n767), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n718), .A2(G26), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT97), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT28), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n496), .A2(G128), .ZN(new_n776));
  INV_X1    g351(.A(G140), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n466), .A2(G116), .ZN(new_n778));
  OAI21_X1  g353(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n779));
  OAI221_X1 g354(.A(new_n776), .B1(new_n487), .B2(new_n777), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n775), .B1(new_n780), .B2(G29), .ZN(new_n781));
  INV_X1    g356(.A(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n765), .A2(new_n442), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT98), .Z(new_n785));
  OR4_X1    g360(.A1(new_n740), .A2(new_n772), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n698), .A2(G4), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n622), .B2(new_n698), .ZN(new_n788));
  INV_X1    g363(.A(G1348), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n718), .A2(G35), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G162), .B2(new_n718), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT29), .ZN(new_n793));
  INV_X1    g368(.A(G2090), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n698), .A2(G20), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT23), .Z(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G299), .B2(G16), .ZN(new_n798));
  INV_X1    g373(.A(G1956), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(G27), .A2(G29), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G164), .B2(G29), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n800), .B1(G2078), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n790), .A2(new_n795), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n698), .A2(G5), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G171), .B2(new_n698), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT99), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G1961), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n769), .A2(G1341), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n698), .A2(G21), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G168), .B2(new_n698), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n809), .B1(G1966), .B2(new_n811), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n808), .B(new_n812), .C1(G1966), .C2(new_n811), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n807), .A2(G1961), .B1(G2078), .B2(new_n802), .ZN(new_n814));
  NOR4_X1   g389(.A1(new_n786), .A2(new_n804), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n733), .A2(new_n734), .A3(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  NAND2_X1  g392(.A1(new_n622), .A2(G559), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT38), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n521), .A2(G93), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n545), .A2(G55), .ZN(new_n821));
  NAND2_X1  g396(.A1(G80), .A2(G543), .ZN(new_n822));
  INV_X1    g397(.A(G67), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n570), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(KEYINPUT100), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(KEYINPUT100), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G651), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n820), .B(new_n821), .C1(new_n825), .C2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n560), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n819), .B(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n832), .A2(new_n833), .A3(G860), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n828), .A2(G860), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT101), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  OR2_X1    g412(.A1(new_n834), .A2(new_n837), .ZN(G145));
  XNOR2_X1  g413(.A(new_n780), .B(KEYINPUT103), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n764), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n724), .B(KEYINPUT104), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n635), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n840), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n513), .B(new_n748), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n496), .A2(G130), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n466), .A2(G118), .ZN(new_n846));
  OAI21_X1  g421(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G142), .B2(new_n488), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n844), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n843), .B(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n645), .B(new_n498), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT102), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G160), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT105), .ZN(new_n856));
  INV_X1    g431(.A(G37), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n856), .B(new_n857), .C1(new_n854), .C2(new_n851), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g434(.A1(new_n828), .A2(new_n609), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n630), .B(new_n829), .ZN(new_n861));
  XNOR2_X1  g436(.A(G299), .B(new_n621), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(G299), .B(new_n621), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT41), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT41), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n863), .B1(new_n861), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT42), .ZN(new_n870));
  XNOR2_X1  g445(.A(G288), .B(G290), .ZN(new_n871));
  XNOR2_X1  g446(.A(G305), .B(G303), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n870), .B(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n860), .B1(new_n875), .B2(new_n609), .ZN(G295));
  OAI21_X1  g451(.A(new_n860), .B1(new_n875), .B2(new_n609), .ZN(G331));
  INV_X1    g452(.A(KEYINPUT110), .ZN(new_n878));
  XNOR2_X1  g453(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(G168), .A2(G171), .ZN(new_n881));
  NOR2_X1   g456(.A1(G286), .A2(G301), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n830), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n829), .B1(new_n881), .B2(new_n882), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(new_n862), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(KEYINPUT107), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT107), .B1(new_n883), .B2(new_n830), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n887), .B1(new_n891), .B2(new_n868), .ZN(new_n892));
  AOI21_X1  g467(.A(G37), .B1(new_n892), .B2(new_n873), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n888), .A2(new_n864), .A3(new_n890), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n868), .A2(new_n886), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n873), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n897), .A2(KEYINPUT108), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n899));
  AOI211_X1 g474(.A(new_n899), .B(new_n873), .C1(new_n895), .C2(new_n896), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n893), .B(new_n894), .C1(new_n898), .C2(new_n900), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n892), .A2(new_n873), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n893), .ZN(new_n903));
  AOI22_X1  g478(.A1(new_n901), .A2(KEYINPUT109), .B1(KEYINPUT43), .B2(new_n903), .ZN(new_n904));
  AOI211_X1 g479(.A(new_n862), .B(new_n889), .C1(new_n886), .C2(KEYINPUT107), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n886), .A2(new_n867), .A3(new_n865), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n874), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n899), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n897), .A2(KEYINPUT108), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n910), .A2(new_n911), .A3(new_n894), .A4(new_n893), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n880), .B1(new_n904), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n902), .A2(new_n893), .A3(new_n894), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT44), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n893), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(KEYINPUT43), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n878), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n901), .A2(KEYINPUT109), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n903), .A2(KEYINPUT43), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n912), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n879), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(KEYINPUT44), .A3(new_n914), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(KEYINPUT110), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n918), .A2(new_n925), .ZN(G397));
  INV_X1    g501(.A(G1384), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n513), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n470), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n479), .A2(KEYINPUT73), .A3(new_n481), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT73), .B1(new_n479), .B2(new_n481), .ZN(new_n933));
  OAI211_X1 g508(.A(G40), .B(new_n931), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G1996), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT111), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n938), .A2(new_n748), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n935), .B(KEYINPUT112), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n780), .B(new_n782), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n936), .B2(new_n749), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n726), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n724), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n939), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  NOR4_X1   g522(.A1(G290), .A2(new_n930), .A3(G1986), .A4(new_n934), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT48), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n941), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n940), .B1(new_n748), .B2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n938), .A2(KEYINPUT46), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n938), .A2(KEYINPUT46), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT47), .Z(new_n956));
  NAND2_X1  g531(.A1(new_n939), .A2(new_n943), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n957), .A2(new_n724), .A3(new_n944), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n780), .A2(G2067), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI211_X1 g535(.A(new_n950), .B(new_n956), .C1(new_n940), .C2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1976), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT52), .B1(G288), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n928), .A2(new_n934), .ZN(new_n964));
  INV_X1    g539(.A(G8), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n963), .B(new_n966), .C1(new_n962), .C2(G288), .ZN(new_n967));
  INV_X1    g542(.A(new_n964), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n968), .B(G8), .C1(G288), .C2(new_n962), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT52), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n589), .A2(new_n595), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(G1981), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(G305), .B2(G1981), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT49), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n972), .B(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(new_n966), .A3(new_n976), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n967), .A2(new_n970), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n928), .A2(KEYINPUT50), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n511), .B1(new_n510), .B2(new_n504), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n478), .A2(new_n506), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(KEYINPUT74), .A3(KEYINPUT4), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n980), .A2(new_n982), .A3(new_n507), .ZN(new_n983));
  AOI21_X1  g558(.A(G1384), .B1(new_n983), .B2(new_n503), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n934), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n979), .A2(new_n794), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n927), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n987), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT113), .B1(new_n984), .B2(KEYINPUT45), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n928), .A2(new_n992), .A3(new_n929), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n990), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n988), .B1(new_n994), .B2(G1971), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(G8), .ZN(new_n996));
  NAND2_X1  g571(.A1(G303), .A2(G8), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n997), .B(KEYINPUT55), .Z(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n978), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n993), .A2(new_n991), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n934), .B1(new_n984), .B2(KEYINPUT45), .ZN(new_n1003));
  AOI21_X1  g578(.A(G1971), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n988), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT114), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n988), .B(new_n1007), .C1(new_n994), .C2(G1971), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1006), .A2(G8), .A3(new_n998), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n965), .B1(new_n995), .B2(KEYINPUT114), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1012), .A2(KEYINPUT115), .A3(new_n998), .A4(new_n1008), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1001), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1966), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n984), .A2(KEYINPUT45), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT117), .B(new_n1015), .C1(new_n990), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G2084), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n979), .A2(new_n1018), .A3(new_n986), .A4(new_n987), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1003), .A2(new_n930), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT117), .B1(new_n1021), .B2(new_n1015), .ZN(new_n1022));
  OAI21_X1  g597(.A(G286), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1015), .B1(new_n990), .B2(new_n1016), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1026), .A2(G168), .A3(new_n1019), .A4(new_n1017), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1023), .A2(G8), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT51), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(new_n1030), .A3(G8), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT53), .B1(new_n994), .B2(new_n443), .ZN(new_n1033));
  INV_X1    g608(.A(G1961), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n987), .B1(new_n985), .B2(new_n984), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n928), .A2(KEYINPUT50), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(G2078), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1003), .A2(new_n930), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1033), .A2(G171), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n992), .B1(new_n928), .B2(new_n929), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n984), .A2(KEYINPUT113), .A3(KEYINPUT45), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n443), .B(new_n1003), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n1038), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n990), .A2(new_n1016), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n979), .A2(new_n987), .A3(new_n986), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1047), .A2(new_n1039), .B1(new_n1048), .B2(new_n1034), .ZN(new_n1049));
  AOI21_X1  g624(.A(G301), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT54), .B1(new_n1042), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(G171), .B1(new_n1033), .B2(new_n1041), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1046), .A2(new_n1049), .A3(G301), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1032), .A2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT56), .B(G2072), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1003), .B(new_n1058), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n799), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT57), .ZN(new_n1063));
  XOR2_X1   g638(.A(new_n1063), .B(KEYINPUT121), .Z(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1062), .A2(KEYINPUT57), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1065), .B1(G299), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1066), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n576), .A2(new_n580), .A3(new_n1068), .A4(new_n1064), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1061), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1059), .A2(new_n1070), .A3(new_n1060), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1059), .A2(new_n1070), .A3(KEYINPUT124), .A4(new_n1060), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1076), .A2(KEYINPUT61), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1074), .A2(KEYINPUT122), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1059), .A2(new_n1070), .A3(new_n1080), .A4(new_n1060), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT61), .B1(new_n1061), .B2(new_n1071), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1078), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n936), .B(new_n1003), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT58), .B(G1341), .Z(new_n1088));
  NAND2_X1  g663(.A1(new_n968), .A2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1086), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1087), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n561), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT59), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1094), .B(new_n561), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT126), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT60), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n928), .A2(G2067), .A3(new_n934), .ZN(new_n1099));
  AOI211_X1 g674(.A(new_n1098), .B(new_n1099), .C1(new_n1048), .C2(new_n789), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1097), .B1(new_n1100), .B2(new_n621), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(new_n1102), .A3(new_n621), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1048), .A2(new_n789), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1099), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1104), .A2(KEYINPUT60), .A3(new_n621), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT125), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1108));
  OAI211_X1 g683(.A(KEYINPUT60), .B(new_n1105), .C1(new_n1108), .C2(G1348), .ZN(new_n1109));
  INV_X1    g684(.A(new_n621), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(KEYINPUT126), .A3(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1101), .A2(new_n1103), .A3(new_n1107), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1099), .B1(new_n1048), .B2(new_n789), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1113), .A2(KEYINPUT60), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1085), .A2(new_n1096), .A3(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1072), .B1(new_n621), .B2(new_n1113), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n1082), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1057), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1029), .A2(new_n1120), .A3(new_n1031), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1121), .A2(new_n1122), .A3(new_n1052), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1014), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1126), .A2(new_n965), .A3(G286), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1001), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT63), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1128), .B1(new_n1014), .B2(new_n1127), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1012), .A2(new_n1008), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n999), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1134), .B1(new_n1136), .B2(new_n978), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n967), .A2(new_n970), .A3(new_n977), .ZN(new_n1138));
  AOI211_X1 g713(.A(KEYINPUT119), .B(new_n1138), .C1(new_n1135), .C2(new_n999), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1125), .A2(KEYINPUT63), .A3(new_n1127), .ZN(new_n1141));
  OAI22_X1  g716(.A1(new_n1132), .A2(new_n1133), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1125), .A2(new_n1138), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n977), .A2(new_n962), .A3(new_n703), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(G1981), .B2(G305), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT116), .ZN(new_n1146));
  AOI211_X1 g721(.A(new_n965), .B(new_n964), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1143), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1124), .A2(new_n1142), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n1151));
  XNOR2_X1  g726(.A(G290), .B(G1986), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n947), .B1(new_n935), .B2(new_n1152), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1151), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n961), .B1(new_n1154), .B2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g731(.A1(new_n680), .A2(G319), .ZN(new_n1158));
  NOR3_X1   g732(.A1(G229), .A2(G401), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g733(.A1(new_n921), .A2(new_n858), .A3(new_n1159), .ZN(G225));
  INV_X1    g734(.A(G225), .ZN(G308));
endmodule


