

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755;

  NOR2_X1 U371 ( .A1(n677), .A2(n584), .ZN(n675) );
  XNOR2_X1 U372 ( .A(n377), .B(n376), .ZN(n375) );
  XNOR2_X1 U373 ( .A(n532), .B(n400), .ZN(n376) );
  XNOR2_X1 U374 ( .A(n733), .B(n416), .ZN(n532) );
  AND2_X1 U375 ( .A1(n674), .A2(n675), .ZN(n599) );
  XNOR2_X1 U376 ( .A(n535), .B(G469), .ZN(n557) );
  XNOR2_X2 U377 ( .A(G128), .B(G143), .ZN(n457) );
  INV_X2 U378 ( .A(G953), .ZN(n741) );
  XNOR2_X1 U379 ( .A(G116), .B(G107), .ZN(n404) );
  NOR2_X1 U380 ( .A1(n622), .A2(n740), .ZN(n625) );
  AND2_X1 U381 ( .A1(n395), .A2(n355), .ZN(n621) );
  NOR2_X1 U382 ( .A1(n668), .A2(n667), .ZN(n388) );
  NAND2_X1 U383 ( .A1(n384), .A2(n675), .ZN(n596) );
  XNOR2_X1 U384 ( .A(n404), .B(G122), .ZN(n399) );
  XNOR2_X1 U385 ( .A(G119), .B(KEYINPUT69), .ZN(n492) );
  XNOR2_X1 U386 ( .A(n621), .B(KEYINPUT85), .ZN(n740) );
  NAND2_X1 U387 ( .A1(n363), .A2(n408), .ZN(n640) );
  XNOR2_X1 U388 ( .A(n441), .B(n440), .ZN(n439) );
  OR2_X1 U389 ( .A1(n750), .A2(n751), .ZN(n441) );
  AND2_X1 U390 ( .A1(n572), .A2(n647), .ZN(n549) );
  INV_X1 U391 ( .A(n405), .ZN(n645) );
  AND2_X1 U392 ( .A1(n431), .A2(n429), .ZN(n428) );
  XNOR2_X1 U393 ( .A(n596), .B(n546), .ZN(n551) );
  NOR2_X1 U394 ( .A1(n419), .A2(n417), .ZN(n589) );
  AND2_X1 U395 ( .A1(n426), .A2(n425), .ZN(n424) );
  XNOR2_X1 U396 ( .A(n558), .B(n412), .ZN(n606) );
  NAND2_X1 U397 ( .A1(n434), .A2(KEYINPUT88), .ZN(n421) );
  XNOR2_X1 U398 ( .A(n373), .B(n371), .ZN(n377) );
  XNOR2_X1 U399 ( .A(n382), .B(n372), .ZN(n371) );
  NAND2_X1 U400 ( .A1(n370), .A2(n369), .ZN(n382) );
  XNOR2_X1 U401 ( .A(n381), .B(n380), .ZN(n383) );
  XNOR2_X1 U402 ( .A(n399), .B(n379), .ZN(n378) );
  XNOR2_X1 U403 ( .A(n494), .B(n492), .ZN(n381) );
  XNOR2_X1 U404 ( .A(n403), .B(n402), .ZN(n379) );
  XNOR2_X1 U405 ( .A(G110), .B(G104), .ZN(n733) );
  XNOR2_X1 U406 ( .A(KEYINPUT90), .B(KEYINPUT18), .ZN(n372) );
  XNOR2_X1 U407 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n374) );
  XNOR2_X1 U408 ( .A(KEYINPUT74), .B(KEYINPUT16), .ZN(n403) );
  XNOR2_X1 U409 ( .A(G113), .B(G101), .ZN(n494) );
  XOR2_X1 U410 ( .A(G902), .B(KEYINPUT15), .Z(n623) );
  NOR2_X1 U411 ( .A1(n661), .A2(n626), .ZN(n349) );
  NOR2_X2 U412 ( .A1(n661), .A2(n626), .ZN(n722) );
  BUF_X1 U413 ( .A(n401), .Z(n350) );
  NAND2_X1 U414 ( .A1(n428), .A2(n424), .ZN(n401) );
  NAND2_X1 U415 ( .A1(n427), .A2(n361), .ZN(n426) );
  BUF_X1 U416 ( .A(n600), .Z(n351) );
  BUF_X1 U417 ( .A(n353), .Z(n352) );
  XNOR2_X1 U418 ( .A(n732), .B(n375), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n732), .B(n375), .ZN(n703) );
  XNOR2_X1 U420 ( .A(n396), .B(n566), .ZN(n395) );
  XNOR2_X1 U421 ( .A(KEYINPUT67), .B(KEYINPUT48), .ZN(n566) );
  NAND2_X1 U422 ( .A1(n442), .A2(n439), .ZN(n396) );
  XNOR2_X1 U423 ( .A(n443), .B(n359), .ZN(n558) );
  OR2_X1 U424 ( .A1(n627), .A2(G902), .ZN(n443) );
  XNOR2_X1 U425 ( .A(n591), .B(KEYINPUT87), .ZN(n455) );
  XNOR2_X1 U426 ( .A(G128), .B(G137), .ZN(n514) );
  XNOR2_X1 U427 ( .A(G119), .B(G110), .ZN(n511) );
  NOR2_X1 U428 ( .A1(G953), .A2(G237), .ZN(n501) );
  XNOR2_X1 U429 ( .A(n493), .B(n411), .ZN(n380) );
  INV_X1 U430 ( .A(KEYINPUT3), .ZN(n493) );
  NAND2_X1 U431 ( .A1(n459), .A2(n664), .ZN(n668) );
  NAND2_X1 U432 ( .A1(n395), .A2(n356), .ZN(n574) );
  NOR2_X1 U433 ( .A1(n393), .A2(n394), .ZN(n392) );
  INV_X1 U434 ( .A(KEYINPUT2), .ZN(n394) );
  XNOR2_X1 U435 ( .A(n524), .B(n523), .ZN(n677) );
  XNOR2_X1 U436 ( .A(n522), .B(n521), .ZN(n523) );
  INV_X1 U437 ( .A(KEYINPUT25), .ZN(n521) );
  XOR2_X1 U438 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n465) );
  INV_X1 U439 ( .A(G134), .ZN(n462) );
  XNOR2_X1 U440 ( .A(n449), .B(n468), .ZN(n448) );
  XNOR2_X1 U441 ( .A(n534), .B(n454), .ZN(n708) );
  XNOR2_X1 U442 ( .A(n533), .B(n360), .ZN(n454) );
  XNOR2_X1 U443 ( .A(KEYINPUT89), .B(KEYINPUT33), .ZN(n581) );
  NAND2_X1 U444 ( .A1(n418), .A2(n414), .ZN(n417) );
  INV_X1 U445 ( .A(n606), .ZN(n418) );
  XNOR2_X1 U446 ( .A(n587), .B(n367), .ZN(n456) );
  XNOR2_X1 U447 ( .A(n401), .B(n358), .ZN(n406) );
  OR2_X1 U448 ( .A1(n390), .A2(n357), .ZN(n550) );
  INV_X1 U449 ( .A(KEYINPUT28), .ZN(n391) );
  BUF_X1 U450 ( .A(n558), .Z(n681) );
  BUF_X1 U451 ( .A(n677), .Z(n414) );
  INV_X1 U452 ( .A(KEYINPUT46), .ZN(n440) );
  INV_X1 U453 ( .A(KEYINPUT68), .ZN(n411) );
  NOR2_X1 U454 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U455 ( .A(KEYINPUT21), .B(n526), .ZN(n678) );
  OR2_X1 U456 ( .A1(G237), .A2(G902), .ZN(n497) );
  NAND2_X1 U457 ( .A1(n354), .A2(n623), .ZN(n434) );
  INV_X1 U458 ( .A(KEYINPUT107), .ZN(n450) );
  XNOR2_X1 U459 ( .A(G107), .B(G140), .ZN(n458) );
  INV_X1 U460 ( .A(KEYINPUT38), .ZN(n436) );
  INV_X1 U461 ( .A(KEYINPUT88), .ZN(n430) );
  XNOR2_X1 U462 ( .A(n579), .B(KEYINPUT94), .ZN(n580) );
  XNOR2_X1 U463 ( .A(n364), .B(n504), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n415), .B(n513), .ZN(n516) );
  XNOR2_X1 U465 ( .A(n511), .B(n510), .ZN(n513) );
  XNOR2_X1 U466 ( .A(n512), .B(n514), .ZN(n415) );
  XOR2_X1 U467 ( .A(G104), .B(G113), .Z(n483) );
  XNOR2_X1 U468 ( .A(G140), .B(KEYINPUT10), .ZN(n481) );
  XNOR2_X1 U469 ( .A(n457), .B(n374), .ZN(n373) );
  INV_X1 U470 ( .A(KEYINPUT71), .ZN(n416) );
  NAND2_X1 U471 ( .A1(n741), .A2(G224), .ZN(n400) );
  INV_X1 U472 ( .A(KEYINPUT73), .ZN(n402) );
  XNOR2_X1 U473 ( .A(n388), .B(KEYINPUT41), .ZN(n695) );
  INV_X1 U474 ( .A(KEYINPUT86), .ZN(n573) );
  INV_X1 U475 ( .A(n695), .ZN(n387) );
  INV_X1 U476 ( .A(KEYINPUT91), .ZN(n410) );
  INV_X1 U477 ( .A(KEYINPUT6), .ZN(n412) );
  XNOR2_X1 U478 ( .A(n467), .B(n447), .ZN(n720) );
  XNOR2_X1 U479 ( .A(n463), .B(n448), .ZN(n447) );
  NOR2_X1 U480 ( .A1(G952), .A2(n741), .ZN(n726) );
  XNOR2_X1 U481 ( .A(n446), .B(n445), .ZN(n751) );
  XNOR2_X1 U482 ( .A(KEYINPUT117), .B(KEYINPUT42), .ZN(n445) );
  NAND2_X1 U483 ( .A1(n389), .A2(n387), .ZN(n446) );
  INV_X1 U484 ( .A(n550), .ZN(n389) );
  NOR2_X1 U485 ( .A1(n681), .A2(n409), .ZN(n408) );
  INV_X1 U486 ( .A(n414), .ZN(n409) );
  INV_X1 U487 ( .A(n437), .ZN(n656) );
  XOR2_X1 U488 ( .A(n496), .B(n495), .Z(n354) );
  AND2_X1 U489 ( .A1(n437), .A2(n655), .ZN(n355) );
  AND2_X1 U490 ( .A1(n437), .A2(n392), .ZN(n356) );
  XNOR2_X1 U491 ( .A(n384), .B(KEYINPUT115), .ZN(n357) );
  XOR2_X1 U492 ( .A(KEYINPUT19), .B(KEYINPUT76), .Z(n358) );
  XOR2_X1 U493 ( .A(G472), .B(KEYINPUT99), .Z(n359) );
  XOR2_X1 U494 ( .A(n531), .B(n530), .Z(n360) );
  AND2_X1 U495 ( .A1(n664), .A2(n430), .ZN(n361) );
  OR2_X1 U496 ( .A1(n604), .A2(n603), .ZN(n362) );
  AND2_X1 U497 ( .A1(n456), .A2(n588), .ZN(n363) );
  NAND2_X1 U498 ( .A1(n501), .A2(G210), .ZN(n364) );
  AND2_X1 U499 ( .A1(n541), .A2(n540), .ZN(n365) );
  OR2_X1 U500 ( .A1(n354), .A2(n623), .ZN(n366) );
  XOR2_X1 U501 ( .A(KEYINPUT22), .B(KEYINPUT72), .Z(n367) );
  XNOR2_X1 U502 ( .A(KEYINPUT35), .B(KEYINPUT77), .ZN(n368) );
  NAND2_X1 U503 ( .A1(n479), .A2(G146), .ZN(n369) );
  NAND2_X1 U504 ( .A1(n480), .A2(G125), .ZN(n370) );
  XNOR2_X2 U505 ( .A(n383), .B(n378), .ZN(n732) );
  XNOR2_X1 U506 ( .A(n382), .B(n481), .ZN(n739) );
  XNOR2_X1 U507 ( .A(n398), .B(n383), .ZN(n397) );
  XNOR2_X1 U508 ( .A(n535), .B(G469), .ZN(n384) );
  XNOR2_X1 U509 ( .A(G110), .B(G104), .ZN(n385) );
  NAND2_X1 U510 ( .A1(n703), .A2(n354), .ZN(n435) );
  NAND2_X1 U511 ( .A1(n435), .A2(n434), .ZN(n423) );
  BUF_X1 U512 ( .A(n732), .Z(n386) );
  XNOR2_X1 U513 ( .A(n534), .B(n397), .ZN(n627) );
  INV_X1 U514 ( .A(n423), .ZN(n433) );
  XNOR2_X1 U515 ( .A(n529), .B(n391), .ZN(n390) );
  INV_X1 U516 ( .A(n655), .ZN(n393) );
  XNOR2_X1 U517 ( .A(n399), .B(n450), .ZN(n449) );
  NOR2_X1 U518 ( .A1(n562), .A2(n350), .ZN(n563) );
  XNOR2_X1 U519 ( .A(n444), .B(KEYINPUT0), .ZN(n586) );
  INV_X1 U520 ( .A(n586), .ZN(n600) );
  OR2_X2 U521 ( .A1(n708), .A2(G902), .ZN(n535) );
  XNOR2_X2 U522 ( .A(n557), .B(KEYINPUT1), .ZN(n674) );
  NOR2_X2 U523 ( .A1(n406), .A2(n580), .ZN(n444) );
  OR2_X1 U524 ( .A1(n550), .A2(n406), .ZN(n405) );
  NAND2_X1 U525 ( .A1(n547), .A2(n552), .ZN(n413) );
  XNOR2_X1 U526 ( .A(n413), .B(KEYINPUT39), .ZN(n572) );
  NAND2_X1 U527 ( .A1(n456), .A2(n407), .ZN(n590) );
  XNOR2_X1 U528 ( .A(n589), .B(KEYINPUT78), .ZN(n407) );
  NAND2_X1 U529 ( .A1(n599), .A2(n606), .ZN(n582) );
  XNOR2_X1 U530 ( .A(n588), .B(n410), .ZN(n419) );
  NAND2_X1 U531 ( .A1(n586), .A2(n585), .ZN(n587) );
  INV_X1 U532 ( .A(n457), .ZN(n491) );
  NAND2_X1 U533 ( .A1(n420), .A2(n432), .ZN(n431) );
  NOR2_X1 U534 ( .A1(n422), .A2(n421), .ZN(n420) );
  INV_X1 U535 ( .A(n435), .ZN(n422) );
  OR2_X2 U536 ( .A1(n353), .A2(n366), .ZN(n432) );
  NAND2_X1 U537 ( .A1(n423), .A2(n361), .ZN(n429) );
  NAND2_X1 U538 ( .A1(n433), .A2(n432), .ZN(n438) );
  OR2_X1 U539 ( .A1(n664), .A2(n430), .ZN(n425) );
  INV_X1 U540 ( .A(n432), .ZN(n427) );
  XNOR2_X1 U541 ( .A(n438), .B(n436), .ZN(n459) );
  NAND2_X1 U542 ( .A1(n583), .A2(n438), .ZN(n555) );
  OR2_X1 U543 ( .A1(n571), .A2(n438), .ZN(n437) );
  AND2_X1 U544 ( .A1(n565), .A2(n365), .ZN(n442) );
  AND2_X2 U545 ( .A1(n749), .A2(KEYINPUT64), .ZN(n592) );
  XNOR2_X2 U546 ( .A(n582), .B(n581), .ZN(n694) );
  XNOR2_X1 U547 ( .A(n453), .B(KEYINPUT34), .ZN(n452) );
  NAND2_X1 U548 ( .A1(n452), .A2(n583), .ZN(n451) );
  XNOR2_X2 U549 ( .A(n451), .B(n368), .ZN(n749) );
  NOR2_X2 U550 ( .A1(n694), .A2(n600), .ZN(n453) );
  XNOR2_X2 U551 ( .A(n738), .B(G146), .ZN(n534) );
  NAND2_X1 U552 ( .A1(n592), .A2(n455), .ZN(n594) );
  NAND2_X1 U553 ( .A1(n455), .A2(n595), .ZN(n605) );
  NOR2_X1 U554 ( .A1(n717), .A2(n726), .ZN(n718) );
  XNOR2_X2 U555 ( .A(n616), .B(KEYINPUT75), .ZN(n661) );
  XNOR2_X2 U556 ( .A(n500), .B(n499), .ZN(n738) );
  XNOR2_X1 U557 ( .A(n352), .B(n702), .ZN(n704) );
  INV_X1 U558 ( .A(KEYINPUT24), .ZN(n510) );
  INV_X1 U559 ( .A(KEYINPUT84), .ZN(n619) );
  XNOR2_X1 U560 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U561 ( .A(n574), .B(n573), .ZN(n615) );
  INV_X1 U562 ( .A(KEYINPUT114), .ZN(n546) );
  XNOR2_X1 U563 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U564 ( .A(n631), .B(n630), .ZN(n632) );
  XOR2_X1 U565 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n461) );
  XNOR2_X1 U566 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n460) );
  XNOR2_X1 U567 ( .A(n461), .B(n460), .ZN(n468) );
  XNOR2_X2 U568 ( .A(n491), .B(n462), .ZN(n500) );
  XNOR2_X1 U569 ( .A(n500), .B(KEYINPUT106), .ZN(n463) );
  NAND2_X1 U570 ( .A1(G234), .A2(n741), .ZN(n464) );
  XNOR2_X1 U571 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U572 ( .A(KEYINPUT82), .B(n466), .ZN(n517) );
  NAND2_X1 U573 ( .A1(G217), .A2(n517), .ZN(n467) );
  NOR2_X1 U574 ( .A1(G902), .A2(n720), .ZN(n470) );
  XNOR2_X1 U575 ( .A(KEYINPUT110), .B(G478), .ZN(n469) );
  XNOR2_X1 U576 ( .A(n470), .B(n469), .ZN(n554) );
  XOR2_X1 U577 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n472) );
  XNOR2_X1 U578 ( .A(KEYINPUT13), .B(G475), .ZN(n471) );
  XNOR2_X1 U579 ( .A(n472), .B(n471), .ZN(n488) );
  XOR2_X1 U580 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n474) );
  NAND2_X1 U581 ( .A1(G214), .A2(n501), .ZN(n473) );
  XNOR2_X1 U582 ( .A(n474), .B(n473), .ZN(n478) );
  XOR2_X1 U583 ( .A(KEYINPUT103), .B(KEYINPUT11), .Z(n476) );
  XNOR2_X1 U584 ( .A(G122), .B(KEYINPUT12), .ZN(n475) );
  XNOR2_X1 U585 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U586 ( .A(n478), .B(n477), .Z(n486) );
  INV_X1 U587 ( .A(G125), .ZN(n479) );
  INV_X1 U588 ( .A(G146), .ZN(n480) );
  XNOR2_X1 U589 ( .A(G143), .B(G131), .ZN(n482) );
  XNOR2_X1 U590 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U591 ( .A(n739), .B(n484), .ZN(n485) );
  XNOR2_X1 U592 ( .A(n486), .B(n485), .ZN(n714) );
  NOR2_X1 U593 ( .A1(G902), .A2(n714), .ZN(n487) );
  XOR2_X1 U594 ( .A(n488), .B(n487), .Z(n553) );
  INV_X1 U595 ( .A(n553), .ZN(n489) );
  NAND2_X1 U596 ( .A1(n554), .A2(n489), .ZN(n561) );
  INV_X1 U597 ( .A(n561), .ZN(n647) );
  NOR2_X1 U598 ( .A1(n489), .A2(n554), .ZN(n490) );
  XOR2_X1 U599 ( .A(n490), .B(KEYINPUT111), .Z(n650) );
  NOR2_X1 U600 ( .A1(n647), .A2(n650), .ZN(n669) );
  INV_X1 U601 ( .A(n669), .ZN(n537) );
  NAND2_X1 U602 ( .A1(G210), .A2(n497), .ZN(n496) );
  INV_X1 U603 ( .A(KEYINPUT79), .ZN(n495) );
  NAND2_X1 U604 ( .A1(G214), .A2(n497), .ZN(n664) );
  XNOR2_X1 U605 ( .A(G131), .B(KEYINPUT4), .ZN(n498) );
  XNOR2_X1 U606 ( .A(n498), .B(G137), .ZN(n499) );
  XNOR2_X1 U607 ( .A(G116), .B(KEYINPUT5), .ZN(n503) );
  INV_X1 U608 ( .A(KEYINPUT98), .ZN(n502) );
  NAND2_X1 U609 ( .A1(G234), .A2(G237), .ZN(n505) );
  XNOR2_X1 U610 ( .A(n505), .B(KEYINPUT92), .ZN(n506) );
  XNOR2_X1 U611 ( .A(KEYINPUT14), .B(n506), .ZN(n507) );
  NAND2_X1 U612 ( .A1(G952), .A2(n507), .ZN(n693) );
  NOR2_X1 U613 ( .A1(G953), .A2(n693), .ZN(n578) );
  NAND2_X1 U614 ( .A1(G902), .A2(n507), .ZN(n576) );
  OR2_X1 U615 ( .A1(n741), .A2(n576), .ZN(n508) );
  NOR2_X1 U616 ( .A1(G900), .A2(n508), .ZN(n509) );
  NOR2_X1 U617 ( .A1(n578), .A2(n509), .ZN(n544) );
  XOR2_X1 U618 ( .A(KEYINPUT23), .B(KEYINPUT70), .Z(n512) );
  INV_X1 U619 ( .A(n739), .ZN(n515) );
  XNOR2_X1 U620 ( .A(n516), .B(n515), .ZN(n519) );
  NAND2_X1 U621 ( .A1(G221), .A2(n517), .ZN(n518) );
  XNOR2_X1 U622 ( .A(n519), .B(n518), .ZN(n724) );
  NOR2_X1 U623 ( .A1(G902), .A2(n724), .ZN(n524) );
  INV_X1 U624 ( .A(n623), .ZN(n617) );
  NAND2_X1 U625 ( .A1(n617), .A2(G234), .ZN(n520) );
  XNOR2_X1 U626 ( .A(n520), .B(KEYINPUT20), .ZN(n525) );
  NAND2_X1 U627 ( .A1(n525), .A2(G217), .ZN(n522) );
  NAND2_X1 U628 ( .A1(n525), .A2(G221), .ZN(n526) );
  INV_X1 U629 ( .A(n678), .ZN(n527) );
  NAND2_X1 U630 ( .A1(n677), .A2(n527), .ZN(n528) );
  NOR2_X1 U631 ( .A1(n544), .A2(n528), .ZN(n559) );
  AND2_X1 U632 ( .A1(n681), .A2(n559), .ZN(n529) );
  XOR2_X1 U633 ( .A(G101), .B(KEYINPUT95), .Z(n531) );
  NAND2_X1 U634 ( .A1(G227), .A2(n741), .ZN(n530) );
  XNOR2_X1 U635 ( .A(n532), .B(n458), .ZN(n533) );
  NAND2_X1 U636 ( .A1(n537), .A2(n645), .ZN(n536) );
  NAND2_X1 U637 ( .A1(n536), .A2(KEYINPUT47), .ZN(n541) );
  XNOR2_X1 U638 ( .A(KEYINPUT81), .B(n537), .ZN(n604) );
  XOR2_X1 U639 ( .A(KEYINPUT65), .B(KEYINPUT47), .Z(n538) );
  NOR2_X1 U640 ( .A1(n604), .A2(n538), .ZN(n539) );
  NAND2_X1 U641 ( .A1(n539), .A2(n645), .ZN(n540) );
  INV_X1 U642 ( .A(KEYINPUT30), .ZN(n543) );
  AND2_X1 U643 ( .A1(n558), .A2(n664), .ZN(n542) );
  XNOR2_X1 U644 ( .A(n543), .B(n542), .ZN(n545) );
  NOR2_X1 U645 ( .A1(n545), .A2(n544), .ZN(n552) );
  XNOR2_X1 U646 ( .A(KEYINPUT96), .B(n678), .ZN(n584) );
  AND2_X1 U647 ( .A1(n551), .A2(n459), .ZN(n547) );
  XNOR2_X1 U648 ( .A(KEYINPUT40), .B(KEYINPUT116), .ZN(n548) );
  XNOR2_X1 U649 ( .A(n549), .B(n548), .ZN(n750) );
  NAND2_X1 U650 ( .A1(n554), .A2(n553), .ZN(n667) );
  NAND2_X1 U651 ( .A1(n552), .A2(n551), .ZN(n556) );
  NOR2_X1 U652 ( .A1(n554), .A2(n553), .ZN(n583) );
  NOR2_X1 U653 ( .A1(n556), .A2(n555), .ZN(n644) );
  NAND2_X1 U654 ( .A1(n606), .A2(n559), .ZN(n560) );
  NOR2_X1 U655 ( .A1(n561), .A2(n560), .ZN(n567) );
  INV_X1 U656 ( .A(n567), .ZN(n562) );
  XOR2_X1 U657 ( .A(KEYINPUT36), .B(n563), .Z(n564) );
  NOR2_X1 U658 ( .A1(n419), .A2(n564), .ZN(n653) );
  NOR2_X1 U659 ( .A1(n644), .A2(n653), .ZN(n565) );
  NAND2_X1 U660 ( .A1(n567), .A2(n664), .ZN(n568) );
  XOR2_X1 U661 ( .A(KEYINPUT113), .B(n568), .Z(n569) );
  NOR2_X1 U662 ( .A1(n674), .A2(n569), .ZN(n570) );
  XNOR2_X1 U663 ( .A(n570), .B(KEYINPUT43), .ZN(n571) );
  NAND2_X1 U664 ( .A1(n650), .A2(n572), .ZN(n655) );
  NOR2_X1 U665 ( .A1(G898), .A2(n741), .ZN(n575) );
  XNOR2_X1 U666 ( .A(KEYINPUT93), .B(n575), .ZN(n735) );
  NOR2_X1 U667 ( .A1(n735), .A2(n576), .ZN(n577) );
  NOR2_X1 U668 ( .A1(n578), .A2(n577), .ZN(n579) );
  INV_X1 U669 ( .A(n674), .ZN(n588) );
  NOR2_X1 U670 ( .A1(n667), .A2(n584), .ZN(n585) );
  XNOR2_X1 U671 ( .A(n590), .B(KEYINPUT32), .ZN(n752) );
  NAND2_X1 U672 ( .A1(n640), .A2(n752), .ZN(n591) );
  INV_X1 U673 ( .A(KEYINPUT44), .ZN(n593) );
  XNOR2_X1 U674 ( .A(n594), .B(n593), .ZN(n612) );
  NOR2_X1 U675 ( .A1(KEYINPUT64), .A2(n749), .ZN(n595) );
  NOR2_X1 U676 ( .A1(n600), .A2(n596), .ZN(n597) );
  XNOR2_X1 U677 ( .A(n597), .B(KEYINPUT97), .ZN(n598) );
  NOR2_X1 U678 ( .A1(n681), .A2(n598), .ZN(n636) );
  NAND2_X1 U679 ( .A1(n681), .A2(n599), .ZN(n686) );
  NOR2_X1 U680 ( .A1(n351), .A2(n686), .ZN(n602) );
  XOR2_X1 U681 ( .A(KEYINPUT31), .B(KEYINPUT100), .Z(n601) );
  XNOR2_X1 U682 ( .A(n602), .B(n601), .ZN(n651) );
  NOR2_X1 U683 ( .A1(n636), .A2(n651), .ZN(n603) );
  NAND2_X1 U684 ( .A1(n605), .A2(n362), .ZN(n610) );
  NOR2_X1 U685 ( .A1(n606), .A2(n414), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n363), .A2(n607), .ZN(n608) );
  XNOR2_X1 U687 ( .A(KEYINPUT112), .B(n608), .ZN(n755) );
  INV_X1 U688 ( .A(n755), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n614) );
  INV_X1 U690 ( .A(KEYINPUT45), .ZN(n613) );
  XNOR2_X1 U691 ( .A(n614), .B(n613), .ZN(n618) );
  BUF_X1 U692 ( .A(n618), .Z(n657) );
  INV_X1 U693 ( .A(n657), .ZN(n729) );
  NAND2_X1 U694 ( .A1(n615), .A2(n729), .ZN(n616) );
  NOR2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n620) );
  XNOR2_X1 U696 ( .A(n620), .B(n619), .ZN(n622) );
  AND2_X1 U697 ( .A1(n623), .A2(KEYINPUT2), .ZN(n624) );
  NOR2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U699 ( .A1(n722), .A2(G472), .ZN(n631) );
  XNOR2_X1 U700 ( .A(n627), .B(KEYINPUT119), .ZN(n629) );
  XOR2_X1 U701 ( .A(KEYINPUT62), .B(KEYINPUT118), .Z(n628) );
  NOR2_X1 U702 ( .A1(n632), .A2(n726), .ZN(n634) );
  INV_X1 U703 ( .A(KEYINPUT63), .ZN(n633) );
  XNOR2_X1 U704 ( .A(n634), .B(n633), .ZN(G57) );
  NAND2_X1 U705 ( .A1(n647), .A2(n636), .ZN(n635) );
  XNOR2_X1 U706 ( .A(G104), .B(n635), .ZN(G6) );
  XOR2_X1 U707 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n638) );
  NAND2_X1 U708 ( .A1(n636), .A2(n650), .ZN(n637) );
  XNOR2_X1 U709 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U710 ( .A(G107), .B(n639), .ZN(G9) );
  XNOR2_X1 U711 ( .A(n640), .B(G110), .ZN(G12) );
  XOR2_X1 U712 ( .A(KEYINPUT120), .B(KEYINPUT29), .Z(n642) );
  NAND2_X1 U713 ( .A1(n645), .A2(n650), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U715 ( .A(G128), .B(n643), .ZN(G30) );
  XOR2_X1 U716 ( .A(G143), .B(n644), .Z(G45) );
  NAND2_X1 U717 ( .A1(n645), .A2(n647), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n646), .B(G146), .ZN(G48) );
  XOR2_X1 U719 ( .A(G113), .B(KEYINPUT121), .Z(n649) );
  NAND2_X1 U720 ( .A1(n647), .A2(n651), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n649), .B(n648), .ZN(G15) );
  NAND2_X1 U722 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n652), .B(G116), .ZN(G18) );
  XNOR2_X1 U724 ( .A(G125), .B(n653), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n654), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U726 ( .A(G134), .B(n655), .ZN(G36) );
  XOR2_X1 U727 ( .A(G140), .B(n656), .Z(G42) );
  XOR2_X1 U728 ( .A(KEYINPUT80), .B(KEYINPUT2), .Z(n658) );
  NAND2_X1 U729 ( .A1(n657), .A2(n658), .ZN(n663) );
  NAND2_X1 U730 ( .A1(n658), .A2(n740), .ZN(n659) );
  XNOR2_X1 U731 ( .A(KEYINPUT83), .B(n659), .ZN(n660) );
  NOR2_X1 U732 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U733 ( .A1(n663), .A2(n662), .ZN(n699) );
  NOR2_X1 U734 ( .A1(n459), .A2(n664), .ZN(n665) );
  XOR2_X1 U735 ( .A(KEYINPUT123), .B(n665), .Z(n666) );
  NOR2_X1 U736 ( .A1(n667), .A2(n666), .ZN(n671) );
  NOR2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n672), .B(KEYINPUT124), .ZN(n673) );
  NOR2_X1 U740 ( .A1(n694), .A2(n673), .ZN(n690) );
  NOR2_X1 U741 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U742 ( .A(KEYINPUT50), .B(n676), .Z(n684) );
  NAND2_X1 U743 ( .A1(n678), .A2(n414), .ZN(n679) );
  XNOR2_X1 U744 ( .A(KEYINPUT49), .B(n679), .ZN(n680) );
  NOR2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U746 ( .A(KEYINPUT122), .B(n682), .ZN(n683) );
  NAND2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U748 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U749 ( .A(KEYINPUT51), .B(n687), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n695), .A2(n688), .ZN(n689) );
  NOR2_X1 U751 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U752 ( .A(n691), .B(KEYINPUT52), .ZN(n692) );
  NOR2_X1 U753 ( .A1(n693), .A2(n692), .ZN(n697) );
  NOR2_X1 U754 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U755 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U756 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U757 ( .A1(n700), .A2(G953), .ZN(n701) );
  XNOR2_X1 U758 ( .A(n701), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U759 ( .A1(n722), .A2(G210), .ZN(n705) );
  XOR2_X1 U760 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n702) );
  XNOR2_X1 U761 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U762 ( .A1(n706), .A2(n726), .ZN(n707) );
  XNOR2_X1 U763 ( .A(n707), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U764 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n710) );
  XNOR2_X1 U765 ( .A(n708), .B(KEYINPUT125), .ZN(n709) );
  XNOR2_X1 U766 ( .A(n710), .B(n709), .ZN(n712) );
  NAND2_X1 U767 ( .A1(n349), .A2(G469), .ZN(n711) );
  XOR2_X1 U768 ( .A(n712), .B(n711), .Z(n713) );
  NOR2_X1 U769 ( .A1(n726), .A2(n713), .ZN(G54) );
  XOR2_X1 U770 ( .A(n714), .B(KEYINPUT59), .Z(n716) );
  NAND2_X1 U771 ( .A1(n722), .A2(G475), .ZN(n715) );
  XNOR2_X1 U772 ( .A(n715), .B(n716), .ZN(n717) );
  XNOR2_X1 U773 ( .A(n718), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U774 ( .A1(G478), .A2(n349), .ZN(n719) );
  XNOR2_X1 U775 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U776 ( .A1(n726), .A2(n721), .ZN(G63) );
  NAND2_X1 U777 ( .A1(G217), .A2(n349), .ZN(n723) );
  XNOR2_X1 U778 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U779 ( .A1(n726), .A2(n725), .ZN(G66) );
  NAND2_X1 U780 ( .A1(G953), .A2(G224), .ZN(n727) );
  XNOR2_X1 U781 ( .A(KEYINPUT61), .B(n727), .ZN(n728) );
  NAND2_X1 U782 ( .A1(n728), .A2(G898), .ZN(n731) );
  NAND2_X1 U783 ( .A1(n729), .A2(n741), .ZN(n730) );
  NAND2_X1 U784 ( .A1(n731), .A2(n730), .ZN(n737) );
  XNOR2_X1 U785 ( .A(n385), .B(n386), .ZN(n734) );
  NAND2_X1 U786 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U787 ( .A(n737), .B(n736), .Z(G69) );
  XNOR2_X1 U788 ( .A(n738), .B(n739), .ZN(n743) );
  XNOR2_X1 U789 ( .A(n740), .B(n743), .ZN(n742) );
  NAND2_X1 U790 ( .A1(n742), .A2(n741), .ZN(n747) );
  XNOR2_X1 U791 ( .A(G227), .B(n743), .ZN(n744) );
  NAND2_X1 U792 ( .A1(n744), .A2(G900), .ZN(n745) );
  NAND2_X1 U793 ( .A1(n745), .A2(G953), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U795 ( .A(KEYINPUT126), .B(n748), .ZN(G72) );
  XNOR2_X1 U796 ( .A(n749), .B(G122), .ZN(G24) );
  XOR2_X1 U797 ( .A(G131), .B(n750), .Z(G33) );
  XOR2_X1 U798 ( .A(G137), .B(n751), .Z(G39) );
  BUF_X1 U799 ( .A(n752), .Z(n753) );
  XOR2_X1 U800 ( .A(G119), .B(n753), .Z(n754) );
  XNOR2_X1 U801 ( .A(KEYINPUT127), .B(n754), .ZN(G21) );
  XNOR2_X1 U802 ( .A(G101), .B(n755), .ZN(G3) );
endmodule

