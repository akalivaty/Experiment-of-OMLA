

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U551 ( .A(KEYINPUT27), .B(n588), .Z(n515) );
  OR2_X1 U552 ( .A1(n689), .A2(n688), .ZN(n516) );
  OR2_X1 U553 ( .A1(n682), .A2(n681), .ZN(n517) );
  AND2_X1 U554 ( .A1(n633), .A2(G1996), .ZN(n605) );
  NOR2_X1 U555 ( .A1(n915), .A2(n608), .ZN(n609) );
  INV_X1 U556 ( .A(KEYINPUT89), .ZN(n587) );
  INV_X1 U557 ( .A(KEYINPUT28), .ZN(n591) );
  INV_X1 U558 ( .A(KEYINPUT29), .ZN(n630) );
  XNOR2_X1 U559 ( .A(n631), .B(n630), .ZN(n638) );
  NOR2_X1 U560 ( .A1(n648), .A2(n647), .ZN(n649) );
  AND2_X1 U561 ( .A1(n690), .A2(n516), .ZN(n691) );
  AND2_X1 U562 ( .A1(n522), .A2(G2104), .ZN(n884) );
  NOR2_X1 U563 ( .A1(G651), .A2(n562), .ZN(n775) );
  NOR2_X1 U564 ( .A1(n526), .A2(n525), .ZN(G160) );
  AND2_X1 U565 ( .A1(G2105), .A2(G2104), .ZN(n881) );
  NAND2_X1 U566 ( .A1(n881), .A2(G113), .ZN(n520) );
  INV_X1 U567 ( .A(G2105), .ZN(n522) );
  NAND2_X1 U568 ( .A1(G101), .A2(n884), .ZN(n518) );
  XOR2_X1 U569 ( .A(KEYINPUT23), .B(n518), .Z(n519) );
  NAND2_X1 U570 ( .A1(n520), .A2(n519), .ZN(n526) );
  NOR2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XOR2_X2 U572 ( .A(KEYINPUT17), .B(n521), .Z(n885) );
  NAND2_X1 U573 ( .A1(G137), .A2(n885), .ZN(n524) );
  NOR2_X1 U574 ( .A1(G2104), .A2(n522), .ZN(n880) );
  NAND2_X1 U575 ( .A1(G125), .A2(n880), .ZN(n523) );
  NAND2_X1 U576 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U577 ( .A1(G102), .A2(n884), .ZN(n528) );
  NAND2_X1 U578 ( .A1(G138), .A2(n885), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n532) );
  NAND2_X1 U580 ( .A1(G126), .A2(n880), .ZN(n530) );
  NAND2_X1 U581 ( .A1(G114), .A2(n881), .ZN(n529) );
  NAND2_X1 U582 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U583 ( .A1(n532), .A2(n531), .ZN(G164) );
  INV_X1 U584 ( .A(G651), .ZN(n537) );
  NOR2_X1 U585 ( .A1(G543), .A2(n537), .ZN(n533) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n533), .Z(n774) );
  NAND2_X1 U587 ( .A1(G64), .A2(n774), .ZN(n535) );
  XOR2_X1 U588 ( .A(KEYINPUT0), .B(G543), .Z(n562) );
  NAND2_X1 U589 ( .A1(G52), .A2(n775), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n535), .A2(n534), .ZN(n542) );
  NOR2_X1 U591 ( .A1(G651), .A2(G543), .ZN(n536) );
  XOR2_X1 U592 ( .A(KEYINPUT65), .B(n536), .Z(n770) );
  NAND2_X1 U593 ( .A1(G90), .A2(n770), .ZN(n539) );
  NOR2_X1 U594 ( .A1(n562), .A2(n537), .ZN(n771) );
  NAND2_X1 U595 ( .A1(G77), .A2(n771), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U597 ( .A(KEYINPUT9), .B(n540), .Z(n541) );
  NOR2_X1 U598 ( .A1(n542), .A2(n541), .ZN(G171) );
  NAND2_X1 U599 ( .A1(n770), .A2(G89), .ZN(n543) );
  XNOR2_X1 U600 ( .A(n543), .B(KEYINPUT4), .ZN(n545) );
  NAND2_X1 U601 ( .A1(G76), .A2(n771), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U603 ( .A(n546), .B(KEYINPUT5), .ZN(n551) );
  NAND2_X1 U604 ( .A1(G63), .A2(n774), .ZN(n548) );
  NAND2_X1 U605 ( .A1(G51), .A2(n775), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U607 ( .A(KEYINPUT6), .B(n549), .Z(n550) );
  NAND2_X1 U608 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U609 ( .A(n552), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U610 ( .A1(G88), .A2(n770), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G75), .A2(n771), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G62), .A2(n774), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G50), .A2(n775), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U616 ( .A1(n558), .A2(n557), .ZN(G166) );
  INV_X1 U617 ( .A(G166), .ZN(G303) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U619 ( .A1(G49), .A2(n775), .ZN(n560) );
  NAND2_X1 U620 ( .A1(G74), .A2(G651), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U622 ( .A1(n774), .A2(n561), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n562), .A2(G87), .ZN(n563) );
  NAND2_X1 U624 ( .A1(n564), .A2(n563), .ZN(G288) );
  NAND2_X1 U625 ( .A1(G86), .A2(n770), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G61), .A2(n774), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n771), .A2(G73), .ZN(n567) );
  XOR2_X1 U629 ( .A(KEYINPUT2), .B(n567), .Z(n568) );
  NOR2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U631 ( .A(n570), .B(KEYINPUT72), .ZN(n572) );
  NAND2_X1 U632 ( .A1(G48), .A2(n775), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n572), .A2(n571), .ZN(G305) );
  NAND2_X1 U634 ( .A1(G85), .A2(n770), .ZN(n574) );
  NAND2_X1 U635 ( .A1(G72), .A2(n771), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G60), .A2(n774), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G47), .A2(n775), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n577) );
  OR2_X1 U640 ( .A1(n578), .A2(n577), .ZN(G290) );
  NAND2_X1 U641 ( .A1(G65), .A2(n774), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G53), .A2(n775), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U644 ( .A1(G91), .A2(n770), .ZN(n582) );
  NAND2_X1 U645 ( .A1(G78), .A2(n771), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U647 ( .A1(n584), .A2(n583), .ZN(n921) );
  NAND2_X1 U648 ( .A1(G40), .A2(G160), .ZN(n586) );
  INV_X1 U649 ( .A(KEYINPUT82), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n721) );
  NOR2_X1 U651 ( .A1(G164), .A2(G1384), .ZN(n722) );
  NAND2_X1 U652 ( .A1(n721), .A2(n722), .ZN(n604) );
  XNOR2_X1 U653 ( .A(n604), .B(n587), .ZN(n632) );
  NAND2_X1 U654 ( .A1(n632), .A2(G1956), .ZN(n589) );
  INV_X1 U655 ( .A(n632), .ZN(n617) );
  NAND2_X1 U656 ( .A1(n617), .A2(G2072), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n515), .ZN(n590) );
  XNOR2_X1 U658 ( .A(n590), .B(KEYINPUT91), .ZN(n593) );
  NOR2_X1 U659 ( .A1(n921), .A2(n593), .ZN(n592) );
  XNOR2_X1 U660 ( .A(n592), .B(n591), .ZN(n629) );
  NAND2_X1 U661 ( .A1(n921), .A2(n593), .ZN(n627) );
  XNOR2_X1 U662 ( .A(KEYINPUT67), .B(KEYINPUT13), .ZN(n598) );
  NAND2_X1 U663 ( .A1(n770), .A2(G81), .ZN(n594) );
  XNOR2_X1 U664 ( .A(n594), .B(KEYINPUT12), .ZN(n596) );
  NAND2_X1 U665 ( .A1(G68), .A2(n771), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U667 ( .A(n598), .B(n597), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n774), .A2(G56), .ZN(n599) );
  XOR2_X1 U669 ( .A(KEYINPUT14), .B(n599), .Z(n600) );
  NOR2_X1 U670 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U671 ( .A1(n775), .A2(G43), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n603), .A2(n602), .ZN(n915) );
  INV_X1 U673 ( .A(n604), .ZN(n633) );
  XOR2_X1 U674 ( .A(n605), .B(KEYINPUT26), .Z(n607) );
  INV_X1 U675 ( .A(n633), .ZN(n653) );
  NAND2_X1 U676 ( .A1(n653), .A2(G1341), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U678 ( .A(KEYINPUT64), .B(n609), .Z(n623) );
  NAND2_X1 U679 ( .A1(G92), .A2(n770), .ZN(n611) );
  NAND2_X1 U680 ( .A1(G79), .A2(n771), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U682 ( .A1(G66), .A2(n774), .ZN(n613) );
  NAND2_X1 U683 ( .A1(G54), .A2(n775), .ZN(n612) );
  NAND2_X1 U684 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U686 ( .A(KEYINPUT15), .B(n616), .Z(n899) );
  INV_X1 U687 ( .A(n899), .ZN(n929) );
  OR2_X1 U688 ( .A1(n623), .A2(n929), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G2067), .A2(n617), .ZN(n619) );
  NAND2_X1 U690 ( .A1(G1348), .A2(n653), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U692 ( .A(n620), .B(KEYINPUT92), .ZN(n621) );
  NAND2_X1 U693 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U694 ( .A1(n623), .A2(n929), .ZN(n624) );
  NAND2_X1 U695 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U697 ( .A1(n629), .A2(n628), .ZN(n631) );
  XOR2_X1 U698 ( .A(G2078), .B(KEYINPUT25), .Z(n966) );
  NOR2_X1 U699 ( .A1(n966), .A2(n632), .ZN(n635) );
  NOR2_X1 U700 ( .A1(n633), .A2(G1961), .ZN(n634) );
  NOR2_X1 U701 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U702 ( .A(KEYINPUT90), .B(n636), .Z(n639) );
  NAND2_X1 U703 ( .A1(G171), .A2(n639), .ZN(n637) );
  NAND2_X1 U704 ( .A1(n638), .A2(n637), .ZN(n660) );
  OR2_X1 U705 ( .A1(G171), .A2(n639), .ZN(n640) );
  XNOR2_X1 U706 ( .A(n640), .B(KEYINPUT93), .ZN(n645) );
  NOR2_X1 U707 ( .A1(G2084), .A2(n653), .ZN(n650) );
  NAND2_X1 U708 ( .A1(G8), .A2(n653), .ZN(n689) );
  NOR2_X1 U709 ( .A1(G1966), .A2(n689), .ZN(n647) );
  NOR2_X1 U710 ( .A1(n650), .A2(n647), .ZN(n641) );
  NAND2_X1 U711 ( .A1(G8), .A2(n641), .ZN(n642) );
  XNOR2_X1 U712 ( .A(KEYINPUT30), .B(n642), .ZN(n643) );
  NOR2_X1 U713 ( .A1(n643), .A2(G168), .ZN(n644) );
  NOR2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U715 ( .A(KEYINPUT31), .B(n646), .Z(n658) );
  AND2_X1 U716 ( .A1(n660), .A2(n658), .ZN(n648) );
  XNOR2_X1 U717 ( .A(n649), .B(KEYINPUT94), .ZN(n652) );
  NAND2_X1 U718 ( .A1(n650), .A2(G8), .ZN(n651) );
  NAND2_X1 U719 ( .A1(n652), .A2(n651), .ZN(n668) );
  NOR2_X1 U720 ( .A1(G1971), .A2(n689), .ZN(n655) );
  NOR2_X1 U721 ( .A1(G2090), .A2(n653), .ZN(n654) );
  NOR2_X1 U722 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U723 ( .A(KEYINPUT95), .B(n656), .Z(n657) );
  NAND2_X1 U724 ( .A1(n657), .A2(G303), .ZN(n661) );
  AND2_X1 U725 ( .A1(n658), .A2(n661), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n660), .A2(n659), .ZN(n665) );
  INV_X1 U727 ( .A(n661), .ZN(n662) );
  OR2_X1 U728 ( .A1(n662), .A2(G286), .ZN(n663) );
  AND2_X1 U729 ( .A1(G8), .A2(n663), .ZN(n664) );
  NAND2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U731 ( .A(n666), .B(KEYINPUT32), .ZN(n667) );
  NAND2_X1 U732 ( .A1(n668), .A2(n667), .ZN(n685) );
  NOR2_X1 U733 ( .A1(G1976), .A2(G288), .ZN(n677) );
  NOR2_X1 U734 ( .A1(G1971), .A2(G303), .ZN(n669) );
  NOR2_X1 U735 ( .A1(n677), .A2(n669), .ZN(n917) );
  INV_X1 U736 ( .A(KEYINPUT33), .ZN(n673) );
  AND2_X1 U737 ( .A1(n917), .A2(n673), .ZN(n670) );
  NAND2_X1 U738 ( .A1(n685), .A2(n670), .ZN(n675) );
  NAND2_X1 U739 ( .A1(G1976), .A2(G288), .ZN(n916) );
  INV_X1 U740 ( .A(n689), .ZN(n671) );
  NAND2_X1 U741 ( .A1(n916), .A2(n671), .ZN(n672) );
  NAND2_X1 U742 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n682) );
  XNOR2_X1 U744 ( .A(G1981), .B(KEYINPUT97), .ZN(n676) );
  XNOR2_X1 U745 ( .A(n676), .B(G305), .ZN(n912) );
  NAND2_X1 U746 ( .A1(KEYINPUT33), .A2(n677), .ZN(n678) );
  NOR2_X1 U747 ( .A1(n689), .A2(n678), .ZN(n679) );
  XOR2_X1 U748 ( .A(KEYINPUT96), .B(n679), .Z(n680) );
  NAND2_X1 U749 ( .A1(n912), .A2(n680), .ZN(n681) );
  NOR2_X1 U750 ( .A1(G2090), .A2(G303), .ZN(n683) );
  NAND2_X1 U751 ( .A1(G8), .A2(n683), .ZN(n684) );
  NAND2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U753 ( .A1(n689), .A2(n686), .ZN(n690) );
  NOR2_X1 U754 ( .A1(G1981), .A2(G305), .ZN(n687) );
  XOR2_X1 U755 ( .A(n687), .B(KEYINPUT24), .Z(n688) );
  NAND2_X1 U756 ( .A1(n517), .A2(n691), .ZN(n726) );
  NAND2_X1 U757 ( .A1(G104), .A2(n884), .ZN(n693) );
  NAND2_X1 U758 ( .A1(G140), .A2(n885), .ZN(n692) );
  NAND2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U760 ( .A(KEYINPUT34), .B(n694), .ZN(n700) );
  NAND2_X1 U761 ( .A1(n880), .A2(G128), .ZN(n695) );
  XNOR2_X1 U762 ( .A(n695), .B(KEYINPUT84), .ZN(n697) );
  NAND2_X1 U763 ( .A1(G116), .A2(n881), .ZN(n696) );
  NAND2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U765 ( .A(n698), .B(KEYINPUT35), .Z(n699) );
  NOR2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U767 ( .A(KEYINPUT36), .B(n701), .Z(n702) );
  XNOR2_X1 U768 ( .A(KEYINPUT85), .B(n702), .ZN(n870) );
  XOR2_X1 U769 ( .A(G2067), .B(KEYINPUT37), .Z(n703) );
  XNOR2_X1 U770 ( .A(KEYINPUT83), .B(n703), .ZN(n739) );
  NOR2_X1 U771 ( .A1(n870), .A2(n739), .ZN(n736) );
  XOR2_X1 U772 ( .A(KEYINPUT87), .B(G1991), .Z(n973) );
  NAND2_X1 U773 ( .A1(G119), .A2(n880), .ZN(n705) );
  NAND2_X1 U774 ( .A1(G107), .A2(n881), .ZN(n704) );
  NAND2_X1 U775 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U776 ( .A(KEYINPUT86), .B(n706), .Z(n710) );
  NAND2_X1 U777 ( .A1(G95), .A2(n884), .ZN(n708) );
  NAND2_X1 U778 ( .A1(G131), .A2(n885), .ZN(n707) );
  AND2_X1 U779 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U780 ( .A1(n710), .A2(n709), .ZN(n893) );
  NAND2_X1 U781 ( .A1(n973), .A2(n893), .ZN(n720) );
  NAND2_X1 U782 ( .A1(G129), .A2(n880), .ZN(n712) );
  NAND2_X1 U783 ( .A1(G117), .A2(n881), .ZN(n711) );
  NAND2_X1 U784 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U785 ( .A1(n884), .A2(G105), .ZN(n713) );
  XOR2_X1 U786 ( .A(KEYINPUT38), .B(n713), .Z(n714) );
  NOR2_X1 U787 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U788 ( .A(n716), .B(KEYINPUT88), .ZN(n718) );
  NAND2_X1 U789 ( .A1(G141), .A2(n885), .ZN(n717) );
  NAND2_X1 U790 ( .A1(n718), .A2(n717), .ZN(n872) );
  NAND2_X1 U791 ( .A1(G1996), .A2(n872), .ZN(n719) );
  NAND2_X1 U792 ( .A1(n720), .A2(n719), .ZN(n731) );
  NOR2_X1 U793 ( .A1(n736), .A2(n731), .ZN(n1009) );
  XOR2_X1 U794 ( .A(G1986), .B(G290), .Z(n932) );
  NAND2_X1 U795 ( .A1(n1009), .A2(n932), .ZN(n724) );
  INV_X1 U796 ( .A(n721), .ZN(n723) );
  NOR2_X1 U797 ( .A1(n723), .A2(n722), .ZN(n741) );
  NAND2_X1 U798 ( .A1(n724), .A2(n741), .ZN(n725) );
  NAND2_X1 U799 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U800 ( .A(n727), .B(KEYINPUT98), .ZN(n744) );
  NOR2_X1 U801 ( .A1(G1996), .A2(n872), .ZN(n728) );
  XOR2_X1 U802 ( .A(KEYINPUT99), .B(n728), .Z(n1004) );
  NOR2_X1 U803 ( .A1(n973), .A2(n893), .ZN(n993) );
  NOR2_X1 U804 ( .A1(G1986), .A2(G290), .ZN(n729) );
  XNOR2_X1 U805 ( .A(KEYINPUT100), .B(n729), .ZN(n730) );
  NOR2_X1 U806 ( .A1(n993), .A2(n730), .ZN(n732) );
  NOR2_X1 U807 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U808 ( .A1(n1004), .A2(n733), .ZN(n734) );
  XOR2_X1 U809 ( .A(n734), .B(KEYINPUT101), .Z(n735) );
  XNOR2_X1 U810 ( .A(KEYINPUT39), .B(n735), .ZN(n738) );
  INV_X1 U811 ( .A(n736), .ZN(n737) );
  NAND2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n740) );
  NAND2_X1 U813 ( .A1(n870), .A2(n739), .ZN(n998) );
  NAND2_X1 U814 ( .A1(n740), .A2(n998), .ZN(n742) );
  NAND2_X1 U815 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U816 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U817 ( .A(n745), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U818 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U819 ( .A(G132), .ZN(G219) );
  INV_X1 U820 ( .A(G82), .ZN(G220) );
  NAND2_X1 U821 ( .A1(G7), .A2(G661), .ZN(n746) );
  XNOR2_X1 U822 ( .A(n746), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U823 ( .A(G223), .ZN(n826) );
  NAND2_X1 U824 ( .A1(n826), .A2(G567), .ZN(n747) );
  XOR2_X1 U825 ( .A(KEYINPUT11), .B(n747), .Z(G234) );
  INV_X1 U826 ( .A(G860), .ZN(n753) );
  OR2_X1 U827 ( .A1(n915), .A2(n753), .ZN(G153) );
  INV_X1 U828 ( .A(G171), .ZN(G301) );
  NAND2_X1 U829 ( .A1(G868), .A2(G301), .ZN(n749) );
  INV_X1 U830 ( .A(G868), .ZN(n750) );
  NAND2_X1 U831 ( .A1(n929), .A2(n750), .ZN(n748) );
  NAND2_X1 U832 ( .A1(n749), .A2(n748), .ZN(G284) );
  INV_X1 U833 ( .A(n921), .ZN(G299) );
  NOR2_X1 U834 ( .A1(G286), .A2(n750), .ZN(n752) );
  NOR2_X1 U835 ( .A1(G868), .A2(G299), .ZN(n751) );
  NOR2_X1 U836 ( .A1(n752), .A2(n751), .ZN(G297) );
  NAND2_X1 U837 ( .A1(n753), .A2(G559), .ZN(n754) );
  NAND2_X1 U838 ( .A1(n754), .A2(n899), .ZN(n755) );
  XNOR2_X1 U839 ( .A(n755), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U840 ( .A1(G868), .A2(n915), .ZN(n758) );
  NAND2_X1 U841 ( .A1(G868), .A2(n899), .ZN(n756) );
  NOR2_X1 U842 ( .A1(G559), .A2(n756), .ZN(n757) );
  NOR2_X1 U843 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U844 ( .A(KEYINPUT68), .B(n759), .ZN(G282) );
  NAND2_X1 U845 ( .A1(G111), .A2(n881), .ZN(n761) );
  NAND2_X1 U846 ( .A1(G99), .A2(n884), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n767) );
  NAND2_X1 U848 ( .A1(n880), .A2(G123), .ZN(n762) );
  XNOR2_X1 U849 ( .A(n762), .B(KEYINPUT18), .ZN(n764) );
  NAND2_X1 U850 ( .A1(G135), .A2(n885), .ZN(n763) );
  NAND2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U852 ( .A(KEYINPUT69), .B(n765), .Z(n766) );
  NOR2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n992) );
  XNOR2_X1 U854 ( .A(n992), .B(G2096), .ZN(n769) );
  INV_X1 U855 ( .A(G2100), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n769), .A2(n768), .ZN(G156) );
  NAND2_X1 U857 ( .A1(G93), .A2(n770), .ZN(n773) );
  NAND2_X1 U858 ( .A1(G80), .A2(n771), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n779) );
  NAND2_X1 U860 ( .A1(G67), .A2(n774), .ZN(n777) );
  NAND2_X1 U861 ( .A1(G55), .A2(n775), .ZN(n776) );
  NAND2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U863 ( .A1(n779), .A2(n778), .ZN(n793) );
  XNOR2_X1 U864 ( .A(n915), .B(KEYINPUT70), .ZN(n781) );
  NAND2_X1 U865 ( .A1(n899), .A2(G559), .ZN(n780) );
  XNOR2_X1 U866 ( .A(n781), .B(n780), .ZN(n791) );
  NOR2_X1 U867 ( .A1(n791), .A2(G860), .ZN(n782) );
  XOR2_X1 U868 ( .A(KEYINPUT71), .B(n782), .Z(n783) );
  XNOR2_X1 U869 ( .A(n793), .B(n783), .ZN(G145) );
  XNOR2_X1 U870 ( .A(G166), .B(G305), .ZN(n784) );
  XNOR2_X1 U871 ( .A(n784), .B(G288), .ZN(n788) );
  XNOR2_X1 U872 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n786) );
  XNOR2_X1 U873 ( .A(G290), .B(KEYINPUT73), .ZN(n785) );
  XNOR2_X1 U874 ( .A(n786), .B(n785), .ZN(n787) );
  XOR2_X1 U875 ( .A(n788), .B(n787), .Z(n790) );
  XNOR2_X1 U876 ( .A(n921), .B(n793), .ZN(n789) );
  XNOR2_X1 U877 ( .A(n790), .B(n789), .ZN(n898) );
  XNOR2_X1 U878 ( .A(n791), .B(n898), .ZN(n792) );
  NAND2_X1 U879 ( .A1(n792), .A2(G868), .ZN(n795) );
  OR2_X1 U880 ( .A1(G868), .A2(n793), .ZN(n794) );
  NAND2_X1 U881 ( .A1(n795), .A2(n794), .ZN(G295) );
  NAND2_X1 U882 ( .A1(G2084), .A2(G2078), .ZN(n796) );
  XNOR2_X1 U883 ( .A(n796), .B(KEYINPUT20), .ZN(n797) );
  XNOR2_X1 U884 ( .A(n797), .B(KEYINPUT75), .ZN(n798) );
  NAND2_X1 U885 ( .A1(n798), .A2(G2090), .ZN(n799) );
  XNOR2_X1 U886 ( .A(n799), .B(KEYINPUT76), .ZN(n800) );
  XNOR2_X1 U887 ( .A(n800), .B(KEYINPUT21), .ZN(n801) );
  NAND2_X1 U888 ( .A1(n801), .A2(G2072), .ZN(n802) );
  XOR2_X1 U889 ( .A(KEYINPUT77), .B(n802), .Z(G158) );
  XOR2_X1 U890 ( .A(KEYINPUT66), .B(G57), .Z(G237) );
  XNOR2_X1 U891 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U892 ( .A1(G108), .A2(G120), .ZN(n803) );
  NOR2_X1 U893 ( .A1(G237), .A2(n803), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G69), .A2(n804), .ZN(n830) );
  NAND2_X1 U895 ( .A1(n830), .A2(G567), .ZN(n812) );
  NOR2_X1 U896 ( .A1(G220), .A2(G219), .ZN(n807) );
  XOR2_X1 U897 ( .A(KEYINPUT22), .B(KEYINPUT79), .Z(n805) );
  XNOR2_X1 U898 ( .A(KEYINPUT78), .B(n805), .ZN(n806) );
  XNOR2_X1 U899 ( .A(n807), .B(n806), .ZN(n808) );
  NAND2_X1 U900 ( .A1(G96), .A2(n808), .ZN(n809) );
  NOR2_X1 U901 ( .A1(G218), .A2(n809), .ZN(n810) );
  XOR2_X1 U902 ( .A(KEYINPUT80), .B(n810), .Z(n831) );
  NAND2_X1 U903 ( .A1(n831), .A2(G2106), .ZN(n811) );
  NAND2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n832) );
  NAND2_X1 U905 ( .A1(G661), .A2(G483), .ZN(n813) );
  XOR2_X1 U906 ( .A(KEYINPUT81), .B(n813), .Z(n814) );
  NOR2_X1 U907 ( .A1(n832), .A2(n814), .ZN(n829) );
  NAND2_X1 U908 ( .A1(n829), .A2(G36), .ZN(G176) );
  XNOR2_X1 U909 ( .A(G2443), .B(G2435), .ZN(n824) );
  XOR2_X1 U910 ( .A(G2454), .B(G2430), .Z(n816) );
  XNOR2_X1 U911 ( .A(G2446), .B(KEYINPUT103), .ZN(n815) );
  XNOR2_X1 U912 ( .A(n816), .B(n815), .ZN(n820) );
  XOR2_X1 U913 ( .A(G2451), .B(G2427), .Z(n818) );
  XNOR2_X1 U914 ( .A(G1341), .B(G1348), .ZN(n817) );
  XNOR2_X1 U915 ( .A(n818), .B(n817), .ZN(n819) );
  XOR2_X1 U916 ( .A(n820), .B(n819), .Z(n822) );
  XNOR2_X1 U917 ( .A(G2438), .B(KEYINPUT102), .ZN(n821) );
  XNOR2_X1 U918 ( .A(n822), .B(n821), .ZN(n823) );
  XNOR2_X1 U919 ( .A(n824), .B(n823), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n825), .A2(G14), .ZN(n906) );
  XOR2_X1 U921 ( .A(KEYINPUT104), .B(n906), .Z(G401) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U924 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U926 ( .A1(n829), .A2(n828), .ZN(G188) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G108), .ZN(G238) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  INV_X1 U931 ( .A(G69), .ZN(G235) );
  NOR2_X1 U932 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  INV_X1 U934 ( .A(n832), .ZN(G319) );
  XOR2_X1 U935 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n834) );
  XNOR2_X1 U936 ( .A(G2678), .B(KEYINPUT43), .ZN(n833) );
  XNOR2_X1 U937 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U938 ( .A(KEYINPUT42), .B(G2090), .Z(n836) );
  XNOR2_X1 U939 ( .A(G2067), .B(G2072), .ZN(n835) );
  XNOR2_X1 U940 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U941 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U942 ( .A(G2096), .B(G2100), .ZN(n839) );
  XNOR2_X1 U943 ( .A(n840), .B(n839), .ZN(n842) );
  XOR2_X1 U944 ( .A(G2084), .B(G2078), .Z(n841) );
  XNOR2_X1 U945 ( .A(n842), .B(n841), .ZN(G227) );
  XOR2_X1 U946 ( .A(G1976), .B(G1981), .Z(n844) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1971), .ZN(n843) );
  XNOR2_X1 U948 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U949 ( .A(G1961), .B(G1966), .Z(n846) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1991), .ZN(n845) );
  XNOR2_X1 U951 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U952 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U953 ( .A(KEYINPUT107), .B(G2474), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n850), .B(n849), .ZN(n852) );
  XOR2_X1 U955 ( .A(G1956), .B(KEYINPUT41), .Z(n851) );
  XNOR2_X1 U956 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G112), .A2(n881), .ZN(n854) );
  NAND2_X1 U958 ( .A1(G100), .A2(n884), .ZN(n853) );
  NAND2_X1 U959 ( .A1(n854), .A2(n853), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G136), .A2(n885), .ZN(n855) );
  XNOR2_X1 U961 ( .A(n855), .B(KEYINPUT108), .ZN(n858) );
  NAND2_X1 U962 ( .A1(G124), .A2(n880), .ZN(n856) );
  XNOR2_X1 U963 ( .A(n856), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U964 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U965 ( .A1(n860), .A2(n859), .ZN(G162) );
  NAND2_X1 U966 ( .A1(G103), .A2(n884), .ZN(n862) );
  NAND2_X1 U967 ( .A1(G139), .A2(n885), .ZN(n861) );
  NAND2_X1 U968 ( .A1(n862), .A2(n861), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n881), .A2(G115), .ZN(n863) );
  XNOR2_X1 U970 ( .A(n863), .B(KEYINPUT110), .ZN(n865) );
  NAND2_X1 U971 ( .A1(G127), .A2(n880), .ZN(n864) );
  NAND2_X1 U972 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U973 ( .A(KEYINPUT47), .B(n866), .Z(n867) );
  NOR2_X1 U974 ( .A1(n868), .A2(n867), .ZN(n999) );
  XOR2_X1 U975 ( .A(n999), .B(n992), .Z(n869) );
  XNOR2_X1 U976 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U977 ( .A(G164), .B(G162), .Z(n871) );
  XNOR2_X1 U978 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U979 ( .A(n874), .B(n873), .Z(n879) );
  XOR2_X1 U980 ( .A(KEYINPUT113), .B(KEYINPUT111), .Z(n876) );
  XNOR2_X1 U981 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n875) );
  XNOR2_X1 U982 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U983 ( .A(KEYINPUT112), .B(n877), .ZN(n878) );
  XNOR2_X1 U984 ( .A(n879), .B(n878), .ZN(n896) );
  NAND2_X1 U985 ( .A1(G130), .A2(n880), .ZN(n883) );
  NAND2_X1 U986 ( .A1(G118), .A2(n881), .ZN(n882) );
  NAND2_X1 U987 ( .A1(n883), .A2(n882), .ZN(n891) );
  NAND2_X1 U988 ( .A1(G106), .A2(n884), .ZN(n887) );
  NAND2_X1 U989 ( .A1(G142), .A2(n885), .ZN(n886) );
  NAND2_X1 U990 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U991 ( .A(KEYINPUT45), .B(n888), .ZN(n889) );
  XNOR2_X1 U992 ( .A(KEYINPUT109), .B(n889), .ZN(n890) );
  NOR2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U994 ( .A(G160), .B(n892), .ZN(n894) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U997 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U998 ( .A(G286), .B(n898), .ZN(n903) );
  XOR2_X1 U999 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n901) );
  XNOR2_X1 U1000 ( .A(G171), .B(n899), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1003 ( .A(n904), .B(n915), .Z(n905) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n905), .ZN(G397) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n906), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n911) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n910) );
  NAND2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1012 ( .A(G16), .B(KEYINPUT56), .Z(n937) );
  XNOR2_X1 U1013 ( .A(G1966), .B(G168), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(n914), .B(KEYINPUT57), .ZN(n928) );
  XNOR2_X1 U1016 ( .A(n915), .B(G1341), .ZN(n926) );
  AND2_X1 U1017 ( .A1(G303), .A2(G1971), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1020 ( .A(KEYINPUT120), .B(n920), .Z(n923) );
  XOR2_X1 U1021 ( .A(n921), .B(G1956), .Z(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(KEYINPUT121), .B(n924), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n935) );
  XNOR2_X1 U1026 ( .A(G301), .B(G1961), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(n929), .B(G1348), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n990) );
  XNOR2_X1 U1032 ( .A(G1966), .B(G21), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(G1961), .B(G5), .ZN(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n953) );
  XNOR2_X1 U1035 ( .A(KEYINPUT60), .B(KEYINPUT125), .ZN(n951) );
  XNOR2_X1 U1036 ( .A(KEYINPUT59), .B(G4), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(n940), .B(KEYINPUT124), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(G1348), .B(n941), .ZN(n949) );
  XNOR2_X1 U1039 ( .A(G1956), .B(G20), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(G1981), .B(G6), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(n942), .B(KEYINPUT122), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(G19), .B(G1341), .ZN(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(KEYINPUT123), .B(n945), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(n951), .B(n950), .ZN(n952) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n960) );
  XNOR2_X1 U1049 ( .A(G1971), .B(G22), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G23), .B(G1976), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n957) );
  XOR2_X1 U1052 ( .A(G1986), .B(G24), .Z(n956) );
  NAND2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(KEYINPUT58), .B(n958), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1056 ( .A(KEYINPUT61), .B(n961), .Z(n962) );
  NOR2_X1 U1057 ( .A1(G16), .A2(n962), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(n963), .B(KEYINPUT126), .ZN(n987) );
  XOR2_X1 U1059 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n984) );
  XNOR2_X1 U1060 ( .A(G2090), .B(G35), .ZN(n978) );
  XNOR2_X1 U1061 ( .A(G2067), .B(G26), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(G32), .B(G1996), .ZN(n964) );
  NOR2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(n966), .B(G27), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(G33), .B(G2072), .ZN(n967) );
  NOR2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(KEYINPUT117), .B(n971), .ZN(n972) );
  NAND2_X1 U1069 ( .A1(n972), .A2(G28), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(G25), .B(n973), .ZN(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1072 ( .A(KEYINPUT53), .B(n976), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n982) );
  XOR2_X1 U1074 ( .A(KEYINPUT118), .B(G34), .Z(n980) );
  XNOR2_X1 U1075 ( .A(G2084), .B(KEYINPUT54), .ZN(n979) );
  XNOR2_X1 U1076 ( .A(n980), .B(n979), .ZN(n981) );
  NAND2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(n984), .B(n983), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(G29), .A2(n985), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(G11), .A2(n988), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(n991), .B(KEYINPUT127), .ZN(n1017) );
  INV_X1 U1084 ( .A(G29), .ZN(n1015) );
  XNOR2_X1 U1085 ( .A(G160), .B(G2084), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1088 ( .A(KEYINPUT116), .B(n996), .Z(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1011) );
  XOR2_X1 U1090 ( .A(G2072), .B(n999), .Z(n1001) );
  XOR2_X1 U1091 ( .A(G164), .B(G2078), .Z(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1093 ( .A(KEYINPUT50), .B(n1002), .Z(n1007) );
  XOR2_X1 U1094 ( .A(G2090), .B(G162), .Z(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(KEYINPUT51), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1100 ( .A(KEYINPUT52), .B(n1012), .Z(n1013) );
  NOR2_X1 U1101 ( .A1(KEYINPUT55), .A2(n1013), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1018), .ZN(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

