//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT31), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT68), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT64), .A3(G116), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G119), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(G119), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n191), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT2), .B(G113), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT2), .B(G113), .Z(new_n199));
  OAI211_X1 g013(.A(new_n199), .B(new_n191), .C1(new_n195), .C2(new_n194), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(KEYINPUT1), .A3(G146), .ZN(new_n209));
  XNOR2_X1  g023(.A(G143), .B(G146), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n208), .B(new_n209), .C1(G128), .C2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G137), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT11), .A3(G134), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(G137), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n214), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n218), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n213), .A2(G137), .ZN(new_n221));
  OAI21_X1  g035(.A(G131), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n211), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n214), .A2(new_n218), .A3(new_n216), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G131), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n219), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n205), .A2(new_n207), .A3(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT0), .B(G128), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n210), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n226), .A2(KEYINPUT65), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT65), .B1(new_n226), .B2(new_n231), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n223), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT30), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n226), .A2(new_n231), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT30), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n236), .A2(new_n223), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n201), .B1(new_n235), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n223), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n226), .A2(KEYINPUT65), .A3(new_n231), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n241), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n201), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(G101), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G237), .ZN(new_n249));
  INV_X1    g063(.A(G953), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n250), .A3(G210), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT67), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n251), .B(KEYINPUT67), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(new_n254), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n248), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n254), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n253), .A2(new_n255), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(new_n247), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n246), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n189), .B1(new_n240), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n263), .B1(new_n245), .B2(new_n201), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n238), .B1(new_n234), .B2(KEYINPUT30), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n267), .B(KEYINPUT68), .C1(new_n268), .C2(new_n201), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n188), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n236), .A2(new_n223), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n201), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OR2_X1    g088(.A1(new_n271), .A2(new_n201), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n274), .B(new_n275), .C1(new_n246), .C2(new_n273), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(new_n264), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n239), .B1(new_n245), .B2(new_n237), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n198), .A2(new_n200), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(new_n188), .A3(new_n267), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n270), .A2(new_n278), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n285));
  NOR2_X1   g099(.A1(G472), .A2(G902), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT68), .B1(new_n281), .B2(new_n267), .ZN(new_n289));
  INV_X1    g103(.A(new_n269), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT31), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n278), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n282), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT69), .B1(new_n293), .B2(new_n286), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n187), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n286), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(new_n187), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n281), .A2(new_n246), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n263), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT29), .B1(new_n277), .B2(new_n264), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G902), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n234), .A2(new_n280), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n246), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT28), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n308), .A2(KEYINPUT29), .A3(new_n264), .A4(new_n274), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(KEYINPUT70), .ZN(new_n310));
  OAI21_X1  g124(.A(G472), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n295), .A2(new_n298), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n313), .A2(G125), .A3(G140), .ZN(new_n314));
  AOI21_X1  g128(.A(G140), .B1(new_n313), .B2(G125), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT16), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT73), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT16), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(G125), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n319), .B1(new_n321), .B2(KEYINPUT72), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n313), .A2(G125), .A3(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT16), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n317), .A2(G146), .A3(new_n320), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT74), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n325), .B1(new_n324), .B2(KEYINPUT16), .ZN(new_n329));
  AOI211_X1 g143(.A(KEYINPUT73), .B(new_n318), .C1(new_n322), .C2(new_n323), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n331), .A2(new_n332), .A3(G146), .A4(new_n320), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n319), .A2(G125), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n321), .A2(G140), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n335), .A2(new_n336), .A3(new_n204), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n202), .A2(G119), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n190), .A2(G128), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(G110), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n339), .A2(new_n342), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT24), .B(G110), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n334), .B(new_n338), .C1(new_n345), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n344), .A2(G110), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n350), .B(KEYINPUT71), .Z(new_n351));
  NOR2_X1   g165(.A1(new_n346), .A2(new_n347), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(G146), .B1(new_n331), .B2(new_n320), .ZN(new_n354));
  INV_X1    g168(.A(new_n327), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n351), .B(new_n353), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n250), .A2(G221), .A3(G234), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT22), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(G137), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(KEYINPUT75), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT76), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n364));
  AOI211_X1 g178(.A(new_n364), .B(new_n361), .C1(new_n349), .C2(new_n356), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n349), .A2(new_n356), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n360), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G217), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(G234), .B2(new_n304), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(G902), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n364), .B1(new_n367), .B2(new_n361), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n357), .A2(KEYINPUT76), .A3(new_n362), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n375), .A2(new_n304), .A3(new_n368), .A4(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n366), .A2(KEYINPUT25), .A3(new_n304), .A4(new_n368), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n374), .B1(new_n381), .B2(new_n371), .ZN(new_n382));
  OAI21_X1  g196(.A(G214), .B1(G237), .B2(G902), .ZN(new_n383));
  NAND2_X1  g197(.A1(G234), .A2(G237), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n384), .A2(G952), .A3(new_n250), .ZN(new_n385));
  XOR2_X1   g199(.A(KEYINPUT21), .B(G898), .Z(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT94), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n384), .A2(G902), .A3(G953), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n230), .A2(G125), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT85), .ZN(new_n395));
  INV_X1    g209(.A(G224), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(G953), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT7), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n211), .A2(G125), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n394), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n403));
  INV_X1    g217(.A(G104), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT3), .B1(new_n404), .B2(G107), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT3), .ZN(new_n406));
  INV_X1    g220(.A(G107), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(G104), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(G107), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G101), .ZN(new_n411));
  INV_X1    g225(.A(G101), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n405), .A2(new_n408), .A3(new_n412), .A4(new_n409), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(KEYINPUT4), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n410), .A2(new_n415), .A3(G101), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n403), .B1(new_n417), .B2(new_n201), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT5), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n195), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g234(.A(G113), .B(new_n420), .C1(new_n196), .C2(new_n419), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n407), .A2(G104), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n404), .A2(G107), .ZN(new_n423));
  OAI21_X1  g237(.A(G101), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n413), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n426), .A3(new_n200), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n280), .A2(new_n414), .A3(KEYINPUT82), .A4(new_n416), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n418), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  XOR2_X1   g243(.A(G110), .B(G122), .Z(new_n430));
  OR2_X1    g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n421), .A2(new_n200), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n425), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n427), .ZN(new_n434));
  XOR2_X1   g248(.A(new_n430), .B(KEYINPUT8), .Z(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n394), .A2(new_n401), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n395), .A3(new_n399), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n402), .A2(new_n431), .A3(new_n436), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(KEYINPUT83), .A2(KEYINPUT6), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n429), .A2(new_n430), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n441), .B1(new_n429), .B2(new_n430), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n429), .A2(new_n430), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n437), .B(new_n398), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n304), .B(new_n439), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G210), .B1(G237), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n429), .A2(new_n430), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n440), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n429), .A2(new_n430), .A3(new_n441), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n431), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n446), .ZN(new_n455));
  AOI21_X1  g269(.A(G902), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n448), .B1(new_n456), .B2(new_n439), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n383), .B(new_n391), .C1(new_n450), .C2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT80), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n414), .A2(new_n231), .A3(new_n416), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT77), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n426), .A2(new_n211), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT10), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n226), .B(KEYINPUT78), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT79), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT12), .B1(new_n226), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n211), .B(new_n425), .ZN(new_n468));
  INV_X1    g282(.A(new_n226), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n468), .A2(new_n469), .A3(new_n467), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n459), .B1(new_n465), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(G110), .B(G140), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n250), .A2(G227), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n479), .B(KEYINPUT80), .C1(new_n472), .C2(new_n471), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n474), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n469), .B1(new_n461), .B2(new_n463), .ZN(new_n482));
  OR3_X1    g296(.A1(new_n465), .A2(new_n482), .A3(new_n478), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(G469), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n478), .B1(new_n465), .B2(new_n482), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT81), .B1(new_n471), .B2(new_n472), .ZN(new_n486));
  OR2_X1    g300(.A1(new_n426), .A2(new_n211), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n469), .B1(new_n487), .B2(new_n462), .ZN(new_n488));
  INV_X1    g302(.A(new_n467), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT81), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n470), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n486), .A2(new_n477), .A3(new_n492), .A4(new_n479), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G469), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n495), .A3(new_n304), .ZN(new_n496));
  NAND2_X1  g310(.A1(G469), .A2(G902), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n484), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G221), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT9), .B(G234), .Z(new_n500));
  AOI21_X1  g314(.A(new_n499), .B1(new_n500), .B2(new_n304), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G113), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(new_n404), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n249), .A2(new_n250), .A3(G214), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT86), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G143), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n206), .A2(KEYINPUT86), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(G237), .A2(G953), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n512), .A2(KEYINPUT86), .A3(new_n206), .A4(G214), .ZN(new_n513));
  AOI21_X1  g327(.A(G131), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n511), .A2(G131), .A3(new_n513), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT88), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT88), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n511), .A2(new_n517), .A3(G131), .A4(new_n513), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n514), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT19), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n335), .A2(new_n336), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT89), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT89), .A4(new_n521), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n524), .B(new_n525), .C1(new_n521), .C2(new_n324), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(G146), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n334), .A2(new_n520), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(KEYINPUT87), .A2(KEYINPUT18), .ZN(new_n530));
  INV_X1    g344(.A(new_n514), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n530), .B1(new_n531), .B2(new_n515), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n511), .A2(new_n513), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n533), .A2(new_n530), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n324), .A2(new_n204), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(new_n337), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n529), .A2(KEYINPUT90), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT90), .B1(new_n529), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n506), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G475), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n354), .A2(new_n355), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n516), .A2(KEYINPUT17), .A3(new_n518), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n543), .B(new_n544), .C1(KEYINPUT17), .C2(new_n520), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n506), .B1(new_n545), .B2(new_n538), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n541), .A2(new_n542), .A3(new_n304), .A4(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT20), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT90), .ZN(new_n551));
  AOI211_X1 g365(.A(new_n527), .B(new_n519), .C1(new_n328), .C2(new_n333), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n551), .B1(new_n552), .B2(new_n537), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n529), .A2(KEYINPUT90), .A3(new_n538), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n546), .B1(new_n555), .B2(new_n506), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n556), .A2(KEYINPUT20), .A3(new_n542), .A4(new_n304), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n500), .A2(G217), .A3(new_n250), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n558), .B(KEYINPUT93), .Z(new_n559));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n560), .B1(new_n202), .B2(G143), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n206), .A2(KEYINPUT92), .A3(G128), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(G128), .B2(new_n206), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n564), .A2(G134), .ZN(new_n565));
  XOR2_X1   g379(.A(G116), .B(G122), .Z(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(G107), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT13), .B1(new_n561), .B2(new_n562), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n561), .A2(KEYINPUT13), .A3(new_n562), .ZN(new_n569));
  AOI211_X1 g383(.A(new_n568), .B(new_n569), .C1(new_n202), .C2(G143), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n565), .B(new_n567), .C1(new_n570), .C2(new_n213), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n564), .B(G134), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n193), .A2(G122), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n407), .B1(new_n573), .B2(KEYINPUT14), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n574), .B(new_n566), .Z(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n559), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n571), .A2(new_n576), .A3(new_n559), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n304), .ZN(new_n581));
  INV_X1    g395(.A(G478), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(KEYINPUT15), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n581), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n545), .A2(new_n538), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n506), .A2(KEYINPUT91), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n304), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n586), .A2(new_n587), .ZN(new_n590));
  OAI21_X1  g404(.A(G475), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n550), .A2(new_n557), .A3(new_n585), .A4(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n458), .A2(new_n503), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n312), .A2(new_n382), .A3(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT95), .B(G101), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G3));
  OAI21_X1  g410(.A(new_n285), .B1(new_n284), .B2(new_n287), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n293), .A2(KEYINPUT69), .A3(new_n286), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(G472), .B1(new_n284), .B2(G902), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n382), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n602), .A2(new_n603), .A3(new_n503), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n550), .A2(new_n557), .A3(new_n591), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n580), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n578), .A2(KEYINPUT33), .A3(new_n579), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n607), .A2(G478), .A3(new_n304), .A4(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n581), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n609), .B1(G478), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n458), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n604), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT34), .B(G104), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n617));
  INV_X1    g431(.A(new_n383), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n447), .A2(new_n449), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n456), .A2(new_n448), .A3(new_n439), .ZN(new_n620));
  AOI211_X1 g434(.A(new_n618), .B(new_n390), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n581), .B(new_n583), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n550), .A2(new_n557), .A3(new_n622), .A4(new_n591), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n617), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n458), .A2(new_n623), .A3(KEYINPUT96), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n604), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  NOR2_X1   g444(.A1(new_n362), .A2(KEYINPUT36), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(new_n357), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n381), .A2(new_n371), .B1(new_n372), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n601), .A2(new_n593), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT37), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n636), .B(G110), .Z(G12));
  AOI21_X1  g451(.A(new_n297), .B1(new_n599), .B2(new_n187), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n633), .B1(new_n638), .B2(new_n311), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n550), .A2(new_n557), .A3(new_n591), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT97), .ZN(new_n642));
  INV_X1    g456(.A(new_n389), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n642), .B1(new_n643), .B2(G900), .ZN(new_n644));
  INV_X1    g458(.A(new_n385), .ZN(new_n645));
  INV_X1    g459(.A(G900), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n389), .A2(KEYINPUT97), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n641), .A2(KEYINPUT98), .A3(new_n622), .A4(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT98), .ZN(new_n650));
  INV_X1    g464(.A(new_n648), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n650), .B1(new_n623), .B2(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n498), .A2(new_n502), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n649), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n639), .A2(new_n640), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT99), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  XNOR2_X1  g471(.A(new_n648), .B(KEYINPUT101), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT39), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n660), .B(KEYINPUT40), .Z(new_n661));
  NAND2_X1  g475(.A1(new_n619), .A2(new_n620), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT38), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n307), .A2(new_n263), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT100), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n266), .A2(new_n269), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n304), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(G472), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n638), .A2(new_n669), .ZN(new_n670));
  NOR4_X1   g484(.A1(new_n634), .A2(new_n618), .A3(new_n585), .A4(new_n641), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n661), .A2(new_n663), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G143), .ZN(G45));
  NAND3_X1  g487(.A1(new_n605), .A2(new_n611), .A3(new_n648), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n639), .A2(new_n653), .A3(new_n640), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT102), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n204), .ZN(G48));
  NAND2_X1  g492(.A1(new_n494), .A2(new_n304), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G469), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n496), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n501), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n312), .A2(new_n382), .A3(new_n613), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT41), .B(G113), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G15));
  NAND4_X1  g499(.A1(new_n627), .A2(new_n312), .A3(new_n382), .A4(new_n682), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G116), .ZN(G18));
  NOR4_X1   g501(.A1(new_n592), .A2(new_n681), .A3(new_n501), .A4(new_n390), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n312), .A2(new_n688), .A3(new_n640), .A4(new_n634), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  NAND2_X1  g504(.A1(new_n308), .A2(new_n274), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n264), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n692), .B2(new_n691), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n270), .A2(new_n283), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n286), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n382), .A2(new_n682), .A3(new_n600), .A4(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n699), .A2(new_n621), .A3(new_n622), .A4(new_n605), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G122), .ZN(G24));
  NAND2_X1  g515(.A1(new_n682), .A2(new_n640), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n697), .A2(new_n600), .ZN(new_n703));
  NOR4_X1   g517(.A1(new_n702), .A2(new_n703), .A3(new_n633), .A4(new_n674), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n321), .ZN(G27));
  NAND3_X1  g519(.A1(new_n296), .A2(KEYINPUT104), .A3(new_n187), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n287), .B1(new_n695), .B2(new_n292), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n707), .B1(new_n708), .B2(KEYINPUT32), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(KEYINPUT32), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n311), .B(new_n706), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n619), .A2(new_n383), .A3(new_n620), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n503), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n711), .A2(new_n382), .A3(new_n713), .A4(new_n675), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT42), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n674), .A2(KEYINPUT42), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n312), .A2(new_n382), .A3(new_n713), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n217), .ZN(G33));
  AND2_X1   g533(.A1(new_n649), .A2(new_n652), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n720), .A2(new_n312), .A3(new_n382), .A4(new_n713), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G134), .ZN(G36));
  INV_X1    g536(.A(new_n611), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n605), .A2(new_n723), .A3(KEYINPUT43), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n605), .B(KEYINPUT105), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n611), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n724), .B1(new_n726), .B2(KEYINPUT43), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n602), .A3(new_n634), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n712), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n728), .A2(new_n729), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n481), .A2(new_n483), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT45), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(G469), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(KEYINPUT46), .A3(new_n497), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n738), .B(G469), .C1(new_n735), .C2(G902), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n737), .A2(new_n496), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n502), .A3(new_n659), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n733), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G137), .ZN(G39));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n502), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n740), .A2(new_n746), .A3(new_n502), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n748), .A2(new_n674), .A3(new_n712), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(new_n638), .A3(new_n311), .A4(new_n603), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G140), .ZN(G42));
  INV_X1    g565(.A(new_n704), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n605), .A2(new_n662), .A3(new_n383), .A4(new_n622), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n633), .A2(new_n653), .A3(new_n648), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n633), .A2(new_n653), .A3(KEYINPUT110), .A4(new_n648), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n670), .A3(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n676), .A2(new_n655), .A3(new_n752), .A4(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n312), .A2(new_n640), .A3(new_n634), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n704), .B1(new_n762), .B2(new_n654), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n763), .A2(KEYINPUT52), .A3(new_n676), .A4(new_n758), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NOR4_X1   g579(.A1(new_n503), .A2(new_n592), .A3(new_n712), .A4(new_n651), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n312), .A2(new_n634), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT108), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n703), .A2(new_n633), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n675), .A3(new_n713), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n312), .A2(KEYINPUT108), .A3(new_n766), .A4(new_n634), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n769), .A2(new_n721), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT109), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n721), .A2(new_n771), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n769), .A4(new_n772), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n623), .A2(KEYINPUT107), .ZN(new_n779));
  MUX2_X1   g593(.A(KEYINPUT107), .B(new_n779), .S(new_n612), .Z(new_n780));
  NAND3_X1  g594(.A1(new_n604), .A2(new_n621), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n594), .A3(new_n635), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n765), .A2(new_n778), .A3(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n686), .A2(new_n700), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n312), .A2(new_n382), .A3(new_n713), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n786), .A2(new_n716), .B1(new_n714), .B2(KEYINPUT42), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n683), .A2(new_n689), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n785), .A2(new_n787), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n686), .A2(new_n683), .A3(new_n700), .A4(new_n689), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT113), .B1(new_n791), .B2(new_n718), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(new_n792), .A3(KEYINPUT53), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT114), .B1(new_n784), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n791), .A2(new_n718), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n765), .A2(new_n778), .A3(new_n795), .A4(new_n783), .ZN(new_n796));
  XOR2_X1   g610(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n790), .A2(new_n792), .A3(KEYINPUT53), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n782), .B1(new_n774), .B2(new_n777), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n800), .A2(new_n801), .A3(new_n765), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n794), .A2(new_n799), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  OR3_X1    g620(.A1(new_n796), .A2(KEYINPUT112), .A3(new_n798), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n796), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT112), .B1(new_n796), .B2(new_n798), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n806), .B1(KEYINPUT54), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n813));
  NOR4_X1   g627(.A1(new_n712), .A2(new_n681), .A3(new_n501), .A4(new_n645), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n727), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n770), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n670), .A2(new_n603), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n723), .A3(new_n814), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n727), .A2(new_n385), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n820), .A2(new_n383), .A3(new_n663), .A4(new_n698), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(KEYINPUT50), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(KEYINPUT50), .ZN(new_n823));
  OAI221_X1 g637(.A(new_n817), .B1(new_n605), .B2(new_n819), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  OR4_X1    g638(.A1(new_n603), .A2(new_n820), .A3(new_n703), .A4(new_n712), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n748), .B1(new_n502), .B2(new_n681), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n813), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n711), .A2(new_n382), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n816), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT48), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n250), .A2(G952), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n820), .A2(new_n698), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n833), .B1(new_n834), .B2(new_n640), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n829), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n827), .A2(KEYINPUT116), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n827), .A2(KEYINPUT116), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n826), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT51), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n824), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n818), .A2(new_n814), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n812), .B(new_n842), .C1(new_n612), .C2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(G952), .B2(G953), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n726), .A2(new_n501), .A3(new_n663), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n681), .A2(KEYINPUT49), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT106), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n618), .B1(new_n681), .B2(KEYINPUT49), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n846), .A2(new_n818), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n845), .A2(new_n850), .ZN(G75));
  INV_X1    g665(.A(KEYINPUT56), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n794), .A2(new_n799), .A3(new_n803), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(G902), .ZN(new_n854));
  INV_X1    g668(.A(G210), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n454), .B(new_n455), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT55), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n856), .A2(KEYINPUT117), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT117), .B1(new_n856), .B2(new_n858), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n854), .A2(KEYINPUT118), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n853), .A2(new_n862), .A3(G902), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n448), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n865));
  OAI22_X1  g679(.A1(new_n859), .A2(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n250), .A2(G952), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT119), .Z(new_n868));
  NOR2_X1   g682(.A1(new_n866), .A2(new_n868), .ZN(G51));
  INV_X1    g683(.A(new_n867), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n736), .B1(new_n861), .B2(new_n863), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n494), .B(KEYINPUT120), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n853), .A2(KEYINPUT54), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n805), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n497), .B(KEYINPUT57), .Z(new_n875));
  AOI21_X1  g689(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n870), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(KEYINPUT121), .B(new_n870), .C1(new_n871), .C2(new_n876), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(G54));
  NAND2_X1  g695(.A1(new_n861), .A2(new_n863), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n882), .A2(KEYINPUT58), .A3(G475), .ZN(new_n883));
  INV_X1    g697(.A(new_n556), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n882), .A2(KEYINPUT58), .A3(G475), .A4(new_n556), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n885), .A2(new_n870), .A3(new_n886), .ZN(G60));
  NAND2_X1  g701(.A1(new_n607), .A2(new_n608), .ZN(new_n888));
  NAND2_X1  g702(.A1(G478), .A2(G902), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT59), .Z(new_n890));
  OAI21_X1  g704(.A(new_n888), .B1(new_n812), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n868), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n888), .B1(new_n873), .B2(new_n805), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n894));
  INV_X1    g708(.A(new_n890), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n894), .B1(new_n893), .B2(new_n895), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n891), .B(new_n892), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(G63));
  NAND2_X1  g713(.A1(G217), .A2(G902), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT123), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT60), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n853), .A2(new_n632), .A3(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n853), .A2(new_n902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n369), .B(KEYINPUT124), .Z(new_n905));
  OAI211_X1 g719(.A(new_n892), .B(new_n903), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g721(.A(G953), .B1(new_n388), .B2(new_n396), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n782), .A2(new_n791), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(G953), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n445), .B1(G898), .B2(new_n250), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(G69));
  XNOR2_X1  g726(.A(new_n279), .B(new_n526), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(G227), .A3(G953), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n763), .A2(new_n676), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n672), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT62), .Z(new_n918));
  NAND3_X1  g732(.A1(new_n786), .A2(new_n659), .A3(new_n780), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n918), .A2(new_n742), .A3(new_n750), .A4(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n250), .B1(new_n920), .B2(new_n914), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n750), .A2(new_n787), .ZN(new_n922));
  INV_X1    g736(.A(new_n753), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n830), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n741), .B1(new_n733), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n916), .A2(new_n721), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n913), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n915), .B1(new_n921), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(G227), .B1(new_n914), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g747(.A(G953), .B1(new_n933), .B2(new_n646), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(G72));
  NAND2_X1  g749(.A1(G472), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT63), .Z(new_n937));
  INV_X1    g751(.A(new_n909), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n920), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n264), .A3(new_n300), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n301), .A2(new_n666), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n811), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n926), .A2(new_n909), .A3(new_n928), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n937), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n299), .A2(new_n263), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT126), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n870), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n949), .A2(KEYINPUT127), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(KEYINPUT127), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n943), .B1(new_n950), .B2(new_n951), .ZN(G57));
endmodule


