

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U548 ( .A(n590), .ZN(n875) );
  NOR2_X1 U549 ( .A1(G2084), .A2(n717), .ZN(n703) );
  INV_X1 U550 ( .A(KEYINPUT17), .ZN(n512) );
  XNOR2_X1 U551 ( .A(n512), .B(KEYINPUT66), .ZN(n513) );
  XNOR2_X1 U552 ( .A(n514), .B(n513), .ZN(n589) );
  NAND2_X1 U553 ( .A1(n811), .A2(n801), .ZN(n802) );
  OR2_X1 U554 ( .A1(n803), .A2(n802), .ZN(n816) );
  NOR2_X1 U555 ( .A1(n524), .A2(n523), .ZN(G160) );
  NOR2_X1 U556 ( .A1(G2105), .A2(G2104), .ZN(n514) );
  NAND2_X1 U557 ( .A1(G137), .A2(n589), .ZN(n515) );
  XOR2_X1 U558 ( .A(KEYINPUT67), .B(n515), .Z(n519) );
  INV_X1 U559 ( .A(G2105), .ZN(n520) );
  AND2_X2 U560 ( .A1(n520), .A2(G2104), .ZN(n874) );
  NAND2_X1 U561 ( .A1(G101), .A2(n874), .ZN(n516) );
  XNOR2_X1 U562 ( .A(n516), .B(KEYINPUT23), .ZN(n517) );
  XNOR2_X1 U563 ( .A(KEYINPUT65), .B(n517), .ZN(n518) );
  NAND2_X1 U564 ( .A1(n519), .A2(n518), .ZN(n524) );
  NOR2_X1 U565 ( .A1(G2104), .A2(n520), .ZN(n869) );
  NAND2_X1 U566 ( .A1(G125), .A2(n869), .ZN(n522) );
  AND2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n870) );
  NAND2_X1 U568 ( .A1(G113), .A2(n870), .ZN(n521) );
  NAND2_X1 U569 ( .A1(n522), .A2(n521), .ZN(n523) );
  INV_X1 U570 ( .A(G651), .ZN(n530) );
  NOR2_X1 U571 ( .A1(G543), .A2(n530), .ZN(n526) );
  XNOR2_X1 U572 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n525) );
  XNOR2_X1 U573 ( .A(n526), .B(n525), .ZN(n631) );
  NAND2_X1 U574 ( .A1(n631), .A2(G64), .ZN(n529) );
  XOR2_X1 U575 ( .A(G543), .B(KEYINPUT0), .Z(n617) );
  NOR2_X1 U576 ( .A1(G651), .A2(n617), .ZN(n527) );
  XNOR2_X1 U577 ( .A(KEYINPUT64), .B(n527), .ZN(n639) );
  NAND2_X1 U578 ( .A1(G52), .A2(n639), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n536) );
  NOR2_X1 U580 ( .A1(G651), .A2(G543), .ZN(n632) );
  NAND2_X1 U581 ( .A1(G90), .A2(n632), .ZN(n532) );
  NOR2_X1 U582 ( .A1(n617), .A2(n530), .ZN(n635) );
  NAND2_X1 U583 ( .A1(G77), .A2(n635), .ZN(n531) );
  NAND2_X1 U584 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U585 ( .A(KEYINPUT9), .B(n533), .Z(n534) );
  XNOR2_X1 U586 ( .A(KEYINPUT70), .B(n534), .ZN(n535) );
  NOR2_X1 U587 ( .A1(n536), .A2(n535), .ZN(G171) );
  AND2_X1 U588 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U589 ( .A(G69), .ZN(G235) );
  INV_X1 U590 ( .A(G132), .ZN(G219) );
  INV_X1 U591 ( .A(G82), .ZN(G220) );
  NAND2_X1 U592 ( .A1(G51), .A2(n639), .ZN(n537) );
  XNOR2_X1 U593 ( .A(n537), .B(KEYINPUT74), .ZN(n539) );
  NAND2_X1 U594 ( .A1(G63), .A2(n631), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U596 ( .A(KEYINPUT6), .B(n540), .ZN(n547) );
  NAND2_X1 U597 ( .A1(n632), .A2(G89), .ZN(n541) );
  XNOR2_X1 U598 ( .A(n541), .B(KEYINPUT4), .ZN(n543) );
  NAND2_X1 U599 ( .A1(G76), .A2(n635), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U601 ( .A(KEYINPUT73), .B(n544), .ZN(n545) );
  XNOR2_X1 U602 ( .A(KEYINPUT5), .B(n545), .ZN(n546) );
  NOR2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U604 ( .A(KEYINPUT7), .B(n548), .Z(G168) );
  XOR2_X1 U605 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U606 ( .A1(G7), .A2(G661), .ZN(n549) );
  XNOR2_X1 U607 ( .A(n549), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U608 ( .A(G223), .ZN(n819) );
  NAND2_X1 U609 ( .A1(n819), .A2(G567), .ZN(n550) );
  XOR2_X1 U610 ( .A(KEYINPUT11), .B(n550), .Z(G234) );
  NAND2_X1 U611 ( .A1(G56), .A2(n631), .ZN(n551) );
  XOR2_X1 U612 ( .A(KEYINPUT14), .B(n551), .Z(n557) );
  NAND2_X1 U613 ( .A1(n632), .A2(G81), .ZN(n552) );
  XNOR2_X1 U614 ( .A(n552), .B(KEYINPUT12), .ZN(n554) );
  NAND2_X1 U615 ( .A1(G68), .A2(n635), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U617 ( .A(KEYINPUT13), .B(n555), .Z(n556) );
  NOR2_X1 U618 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U619 ( .A1(G43), .A2(n639), .ZN(n558) );
  NAND2_X1 U620 ( .A1(n559), .A2(n558), .ZN(n961) );
  INV_X1 U621 ( .A(G860), .ZN(n581) );
  OR2_X1 U622 ( .A1(n961), .A2(n581), .ZN(G153) );
  INV_X1 U623 ( .A(G171), .ZN(G301) );
  NAND2_X1 U624 ( .A1(G868), .A2(G301), .ZN(n570) );
  NAND2_X1 U625 ( .A1(n632), .A2(G92), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n635), .A2(G79), .ZN(n561) );
  NAND2_X1 U627 ( .A1(G54), .A2(n639), .ZN(n560) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT72), .B(n562), .ZN(n565) );
  NAND2_X1 U630 ( .A1(G66), .A2(n631), .ZN(n563) );
  XNOR2_X1 U631 ( .A(KEYINPUT71), .B(n563), .ZN(n564) );
  NOR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT15), .B(n568), .Z(n977) );
  INV_X1 U635 ( .A(G868), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n977), .A2(n577), .ZN(n569) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(G284) );
  NAND2_X1 U638 ( .A1(n631), .A2(G65), .ZN(n572) );
  NAND2_X1 U639 ( .A1(G53), .A2(n639), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G91), .A2(n632), .ZN(n574) );
  NAND2_X1 U642 ( .A1(G78), .A2(n635), .ZN(n573) );
  NAND2_X1 U643 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n958) );
  INV_X1 U645 ( .A(n958), .ZN(G299) );
  NOR2_X1 U646 ( .A1(G868), .A2(G299), .ZN(n579) );
  NOR2_X1 U647 ( .A1(G286), .A2(n577), .ZN(n578) );
  NOR2_X1 U648 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U649 ( .A(KEYINPUT75), .B(n580), .Z(G297) );
  NAND2_X1 U650 ( .A1(n581), .A2(G559), .ZN(n582) );
  INV_X1 U651 ( .A(n977), .ZN(n887) );
  NAND2_X1 U652 ( .A1(n582), .A2(n887), .ZN(n583) );
  XNOR2_X1 U653 ( .A(n583), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U654 ( .A1(G868), .A2(n961), .ZN(n586) );
  NAND2_X1 U655 ( .A1(G868), .A2(n887), .ZN(n584) );
  NOR2_X1 U656 ( .A1(G559), .A2(n584), .ZN(n585) );
  NOR2_X1 U657 ( .A1(n586), .A2(n585), .ZN(G282) );
  NAND2_X1 U658 ( .A1(G99), .A2(n874), .ZN(n587) );
  XNOR2_X1 U659 ( .A(n587), .B(KEYINPUT78), .ZN(n598) );
  NAND2_X1 U660 ( .A1(n869), .A2(G123), .ZN(n588) );
  XNOR2_X1 U661 ( .A(n588), .B(KEYINPUT18), .ZN(n592) );
  INV_X1 U662 ( .A(n589), .ZN(n590) );
  NAND2_X1 U663 ( .A1(G135), .A2(n875), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U665 ( .A(KEYINPUT76), .B(n593), .ZN(n596) );
  NAND2_X1 U666 ( .A1(G111), .A2(n870), .ZN(n594) );
  XNOR2_X1 U667 ( .A(KEYINPUT77), .B(n594), .ZN(n595) );
  NOR2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n1002) );
  XNOR2_X1 U670 ( .A(n1002), .B(G2096), .ZN(n599) );
  XNOR2_X1 U671 ( .A(n599), .B(KEYINPUT79), .ZN(n601) );
  INV_X1 U672 ( .A(G2100), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n601), .A2(n600), .ZN(G156) );
  NAND2_X1 U674 ( .A1(n887), .A2(G559), .ZN(n649) );
  XNOR2_X1 U675 ( .A(n961), .B(n649), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n602), .A2(G860), .ZN(n610) );
  NAND2_X1 U677 ( .A1(G93), .A2(n632), .ZN(n603) );
  XNOR2_X1 U678 ( .A(n603), .B(KEYINPUT80), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n631), .A2(G67), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n635), .A2(G80), .ZN(n607) );
  NAND2_X1 U682 ( .A1(G55), .A2(n639), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n651) );
  XNOR2_X1 U685 ( .A(n610), .B(n651), .ZN(G145) );
  NAND2_X1 U686 ( .A1(G88), .A2(n632), .ZN(n612) );
  NAND2_X1 U687 ( .A1(G75), .A2(n635), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n631), .A2(G62), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G50), .A2(n639), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U692 ( .A1(n616), .A2(n615), .ZN(G166) );
  NAND2_X1 U693 ( .A1(n617), .A2(G87), .ZN(n622) );
  NAND2_X1 U694 ( .A1(G651), .A2(G74), .ZN(n619) );
  NAND2_X1 U695 ( .A1(G49), .A2(n639), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U697 ( .A1(n631), .A2(n620), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U699 ( .A(KEYINPUT81), .B(n623), .Z(G288) );
  NAND2_X1 U700 ( .A1(G61), .A2(n631), .ZN(n625) );
  NAND2_X1 U701 ( .A1(G86), .A2(n632), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n635), .A2(G73), .ZN(n626) );
  XOR2_X1 U704 ( .A(KEYINPUT2), .B(n626), .Z(n627) );
  NOR2_X1 U705 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U706 ( .A1(G48), .A2(n639), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(G305) );
  NAND2_X1 U708 ( .A1(G60), .A2(n631), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G85), .A2(n632), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U711 ( .A1(n635), .A2(G72), .ZN(n636) );
  XOR2_X1 U712 ( .A(KEYINPUT68), .B(n636), .Z(n637) );
  NOR2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U714 ( .A1(G47), .A2(n639), .ZN(n640) );
  NAND2_X1 U715 ( .A1(n641), .A2(n640), .ZN(G290) );
  XNOR2_X1 U716 ( .A(n958), .B(n651), .ZN(n648) );
  XNOR2_X1 U717 ( .A(G166), .B(KEYINPUT19), .ZN(n642) );
  XNOR2_X1 U718 ( .A(n642), .B(KEYINPUT82), .ZN(n643) );
  XNOR2_X1 U719 ( .A(n643), .B(n961), .ZN(n644) );
  XNOR2_X1 U720 ( .A(n644), .B(G288), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n645), .B(G305), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n646), .B(G290), .ZN(n647) );
  XNOR2_X1 U723 ( .A(n648), .B(n647), .ZN(n888) );
  XNOR2_X1 U724 ( .A(n649), .B(n888), .ZN(n650) );
  NAND2_X1 U725 ( .A1(n650), .A2(G868), .ZN(n653) );
  OR2_X1 U726 ( .A1(G868), .A2(n651), .ZN(n652) );
  NAND2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U728 ( .A(KEYINPUT83), .B(n654), .Z(G295) );
  NAND2_X1 U729 ( .A1(G2078), .A2(G2084), .ZN(n655) );
  XOR2_X1 U730 ( .A(KEYINPUT20), .B(n655), .Z(n656) );
  NAND2_X1 U731 ( .A1(G2090), .A2(n656), .ZN(n657) );
  XNOR2_X1 U732 ( .A(KEYINPUT21), .B(n657), .ZN(n658) );
  NAND2_X1 U733 ( .A1(n658), .A2(G2072), .ZN(n659) );
  XNOR2_X1 U734 ( .A(KEYINPUT84), .B(n659), .ZN(G158) );
  XNOR2_X1 U735 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U736 ( .A1(G220), .A2(G219), .ZN(n660) );
  XOR2_X1 U737 ( .A(KEYINPUT22), .B(n660), .Z(n661) );
  NOR2_X1 U738 ( .A1(G218), .A2(n661), .ZN(n662) );
  NAND2_X1 U739 ( .A1(G96), .A2(n662), .ZN(n824) );
  NAND2_X1 U740 ( .A1(G2106), .A2(n824), .ZN(n666) );
  NAND2_X1 U741 ( .A1(G120), .A2(G108), .ZN(n663) );
  NOR2_X1 U742 ( .A1(G235), .A2(n663), .ZN(n664) );
  NAND2_X1 U743 ( .A1(G57), .A2(n664), .ZN(n825) );
  NAND2_X1 U744 ( .A1(G567), .A2(n825), .ZN(n665) );
  NAND2_X1 U745 ( .A1(n666), .A2(n665), .ZN(n826) );
  NAND2_X1 U746 ( .A1(G661), .A2(G483), .ZN(n667) );
  NOR2_X1 U747 ( .A1(n826), .A2(n667), .ZN(n823) );
  NAND2_X1 U748 ( .A1(n823), .A2(G36), .ZN(G176) );
  NAND2_X1 U749 ( .A1(n874), .A2(G102), .ZN(n670) );
  NAND2_X1 U750 ( .A1(G114), .A2(n870), .ZN(n668) );
  XOR2_X1 U751 ( .A(KEYINPUT85), .B(n668), .Z(n669) );
  NAND2_X1 U752 ( .A1(n670), .A2(n669), .ZN(n674) );
  NAND2_X1 U753 ( .A1(n869), .A2(G126), .ZN(n672) );
  NAND2_X1 U754 ( .A1(G138), .A2(n875), .ZN(n671) );
  NAND2_X1 U755 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U756 ( .A1(n674), .A2(n673), .ZN(G164) );
  INV_X1 U757 ( .A(G166), .ZN(G303) );
  NAND2_X1 U758 ( .A1(G160), .A2(G40), .ZN(n768) );
  INV_X1 U759 ( .A(n768), .ZN(n675) );
  NOR2_X1 U760 ( .A1(G164), .A2(G1384), .ZN(n769) );
  NAND2_X1 U761 ( .A1(n675), .A2(n769), .ZN(n717) );
  INV_X1 U762 ( .A(n717), .ZN(n697) );
  NAND2_X1 U763 ( .A1(n697), .A2(G2072), .ZN(n676) );
  XNOR2_X1 U764 ( .A(n676), .B(KEYINPUT27), .ZN(n678) );
  INV_X1 U765 ( .A(G1956), .ZN(n934) );
  NOR2_X1 U766 ( .A1(n934), .A2(n697), .ZN(n677) );
  NOR2_X1 U767 ( .A1(n678), .A2(n677), .ZN(n680) );
  NOR2_X1 U768 ( .A1(n958), .A2(n680), .ZN(n679) );
  XOR2_X1 U769 ( .A(n679), .B(KEYINPUT28), .Z(n695) );
  NAND2_X1 U770 ( .A1(n958), .A2(n680), .ZN(n693) );
  AND2_X1 U771 ( .A1(n697), .A2(G1996), .ZN(n681) );
  XOR2_X1 U772 ( .A(n681), .B(KEYINPUT26), .Z(n683) );
  NAND2_X1 U773 ( .A1(n717), .A2(G1341), .ZN(n682) );
  NAND2_X1 U774 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U775 ( .A1(n961), .A2(n684), .ZN(n688) );
  NAND2_X1 U776 ( .A1(G1348), .A2(n717), .ZN(n686) );
  NAND2_X1 U777 ( .A1(n697), .A2(G2067), .ZN(n685) );
  NAND2_X1 U778 ( .A1(n686), .A2(n685), .ZN(n689) );
  NOR2_X1 U779 ( .A1(n977), .A2(n689), .ZN(n687) );
  OR2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n691) );
  NAND2_X1 U781 ( .A1(n977), .A2(n689), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U783 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U784 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U785 ( .A(n696), .B(KEYINPUT29), .ZN(n702) );
  NAND2_X1 U786 ( .A1(n717), .A2(G1961), .ZN(n699) );
  XOR2_X1 U787 ( .A(G2078), .B(KEYINPUT25), .Z(n911) );
  NAND2_X1 U788 ( .A1(n697), .A2(n911), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U790 ( .A(n700), .B(KEYINPUT92), .Z(n708) );
  AND2_X1 U791 ( .A1(G171), .A2(n708), .ZN(n701) );
  NOR2_X1 U792 ( .A1(n702), .A2(n701), .ZN(n713) );
  XOR2_X1 U793 ( .A(KEYINPUT91), .B(n703), .Z(n729) );
  NAND2_X1 U794 ( .A1(G8), .A2(n717), .ZN(n763) );
  NOR2_X1 U795 ( .A1(G1966), .A2(n763), .ZN(n732) );
  NOR2_X1 U796 ( .A1(n729), .A2(n732), .ZN(n704) );
  XOR2_X1 U797 ( .A(KEYINPUT93), .B(n704), .Z(n705) );
  NAND2_X1 U798 ( .A1(G8), .A2(n705), .ZN(n706) );
  XNOR2_X1 U799 ( .A(KEYINPUT30), .B(n706), .ZN(n707) );
  NOR2_X1 U800 ( .A1(G168), .A2(n707), .ZN(n710) );
  NOR2_X1 U801 ( .A1(G171), .A2(n708), .ZN(n709) );
  NOR2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U803 ( .A(n711), .B(KEYINPUT31), .ZN(n712) );
  NOR2_X1 U804 ( .A1(n713), .A2(n712), .ZN(n715) );
  INV_X1 U805 ( .A(KEYINPUT94), .ZN(n714) );
  XNOR2_X1 U806 ( .A(n715), .B(n714), .ZN(n730) );
  AND2_X1 U807 ( .A1(G286), .A2(G8), .ZN(n716) );
  NAND2_X1 U808 ( .A1(n730), .A2(n716), .ZN(n726) );
  INV_X1 U809 ( .A(G8), .ZN(n724) );
  NOR2_X1 U810 ( .A1(G2090), .A2(n717), .ZN(n718) );
  XOR2_X1 U811 ( .A(KEYINPUT96), .B(n718), .Z(n719) );
  NAND2_X1 U812 ( .A1(n719), .A2(G303), .ZN(n721) );
  NOR2_X1 U813 ( .A1(G1971), .A2(n763), .ZN(n720) );
  NOR2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U815 ( .A(n722), .B(KEYINPUT97), .ZN(n723) );
  OR2_X1 U816 ( .A1(n724), .A2(n723), .ZN(n725) );
  AND2_X1 U817 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U818 ( .A(n727), .B(KEYINPUT98), .ZN(n728) );
  XNOR2_X1 U819 ( .A(n728), .B(KEYINPUT32), .ZN(n736) );
  NAND2_X1 U820 ( .A1(n729), .A2(G8), .ZN(n734) );
  XNOR2_X1 U821 ( .A(KEYINPUT95), .B(n730), .ZN(n731) );
  NOR2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U823 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U824 ( .A1(n736), .A2(n735), .ZN(n754) );
  NOR2_X1 U825 ( .A1(G2090), .A2(G303), .ZN(n737) );
  NAND2_X1 U826 ( .A1(G8), .A2(n737), .ZN(n738) );
  XNOR2_X1 U827 ( .A(n738), .B(KEYINPUT102), .ZN(n743) );
  NOR2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n750) );
  XOR2_X1 U829 ( .A(n750), .B(KEYINPUT100), .Z(n739) );
  NOR2_X1 U830 ( .A1(n763), .A2(n739), .ZN(n741) );
  XOR2_X1 U831 ( .A(KEYINPUT101), .B(G1981), .Z(n740) );
  XNOR2_X1 U832 ( .A(G305), .B(n740), .ZN(n968) );
  NOR2_X1 U833 ( .A1(n741), .A2(n968), .ZN(n742) );
  NAND2_X1 U834 ( .A1(KEYINPUT33), .A2(n742), .ZN(n745) );
  AND2_X1 U835 ( .A1(n743), .A2(n745), .ZN(n744) );
  NAND2_X1 U836 ( .A1(n754), .A2(n744), .ZN(n748) );
  INV_X1 U837 ( .A(n745), .ZN(n746) );
  OR2_X1 U838 ( .A1(n746), .A2(n763), .ZN(n747) );
  AND2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n767) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U841 ( .A1(n750), .A2(n749), .ZN(n976) );
  NOR2_X1 U842 ( .A1(G1981), .A2(G305), .ZN(n751) );
  XNOR2_X1 U843 ( .A(n751), .B(KEYINPUT24), .ZN(n761) );
  INV_X1 U844 ( .A(n761), .ZN(n752) );
  AND2_X1 U845 ( .A1(n976), .A2(n752), .ZN(n753) );
  NAND2_X1 U846 ( .A1(n754), .A2(n753), .ZN(n765) );
  NAND2_X1 U847 ( .A1(G288), .A2(G1976), .ZN(n755) );
  XOR2_X1 U848 ( .A(KEYINPUT99), .B(n755), .Z(n965) );
  INV_X1 U849 ( .A(KEYINPUT33), .ZN(n756) );
  AND2_X1 U850 ( .A1(KEYINPUT100), .A2(n756), .ZN(n758) );
  INV_X1 U851 ( .A(n968), .ZN(n757) );
  AND2_X1 U852 ( .A1(n758), .A2(n757), .ZN(n759) );
  AND2_X1 U853 ( .A1(n965), .A2(n759), .ZN(n760) );
  NOR2_X1 U854 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n764) );
  AND2_X1 U856 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U857 ( .A1(n767), .A2(n766), .ZN(n803) );
  NOR2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n813) );
  XNOR2_X1 U859 ( .A(G2067), .B(KEYINPUT37), .ZN(n804) );
  NAND2_X1 U860 ( .A1(G140), .A2(n875), .ZN(n770) );
  XNOR2_X1 U861 ( .A(KEYINPUT87), .B(n770), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n874), .A2(G104), .ZN(n771) );
  XOR2_X1 U863 ( .A(KEYINPUT86), .B(n771), .Z(n772) );
  NOR2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U865 ( .A(KEYINPUT34), .B(n774), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n869), .A2(G128), .ZN(n775) );
  XNOR2_X1 U867 ( .A(n775), .B(KEYINPUT88), .ZN(n777) );
  NAND2_X1 U868 ( .A1(G116), .A2(n870), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U870 ( .A(KEYINPUT35), .B(n778), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U872 ( .A(n781), .B(KEYINPUT36), .ZN(n782) );
  XNOR2_X1 U873 ( .A(KEYINPUT89), .B(n782), .ZN(n883) );
  NOR2_X1 U874 ( .A1(n804), .A2(n883), .ZN(n1012) );
  NAND2_X1 U875 ( .A1(n813), .A2(n1012), .ZN(n811) );
  NOR2_X1 U876 ( .A1(G1986), .A2(G290), .ZN(n974) );
  XOR2_X1 U877 ( .A(KEYINPUT90), .B(KEYINPUT38), .Z(n784) );
  NAND2_X1 U878 ( .A1(G105), .A2(n874), .ZN(n783) );
  XNOR2_X1 U879 ( .A(n784), .B(n783), .ZN(n788) );
  NAND2_X1 U880 ( .A1(n869), .A2(G129), .ZN(n786) );
  NAND2_X1 U881 ( .A1(G141), .A2(n875), .ZN(n785) );
  NAND2_X1 U882 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U883 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U884 ( .A1(n870), .A2(G117), .ZN(n789) );
  NAND2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n861) );
  NAND2_X1 U886 ( .A1(G1996), .A2(n861), .ZN(n798) );
  NAND2_X1 U887 ( .A1(G95), .A2(n874), .ZN(n792) );
  NAND2_X1 U888 ( .A1(G119), .A2(n869), .ZN(n791) );
  NAND2_X1 U889 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U890 ( .A1(n870), .A2(G107), .ZN(n794) );
  NAND2_X1 U891 ( .A1(G131), .A2(n875), .ZN(n793) );
  NAND2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U893 ( .A1(n796), .A2(n795), .ZN(n862) );
  NAND2_X1 U894 ( .A1(G1991), .A2(n862), .ZN(n797) );
  NAND2_X1 U895 ( .A1(n798), .A2(n797), .ZN(n996) );
  NOR2_X1 U896 ( .A1(n974), .A2(n996), .ZN(n799) );
  NAND2_X1 U897 ( .A1(G1986), .A2(G290), .ZN(n959) );
  NAND2_X1 U898 ( .A1(n799), .A2(n959), .ZN(n800) );
  NAND2_X1 U899 ( .A1(n800), .A2(n813), .ZN(n801) );
  NAND2_X1 U900 ( .A1(n804), .A2(n883), .ZN(n1009) );
  XOR2_X1 U901 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n809) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n861), .ZN(n1005) );
  NOR2_X1 U903 ( .A1(G1991), .A2(n862), .ZN(n997) );
  NOR2_X1 U904 ( .A1(n974), .A2(n997), .ZN(n805) );
  XOR2_X1 U905 ( .A(KEYINPUT103), .B(n805), .Z(n806) );
  NOR2_X1 U906 ( .A1(n996), .A2(n806), .ZN(n807) );
  NOR2_X1 U907 ( .A1(n1005), .A2(n807), .ZN(n808) );
  XOR2_X1 U908 ( .A(n809), .B(n808), .Z(n810) );
  NAND2_X1 U909 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n1009), .A2(n812), .ZN(n814) );
  NAND2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U912 ( .A1(n816), .A2(n815), .ZN(n818) );
  XOR2_X1 U913 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n817) );
  XNOR2_X1 U914 ( .A(n818), .B(n817), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n819), .ZN(G217) );
  NAND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n820) );
  XOR2_X1 U917 ( .A(KEYINPUT108), .B(n820), .Z(n821) );
  NAND2_X1 U918 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n822) );
  NAND2_X1 U920 ( .A1(n823), .A2(n822), .ZN(G188) );
  XNOR2_X1 U921 ( .A(G120), .B(KEYINPUT109), .ZN(G236) );
  XNOR2_X1 U922 ( .A(G108), .B(KEYINPUT115), .ZN(G238) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  NOR2_X1 U925 ( .A1(n825), .A2(n824), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  XOR2_X1 U927 ( .A(KEYINPUT110), .B(n826), .Z(G319) );
  XOR2_X1 U928 ( .A(G2678), .B(G2090), .Z(n828) );
  XNOR2_X1 U929 ( .A(G2078), .B(G2072), .ZN(n827) );
  XNOR2_X1 U930 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U931 ( .A(n829), .B(G2100), .Z(n831) );
  XNOR2_X1 U932 ( .A(G2067), .B(G2084), .ZN(n830) );
  XNOR2_X1 U933 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U934 ( .A(G2096), .B(KEYINPUT111), .Z(n833) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n832) );
  XNOR2_X1 U936 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U937 ( .A(n835), .B(n834), .Z(G227) );
  XOR2_X1 U938 ( .A(G1986), .B(G1976), .Z(n837) );
  XNOR2_X1 U939 ( .A(G1966), .B(G1981), .ZN(n836) );
  XNOR2_X1 U940 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U941 ( .A(n838), .B(G2474), .Z(n840) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n839) );
  XNOR2_X1 U943 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U944 ( .A(KEYINPUT41), .B(G1971), .Z(n842) );
  XNOR2_X1 U945 ( .A(G1961), .B(G1956), .ZN(n841) );
  XNOR2_X1 U946 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U947 ( .A(n844), .B(n843), .ZN(G229) );
  NAND2_X1 U948 ( .A1(G100), .A2(n874), .ZN(n846) );
  NAND2_X1 U949 ( .A1(G112), .A2(n870), .ZN(n845) );
  NAND2_X1 U950 ( .A1(n846), .A2(n845), .ZN(n847) );
  XNOR2_X1 U951 ( .A(KEYINPUT112), .B(n847), .ZN(n852) );
  NAND2_X1 U952 ( .A1(G124), .A2(n869), .ZN(n848) );
  XNOR2_X1 U953 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U954 ( .A1(G136), .A2(n875), .ZN(n849) );
  NAND2_X1 U955 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U956 ( .A1(n852), .A2(n851), .ZN(G162) );
  NAND2_X1 U957 ( .A1(n874), .A2(G103), .ZN(n854) );
  NAND2_X1 U958 ( .A1(G139), .A2(n875), .ZN(n853) );
  NAND2_X1 U959 ( .A1(n854), .A2(n853), .ZN(n859) );
  NAND2_X1 U960 ( .A1(G127), .A2(n869), .ZN(n856) );
  NAND2_X1 U961 ( .A1(G115), .A2(n870), .ZN(n855) );
  NAND2_X1 U962 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U963 ( .A(KEYINPUT47), .B(n857), .Z(n858) );
  NOR2_X1 U964 ( .A1(n859), .A2(n858), .ZN(n991) );
  XOR2_X1 U965 ( .A(G162), .B(n991), .Z(n860) );
  XNOR2_X1 U966 ( .A(n861), .B(n860), .ZN(n866) );
  XNOR2_X1 U967 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n864) );
  XNOR2_X1 U968 ( .A(n862), .B(KEYINPUT46), .ZN(n863) );
  XNOR2_X1 U969 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U970 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U971 ( .A(G160), .B(G164), .ZN(n867) );
  XNOR2_X1 U972 ( .A(n868), .B(n867), .ZN(n885) );
  NAND2_X1 U973 ( .A1(G130), .A2(n869), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G118), .A2(n870), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U976 ( .A(KEYINPUT113), .B(n873), .Z(n880) );
  NAND2_X1 U977 ( .A1(n874), .A2(G106), .ZN(n877) );
  NAND2_X1 U978 ( .A1(G142), .A2(n875), .ZN(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U980 ( .A(n878), .B(KEYINPUT45), .Z(n879) );
  NOR2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U982 ( .A(n881), .B(n1002), .ZN(n882) );
  XOR2_X1 U983 ( .A(n883), .B(n882), .Z(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n886) );
  NOR2_X1 U985 ( .A1(G37), .A2(n886), .ZN(G395) );
  XOR2_X1 U986 ( .A(n888), .B(n887), .Z(n890) );
  XNOR2_X1 U987 ( .A(G286), .B(G171), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U989 ( .A1(G37), .A2(n891), .ZN(G397) );
  XNOR2_X1 U990 ( .A(G2451), .B(G2427), .ZN(n901) );
  XOR2_X1 U991 ( .A(KEYINPUT107), .B(G2443), .Z(n893) );
  XNOR2_X1 U992 ( .A(G2435), .B(G2438), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n893), .B(n892), .ZN(n897) );
  XOR2_X1 U994 ( .A(G2454), .B(G2430), .Z(n895) );
  XNOR2_X1 U995 ( .A(G1341), .B(G1348), .ZN(n894) );
  XNOR2_X1 U996 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U997 ( .A(n897), .B(n896), .Z(n899) );
  XNOR2_X1 U998 ( .A(G2446), .B(KEYINPUT106), .ZN(n898) );
  XNOR2_X1 U999 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n902) );
  NAND2_X1 U1001 ( .A1(n902), .A2(G14), .ZN(n908) );
  NAND2_X1 U1002 ( .A1(n908), .A2(G319), .ZN(n905) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n903), .ZN(n904) );
  NOR2_X1 U1005 ( .A1(n905), .A2(n904), .ZN(n907) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1007 ( .A1(n907), .A2(n906), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G57), .ZN(G237) );
  INV_X1 U1010 ( .A(n908), .ZN(G401) );
  XNOR2_X1 U1011 ( .A(G25), .B(G1991), .ZN(n909) );
  XNOR2_X1 U1012 ( .A(n909), .B(KEYINPUT117), .ZN(n920) );
  XOR2_X1 U1013 ( .A(G2067), .B(G26), .Z(n910) );
  NAND2_X1 U1014 ( .A1(n910), .A2(G28), .ZN(n918) );
  XOR2_X1 U1015 ( .A(G2072), .B(G33), .Z(n916) );
  XNOR2_X1 U1016 ( .A(n911), .B(G27), .ZN(n913) );
  XNOR2_X1 U1017 ( .A(G32), .B(G1996), .ZN(n912) );
  NOR2_X1 U1018 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1019 ( .A(KEYINPUT118), .B(n914), .ZN(n915) );
  NAND2_X1 U1020 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1021 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1023 ( .A(n921), .B(KEYINPUT53), .ZN(n924) );
  XOR2_X1 U1024 ( .A(G2084), .B(G34), .Z(n922) );
  XNOR2_X1 U1025 ( .A(KEYINPUT54), .B(n922), .ZN(n923) );
  NAND2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(G35), .B(G2090), .ZN(n925) );
  NOR2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1029 ( .A(KEYINPUT55), .B(n927), .Z(n928) );
  NOR2_X1 U1030 ( .A1(G29), .A2(n928), .ZN(n957) );
  XOR2_X1 U1031 ( .A(G1961), .B(G5), .Z(n944) );
  XNOR2_X1 U1032 ( .A(G1348), .B(KEYINPUT59), .ZN(n929) );
  XNOR2_X1 U1033 ( .A(n929), .B(G4), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(G1341), .B(G19), .ZN(n931) );
  XNOR2_X1 U1035 ( .A(G6), .B(G1981), .ZN(n930) );
  NOR2_X1 U1036 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1037 ( .A1(n933), .A2(n932), .ZN(n937) );
  XOR2_X1 U1038 ( .A(KEYINPUT124), .B(n934), .Z(n935) );
  XNOR2_X1 U1039 ( .A(G20), .B(n935), .ZN(n936) );
  NOR2_X1 U1040 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1041 ( .A(n938), .B(KEYINPUT125), .ZN(n939) );
  XNOR2_X1 U1042 ( .A(n939), .B(KEYINPUT60), .ZN(n941) );
  XNOR2_X1 U1043 ( .A(G21), .B(G1966), .ZN(n940) );
  NOR2_X1 U1044 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1045 ( .A(KEYINPUT126), .B(n942), .ZN(n943) );
  NAND2_X1 U1046 ( .A1(n944), .A2(n943), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(G1971), .B(G22), .ZN(n946) );
  XNOR2_X1 U1048 ( .A(G23), .B(G1976), .ZN(n945) );
  NOR2_X1 U1049 ( .A1(n946), .A2(n945), .ZN(n948) );
  XOR2_X1 U1050 ( .A(G1986), .B(G24), .Z(n947) );
  NAND2_X1 U1051 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1052 ( .A(KEYINPUT58), .B(n949), .ZN(n950) );
  NOR2_X1 U1053 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1054 ( .A(n952), .B(KEYINPUT61), .ZN(n954) );
  XNOR2_X1 U1055 ( .A(G16), .B(KEYINPUT123), .ZN(n953) );
  NAND2_X1 U1056 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n955), .ZN(n956) );
  NOR2_X1 U1058 ( .A1(n957), .A2(n956), .ZN(n989) );
  XNOR2_X1 U1059 ( .A(n958), .B(G1956), .ZN(n960) );
  NAND2_X1 U1060 ( .A1(n960), .A2(n959), .ZN(n964) );
  XOR2_X1 U1061 ( .A(G1341), .B(n961), .Z(n962) );
  XNOR2_X1 U1062 ( .A(KEYINPUT121), .B(n962), .ZN(n963) );
  NOR2_X1 U1063 ( .A1(n964), .A2(n963), .ZN(n966) );
  NAND2_X1 U1064 ( .A1(n966), .A2(n965), .ZN(n984) );
  XOR2_X1 U1065 ( .A(G168), .B(G1966), .Z(n967) );
  NOR2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1067 ( .A(KEYINPUT57), .B(n969), .ZN(n970) );
  XNOR2_X1 U1068 ( .A(n970), .B(KEYINPUT119), .ZN(n982) );
  XNOR2_X1 U1069 ( .A(G171), .B(G1961), .ZN(n972) );
  NAND2_X1 U1070 ( .A1(G1971), .A2(G303), .ZN(n971) );
  NAND2_X1 U1071 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1072 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(G1348), .B(n977), .ZN(n978) );
  XNOR2_X1 U1075 ( .A(KEYINPUT120), .B(n978), .ZN(n979) );
  NOR2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1079 ( .A(KEYINPUT122), .B(n985), .Z(n987) );
  XNOR2_X1 U1080 ( .A(KEYINPUT56), .B(G16), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(n990), .B(KEYINPUT127), .ZN(n1018) );
  XOR2_X1 U1084 ( .A(G2072), .B(n991), .Z(n993) );
  XOR2_X1 U1085 ( .A(G164), .B(G2078), .Z(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1087 ( .A(KEYINPUT50), .B(n994), .ZN(n995) );
  XNOR2_X1 U1088 ( .A(n995), .B(KEYINPUT116), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XOR2_X1 U1091 ( .A(G160), .B(G2084), .Z(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1008) );
  XOR2_X1 U1094 ( .A(G2090), .B(G162), .Z(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(n1006), .B(KEYINPUT51), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(KEYINPUT52), .B(n1013), .ZN(n1015) );
  INV_X1 U1101 ( .A(KEYINPUT55), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(G29), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1019), .Z(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

