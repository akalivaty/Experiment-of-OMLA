//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1029, new_n1030;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT12), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G229gat), .A2(G233gat), .ZN(new_n209));
  XOR2_X1   g008(.A(new_n209), .B(KEYINPUT13), .Z(new_n210));
  AND2_X1   g009(.A1(G43gat), .A2(G50gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G43gat), .A2(G50gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT15), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT90), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n214), .B(new_n215), .C1(G29gat), .C2(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G29gat), .ZN(new_n220));
  INV_X1    g019(.A(G36gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT90), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n214), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT14), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n213), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G43gat), .ZN(new_n226));
  INV_X1    g025(.A(G50gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT15), .ZN(new_n229));
  NAND2_X1  g028(.A1(G43gat), .A2(G50gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n229), .B1(new_n228), .B2(new_n230), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT91), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n228), .A2(KEYINPUT91), .A3(new_n229), .A4(new_n230), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n234), .A2(new_n224), .A3(new_n219), .A4(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT92), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n225), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G8gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(KEYINPUT94), .ZN(new_n240));
  XNOR2_X1  g039(.A(G15gat), .B(G22gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT16), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G22gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G15gat), .ZN(new_n245));
  INV_X1    g044(.A(G15gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G22gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT93), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G1gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n241), .A2(new_n248), .A3(G1gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n243), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n239), .A2(KEYINPUT94), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n243), .A2(new_n251), .A3(new_n252), .A4(new_n254), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n220), .A2(new_n221), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n215), .B1(new_n259), .B2(new_n214), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n218), .B1(new_n222), .B2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n261), .A2(KEYINPUT92), .A3(new_n234), .A4(new_n235), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n238), .A2(new_n258), .A3(KEYINPUT95), .A4(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n256), .A2(new_n257), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT15), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n265), .B1(KEYINPUT91), .B2(new_n213), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n224), .A2(new_n235), .A3(new_n217), .A4(new_n216), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n237), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n225), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n262), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n268), .A2(new_n262), .A3(new_n269), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT95), .B1(new_n273), .B2(new_n258), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n210), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT96), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT96), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n277), .B(new_n210), .C1(new_n272), .C2(new_n274), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT17), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n270), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n268), .A2(new_n262), .A3(KEYINPUT17), .A4(new_n269), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(new_n258), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(new_n209), .A3(new_n271), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT18), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n258), .B1(new_n238), .B2(new_n262), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n270), .A2(new_n280), .B1(new_n257), .B2(new_n256), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n286), .B1(new_n287), .B2(new_n282), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n285), .B1(G229gat), .B2(G233gat), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n284), .A2(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n208), .B1(new_n279), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n278), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT95), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(new_n264), .B2(new_n270), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(new_n271), .A3(new_n263), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n277), .B1(new_n295), .B2(new_n210), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n207), .B1(new_n288), .B2(new_n289), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n284), .A2(new_n285), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT97), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT18), .B1(new_n288), .B2(new_n209), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n283), .A2(new_n271), .A3(new_n289), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n208), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT97), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n279), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n291), .B1(new_n301), .B2(new_n307), .ZN(new_n308));
  XOR2_X1   g107(.A(KEYINPUT67), .B(G190gat), .Z(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT27), .B(G183gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT26), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n318), .A2(new_n319), .B1(new_n317), .B2(new_n316), .ZN(new_n320));
  OAI211_X1 g119(.A(KEYINPUT69), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n311), .A2(new_n312), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n313), .A2(new_n314), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT23), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n316), .B(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n315), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT65), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT24), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n330), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n331), .A2(KEYINPUT64), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(KEYINPUT64), .ZN(new_n333));
  NAND3_X1  g132(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n334));
  OR2_X1    g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT25), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n326), .A2(KEYINPUT65), .A3(new_n315), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n329), .A2(new_n336), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n315), .B(KEYINPUT66), .Z(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT67), .B(G190gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(G183gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n331), .A2(new_n334), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n340), .B(new_n326), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT25), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n324), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n347), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT73), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G197gat), .B(G204gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT22), .ZN(new_n357));
  INV_X1    g156(.A(G211gat), .ZN(new_n358));
  INV_X1    g157(.A(G218gat), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G211gat), .B(G218gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n349), .A2(new_n351), .ZN(new_n365));
  INV_X1    g164(.A(new_n363), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G8gat), .B(G36gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(G64gat), .B(G92gat), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  NAND3_X1  g169(.A1(new_n364), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT30), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT74), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n366), .B1(new_n352), .B2(new_n354), .ZN(new_n374));
  INV_X1    g173(.A(new_n367), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT74), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT30), .A4(new_n370), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n370), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(new_n374), .B2(new_n375), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT75), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n382), .B1(new_n371), .B2(new_n372), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n371), .A2(new_n382), .A3(new_n372), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n379), .B(new_n381), .C1(new_n383), .C2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT5), .ZN(new_n387));
  INV_X1    g186(.A(G113gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G120gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT71), .B(G120gat), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(new_n388), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT72), .ZN(new_n392));
  INV_X1    g191(.A(G134gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(G127gat), .ZN(new_n394));
  INV_X1    g193(.A(G127gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n395), .A2(G134gat), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n394), .A2(new_n396), .A3(KEYINPUT1), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G113gat), .B(G120gat), .ZN(new_n399));
  OR2_X1    g198(.A1(new_n399), .A2(KEYINPUT1), .ZN(new_n400));
  INV_X1    g199(.A(new_n394), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT70), .B(G134gat), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(new_n395), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G141gat), .B(G148gat), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT2), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n407), .B1(G155gat), .B2(G162gat), .ZN(new_n408));
  INV_X1    g207(.A(G155gat), .ZN(new_n409));
  INV_X1    g208(.A(G162gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI22_X1  g210(.A1(new_n406), .A2(new_n408), .B1(KEYINPUT76), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G155gat), .B(G162gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n412), .B(new_n413), .Z(new_n414));
  INV_X1    g213(.A(KEYINPUT3), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n412), .B(new_n413), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT3), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n405), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n392), .A2(new_n397), .B1(new_n403), .B2(new_n400), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(KEYINPUT4), .A3(new_n414), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n419), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n398), .A2(new_n404), .A3(new_n414), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT77), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n421), .A2(KEYINPUT77), .A3(new_n414), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n387), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n426), .B(new_n428), .C1(new_n421), .C2(new_n414), .ZN(new_n431));
  INV_X1    g230(.A(new_n420), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n427), .B1(new_n426), .B2(new_n428), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n424), .A2(new_n427), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n419), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n438), .A2(KEYINPUT5), .A3(new_n432), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n430), .A2(new_n433), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G1gat), .B(G29gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(KEYINPUT0), .ZN(new_n442));
  XOR2_X1   g241(.A(G57gat), .B(G85gat), .Z(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n444), .B(KEYINPUT85), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT39), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n434), .A2(new_n438), .A3(new_n436), .ZN(new_n449));
  NOR3_X1   g248(.A1(new_n449), .A2(KEYINPUT86), .A3(new_n420), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT86), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n424), .A2(new_n425), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT77), .B1(new_n421), .B2(new_n414), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT4), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(new_n419), .A3(new_n435), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n451), .B1(new_n455), .B2(new_n432), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n448), .B1(new_n450), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT86), .B1(new_n449), .B2(new_n420), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n455), .A2(new_n451), .A3(new_n432), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n431), .A2(new_n432), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n458), .A2(KEYINPUT39), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n461), .A3(new_n446), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT40), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n447), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n457), .A2(new_n461), .A3(KEYINPUT40), .A4(new_n446), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n465), .A2(KEYINPUT87), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(KEYINPUT87), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n386), .B(new_n464), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n417), .A2(KEYINPUT3), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n363), .B1(new_n469), .B2(KEYINPUT29), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT81), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT81), .B(new_n363), .C1(new_n469), .C2(KEYINPUT29), .ZN(new_n473));
  NAND2_X1  g272(.A1(G228gat), .A2(G233gat), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n415), .B1(new_n363), .B2(KEYINPUT29), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n474), .B1(new_n475), .B2(new_n417), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT82), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n472), .A2(KEYINPUT82), .A3(new_n473), .A4(new_n476), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n362), .A2(new_n356), .A3(KEYINPUT80), .A4(new_n360), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n481), .B(new_n350), .C1(new_n366), .C2(KEYINPUT80), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n415), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n417), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n470), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n479), .A2(new_n480), .B1(new_n474), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(G22gat), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT83), .B1(new_n486), .B2(new_n244), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT84), .ZN(new_n490));
  XNOR2_X1  g289(.A(G78gat), .B(G106gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT79), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(KEYINPUT31), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(new_n227), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n489), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n490), .B1(new_n489), .B2(new_n494), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n488), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n489), .A2(new_n494), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT84), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n489), .A2(new_n490), .A3(new_n494), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n487), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n430), .A2(new_n433), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n437), .A2(new_n439), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(new_n504), .A3(new_n444), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n505), .B(new_n506), .C1(new_n440), .C2(new_n446), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n444), .B1(new_n503), .B2(new_n504), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n507), .A2(new_n509), .A3(new_n371), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT37), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n370), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n364), .A2(new_n367), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n381), .A2(new_n513), .B1(new_n514), .B2(KEYINPUT37), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(KEYINPUT89), .A3(KEYINPUT38), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n512), .B1(new_n514), .B2(new_n380), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n355), .A2(new_n366), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n511), .B1(new_n365), .B2(new_n363), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT38), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT88), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n381), .A2(new_n513), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT88), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n525), .A2(new_n526), .A3(new_n522), .A4(new_n521), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(new_n515), .B2(new_n522), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n510), .A2(new_n517), .A3(new_n528), .A4(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n468), .A2(new_n502), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT78), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n506), .B(new_n505), .C1(new_n508), .C2(new_n533), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n440), .A2(KEYINPUT78), .A3(new_n444), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n509), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n381), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n371), .A2(new_n372), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT75), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n539), .B2(new_n384), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n536), .A2(new_n540), .A3(new_n379), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n346), .B(new_n421), .ZN(new_n542));
  INV_X1    g341(.A(G227gat), .ZN(new_n543));
  INV_X1    g342(.A(G233gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT34), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT34), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n542), .A2(new_n549), .A3(new_n546), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n346), .A2(new_n421), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n346), .A2(new_n421), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n545), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT33), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G15gat), .B(G43gat), .Z(new_n556));
  XNOR2_X1  g355(.A(G71gat), .B(G99gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n548), .B(new_n550), .C1(new_n555), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n553), .A2(KEYINPUT32), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n559), .B1(new_n553), .B2(new_n554), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n549), .B1(new_n542), .B2(new_n546), .ZN(new_n564));
  AOI211_X1 g363(.A(KEYINPUT34), .B(new_n545), .C1(new_n551), .C2(new_n552), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n560), .A2(new_n562), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n562), .B1(new_n560), .B2(new_n566), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n569));
  NOR3_X1   g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n566), .ZN(new_n571));
  NOR3_X1   g370(.A1(new_n563), .A2(new_n565), .A3(new_n564), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n561), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n560), .A2(new_n562), .A3(new_n566), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT36), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI221_X1 g374(.A(new_n532), .B1(new_n541), .B2(new_n502), .C1(new_n570), .C2(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n567), .A2(new_n568), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n502), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(new_n386), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT35), .B1(new_n507), .B2(new_n509), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n541), .A2(new_n502), .A3(new_n577), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT35), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n308), .B1(new_n576), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(KEYINPUT98), .A2(G57gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(G64gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  OR2_X1    g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT9), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G57gat), .B(G64gat), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n588), .B(new_n589), .C1(new_n593), .C2(new_n590), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n597), .B(new_n598), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G127gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n595), .B(KEYINPUT99), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n264), .B1(new_n601), .B2(KEYINPUT21), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n600), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT100), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(new_n409), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n605), .B(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n603), .A2(new_n608), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G134gat), .B(G162gat), .Z(new_n612));
  AOI21_X1  g411(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT103), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT7), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT101), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT7), .ZN(new_n619));
  AND2_X1   g418(.A1(G85gat), .A2(G92gat), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G85gat), .A2(G92gat), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(KEYINPUT101), .A3(new_n616), .ZN(new_n623));
  NAND2_X1  g422(.A1(G99gat), .A2(G106gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT8), .ZN(new_n625));
  INV_X1    g424(.A(G85gat), .ZN(new_n626));
  INV_X1    g425(.A(G92gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n623), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(KEYINPUT102), .B1(new_n621), .B2(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(G99gat), .B(G106gat), .Z(new_n631));
  NAND3_X1  g430(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n632));
  AOI22_X1  g431(.A1(KEYINPUT8), .A2(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .A4(new_n623), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n630), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n631), .B1(new_n630), .B2(new_n635), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n615), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n631), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n623), .A2(new_n625), .A3(new_n628), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n634), .B1(new_n640), .B2(new_n632), .ZN(new_n641));
  INV_X1    g440(.A(new_n635), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n630), .A2(new_n631), .A3(new_n635), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(KEYINPUT103), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n646), .A2(new_n282), .A3(new_n281), .ZN(new_n647));
  XNOR2_X1  g446(.A(G190gat), .B(G218gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n638), .A2(new_n270), .A3(new_n645), .ZN(new_n650));
  NAND3_X1  g449(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n647), .A2(new_n649), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n650), .A2(new_n651), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n655), .A2(KEYINPUT104), .A3(new_n649), .A4(new_n647), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n614), .B1(new_n657), .B2(KEYINPUT105), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n647), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n648), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n657), .B(new_n660), .C1(KEYINPUT105), .C2(new_n614), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n638), .A2(new_n645), .A3(KEYINPUT10), .A4(new_n601), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n595), .B1(new_n636), .B2(new_n637), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n643), .A2(new_n644), .A3(new_n596), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT10), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT106), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672));
  AOI211_X1 g471(.A(new_n672), .B(KEYINPUT10), .C1(new_n667), .C2(new_n668), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n666), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(G230gat), .A2(G233gat), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n675), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n667), .A2(new_n677), .A3(new_n668), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(G120gat), .B(G148gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(G176gat), .B(G204gat), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n680), .B(new_n681), .Z(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n676), .A2(new_n678), .A3(new_n682), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n611), .A2(new_n665), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n585), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n536), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(new_n250), .ZN(G1324gat));
  INV_X1    g491(.A(new_n690), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n386), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT107), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(new_n242), .ZN(new_n697));
  OR3_X1    g496(.A1(new_n694), .A2(G8gat), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n695), .ZN(new_n699));
  OAI21_X1  g498(.A(G8gat), .B1(new_n694), .B2(new_n697), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(G1325gat));
  AOI21_X1  g500(.A(G15gat), .B1(new_n693), .B2(new_n577), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT108), .B1(new_n570), .B2(new_n575), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n569), .B1(new_n567), .B2(new_n568), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n573), .A2(KEYINPUT36), .A3(new_n574), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G15gat), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT109), .Z(new_n710));
  AOI21_X1  g509(.A(new_n702), .B1(new_n693), .B2(new_n710), .ZN(G1326gat));
  NOR2_X1   g510(.A1(new_n690), .A2(new_n502), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT43), .B(G22gat), .Z(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  INV_X1    g513(.A(new_n611), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n687), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n665), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n585), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n536), .A2(G29gat), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT110), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n718), .A2(new_n722), .A3(new_n719), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n721), .A2(KEYINPUT45), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT45), .B1(new_n721), .B2(new_n723), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n579), .A2(new_n580), .B1(new_n582), .B2(KEYINPUT35), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n468), .A2(new_n502), .A3(new_n531), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n707), .B(new_n703), .C1(new_n541), .C2(new_n502), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT112), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n386), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n536), .ZN(new_n733));
  INV_X1    g532(.A(new_n502), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n708), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(new_n736), .A3(new_n532), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n728), .B1(new_n731), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n727), .B1(new_n738), .B2(new_n665), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n576), .A2(new_n584), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(KEYINPUT44), .A3(new_n664), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n279), .A2(new_n290), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n207), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n297), .A2(new_n300), .A3(KEYINPUT97), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n306), .B1(new_n305), .B2(new_n279), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT111), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n301), .A2(new_n307), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(new_n750), .A3(new_n744), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n716), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n742), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G29gat), .B1(new_n754), .B2(new_n536), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n726), .A2(new_n755), .ZN(G1328gat));
  NAND4_X1  g555(.A1(new_n739), .A2(new_n386), .A3(new_n741), .A4(new_n753), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G36gat), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n585), .A2(new_n221), .A3(new_n386), .A4(new_n717), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n758), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1329gat));
  NAND2_X1  g563(.A1(new_n585), .A2(new_n717), .ZN(new_n765));
  INV_X1    g564(.A(new_n577), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n765), .A2(G43gat), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT47), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(KEYINPUT114), .B2(new_n768), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n768), .A2(KEYINPUT114), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n739), .A2(new_n708), .A3(new_n741), .A4(new_n753), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G43gat), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n770), .B1(new_n769), .B2(new_n772), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(G1330gat));
  OAI21_X1  g574(.A(new_n227), .B1(new_n765), .B2(new_n502), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n734), .A2(G50gat), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n754), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT48), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT48), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n780), .B(new_n776), .C1(new_n754), .C2(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(G1331gat));
  INV_X1    g581(.A(new_n752), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n665), .A2(new_n611), .A3(new_n686), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n738), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n536), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g587(.A(new_n732), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT115), .ZN(new_n791));
  NOR2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n791), .B(new_n792), .ZN(G1333gat));
  INV_X1    g592(.A(G71gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n785), .A2(new_n794), .A3(new_n577), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n785), .A2(new_n708), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(new_n794), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n797), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g597(.A1(new_n785), .A2(new_n734), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g599(.A1(new_n783), .A2(new_n611), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(new_n687), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n742), .A2(new_n786), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G85gat), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n729), .A2(new_n730), .A3(KEYINPUT112), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n736), .B1(new_n735), .B2(new_n532), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n584), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(new_n664), .A3(new_n801), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n731), .A2(new_n737), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n665), .B1(new_n812), .B2(new_n584), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(KEYINPUT51), .A3(new_n801), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n786), .A2(new_n626), .A3(new_n686), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n805), .B1(new_n816), .B2(new_n817), .ZN(G1336gat));
  NOR3_X1   g617(.A1(new_n732), .A2(G92gat), .A3(new_n687), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n739), .A2(new_n386), .A3(new_n741), .A4(new_n803), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G92gat), .ZN(new_n822));
  XNOR2_X1  g621(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(new_n820), .B2(new_n822), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n824), .A2(new_n825), .ZN(G1337gat));
  NAND3_X1  g625(.A1(new_n742), .A2(new_n708), .A3(new_n803), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(G99gat), .ZN(new_n828));
  OR3_X1    g627(.A1(new_n766), .A2(G99gat), .A3(new_n687), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n828), .B1(new_n816), .B2(new_n829), .ZN(G1338gat));
  NOR2_X1   g629(.A1(new_n502), .A2(new_n687), .ZN(new_n831));
  AOI21_X1  g630(.A(G106gat), .B1(new_n815), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(G106gat), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n502), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n739), .A2(new_n741), .A3(new_n803), .A4(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n836), .A2(new_n837), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n832), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n840), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT51), .B1(new_n813), .B2(new_n801), .ZN(new_n843));
  NOR4_X1   g642(.A1(new_n738), .A2(new_n810), .A3(new_n665), .A4(new_n802), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n831), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n833), .ZN(new_n846));
  INV_X1    g645(.A(new_n839), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n841), .A2(new_n848), .ZN(G1339gat));
  OAI211_X1 g648(.A(new_n666), .B(new_n677), .C1(new_n671), .C2(new_n673), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n676), .A2(KEYINPUT54), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n674), .A2(new_n852), .A3(new_n675), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n851), .A2(KEYINPUT55), .A3(new_n683), .A4(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(new_n685), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n676), .A2(KEYINPUT54), .A3(new_n850), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n853), .A2(new_n683), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n748), .A2(new_n855), .A3(new_n751), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n288), .A2(new_n209), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n295), .A2(new_n210), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n205), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n686), .A2(new_n749), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n664), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n662), .A2(new_n749), .A3(new_n663), .A4(new_n863), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n859), .A2(new_n685), .A3(new_n854), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n715), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n689), .A2(new_n752), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n502), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT118), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n871), .A2(new_n874), .A3(new_n502), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n876), .A2(new_n786), .A3(new_n732), .A4(new_n577), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(new_n388), .A3(new_n308), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n536), .B1(new_n869), .B2(new_n870), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n879), .A2(new_n579), .ZN(new_n880));
  AOI21_X1  g679(.A(G113gat), .B1(new_n880), .B2(new_n783), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n878), .A2(new_n881), .ZN(G1340gat));
  OAI21_X1  g681(.A(G120gat), .B1(new_n877), .B2(new_n687), .ZN(new_n883));
  INV_X1    g682(.A(new_n390), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n880), .A2(new_n884), .A3(new_n686), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(G1341gat));
  OAI21_X1  g685(.A(G127gat), .B1(new_n877), .B2(new_n715), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n880), .A2(new_n395), .A3(new_n611), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1342gat));
  OAI21_X1  g688(.A(G134gat), .B1(new_n877), .B2(new_n665), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n402), .B1(KEYINPUT119), .B2(KEYINPUT56), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n880), .A2(new_n664), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n892), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n890), .A2(new_n894), .ZN(G1343gat));
  NAND2_X1  g694(.A1(new_n871), .A2(new_n734), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(KEYINPUT120), .A3(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n870), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n854), .A2(new_n685), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n636), .A2(new_n637), .A3(new_n595), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n596), .B1(new_n643), .B2(new_n644), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n670), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n672), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n669), .A2(KEYINPUT106), .A3(new_n670), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n677), .B1(new_n906), .B2(new_n666), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n682), .B1(new_n907), .B2(new_n852), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT55), .B1(new_n908), .B2(new_n851), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n900), .A2(new_n308), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n864), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n665), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n866), .A2(new_n867), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n611), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI211_X1 g713(.A(KEYINPUT57), .B(new_n734), .C1(new_n899), .C2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n502), .B1(new_n869), .B2(new_n870), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(KEYINPUT57), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n898), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n732), .A2(new_n786), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(new_n708), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(G141gat), .B1(new_n922), .B2(new_n308), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n708), .A2(new_n386), .A3(new_n502), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n924), .A2(new_n879), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n308), .A2(G141gat), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(KEYINPUT58), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n922), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n783), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n927), .B1(new_n931), .B2(G141gat), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT58), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(G1344gat));
  AOI21_X1  g733(.A(new_n897), .B1(new_n871), .B2(new_n734), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n734), .A2(new_n897), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n912), .A2(new_n937), .A3(new_n913), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n747), .A2(new_n859), .A3(new_n685), .A4(new_n854), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n664), .B1(new_n939), .B2(new_n864), .ZN(new_n940));
  OAI21_X1  g739(.A(KEYINPUT121), .B1(new_n940), .B2(new_n868), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n941), .A3(new_n715), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n689), .A2(new_n308), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n936), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n921), .ZN(new_n945));
  NOR4_X1   g744(.A1(new_n935), .A2(new_n944), .A3(new_n687), .A4(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(G148gat), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT59), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT122), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n896), .A2(KEYINPUT57), .ZN(new_n950));
  INV_X1    g749(.A(new_n944), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n950), .A2(new_n951), .A3(new_n686), .A4(new_n921), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G148gat), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT122), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT59), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n919), .A2(new_n686), .A3(new_n921), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n947), .A2(KEYINPUT59), .ZN(new_n957));
  AOI22_X1  g756(.A1(new_n949), .A2(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n925), .A2(new_n947), .A3(new_n686), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(KEYINPUT123), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n956), .A2(new_n957), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n954), .B1(new_n953), .B2(KEYINPUT59), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT59), .ZN(new_n964));
  AOI211_X1 g763(.A(KEYINPUT122), .B(new_n964), .C1(new_n952), .C2(G148gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n962), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n966), .A2(new_n967), .A3(new_n959), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n961), .A2(new_n968), .ZN(G1345gat));
  OAI21_X1  g768(.A(G155gat), .B1(new_n922), .B2(new_n715), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n925), .A2(new_n409), .A3(new_n611), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1346gat));
  AOI21_X1  g771(.A(G162gat), .B1(new_n925), .B2(new_n664), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n665), .A2(new_n410), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n973), .B1(new_n930), .B2(new_n974), .ZN(G1347gat));
  NAND2_X1  g774(.A1(new_n871), .A2(new_n536), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT124), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n578), .A2(new_n732), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g779(.A(G169gat), .B1(new_n980), .B2(new_n783), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n732), .A2(new_n786), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  AOI211_X1 g782(.A(new_n766), .B(new_n983), .C1(new_n873), .C2(new_n875), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n747), .A2(G169gat), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(G1348gat));
  AND3_X1   g785(.A1(new_n984), .A2(G176gat), .A3(new_n686), .ZN(new_n987));
  AOI21_X1  g786(.A(G176gat), .B1(new_n980), .B2(new_n686), .ZN(new_n988));
  OR2_X1    g787(.A1(new_n988), .A2(KEYINPUT125), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(KEYINPUT125), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n987), .B1(new_n989), .B2(new_n990), .ZN(G1349gat));
  NAND2_X1  g790(.A1(new_n984), .A2(new_n611), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n611), .A2(new_n310), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  AOI22_X1  g793(.A1(G183gat), .A2(new_n992), .B1(new_n980), .B2(new_n994), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT60), .ZN(new_n996));
  XNOR2_X1  g795(.A(new_n995), .B(new_n996), .ZN(G1350gat));
  NAND3_X1  g796(.A1(new_n980), .A2(new_n309), .A3(new_n664), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n984), .A2(new_n664), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(G190gat), .ZN(new_n1000));
  AND2_X1   g799(.A1(new_n1000), .A2(KEYINPUT61), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n1000), .A2(KEYINPUT61), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(G1351gat));
  NOR2_X1   g802(.A1(new_n935), .A2(new_n944), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n983), .A2(new_n708), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g805(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g806(.A(G197gat), .ZN(new_n1008));
  NOR3_X1   g807(.A1(new_n1007), .A2(new_n1008), .A3(new_n308), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n708), .A2(new_n732), .A3(new_n502), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n977), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1011), .A2(KEYINPUT126), .ZN(new_n1012));
  INV_X1    g811(.A(KEYINPUT126), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n977), .A2(new_n1013), .A3(new_n1010), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1012), .A2(new_n783), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g814(.A(new_n1009), .B1(new_n1015), .B2(new_n1008), .ZN(G1352gat));
  OR3_X1    g815(.A1(new_n1011), .A2(G204gat), .A3(new_n687), .ZN(new_n1017));
  OR2_X1    g816(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n1004), .A2(new_n686), .A3(new_n1005), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1019), .A2(G204gat), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .ZN(G1353gat));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n611), .ZN(new_n1023));
  AND3_X1   g822(.A1(new_n1023), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1024));
  AOI21_X1  g823(.A(KEYINPUT63), .B1(new_n1023), .B2(G211gat), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n611), .A2(new_n358), .ZN(new_n1027));
  OAI22_X1  g826(.A1(new_n1024), .A2(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(G1354gat));
  OAI21_X1  g827(.A(G218gat), .B1(new_n1007), .B2(new_n665), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n664), .A2(new_n359), .ZN(new_n1030));
  OAI21_X1  g829(.A(new_n1029), .B1(new_n1026), .B2(new_n1030), .ZN(G1355gat));
endmodule


