//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT78), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G125), .B(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT78), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT18), .A2(G131), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G237), .ZN(new_n202));
  INV_X1    g016(.A(G953), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G214), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n202), .A2(new_n203), .A3(G143), .A4(G214), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT88), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n201), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(new_n207), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n211), .A2(KEYINPUT88), .A3(new_n200), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n199), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT89), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT89), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n215), .B(new_n199), .C1(new_n210), .C2(new_n212), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G113), .B(G122), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n211), .A2(G131), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n206), .A2(new_n223), .A3(new_n207), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT92), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT90), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n229));
  OR3_X1    g043(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n229), .A2(G146), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(G146), .B1(new_n229), .B2(new_n230), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n228), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n230), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n196), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n229), .A2(new_n230), .A3(G146), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(KEYINPUT90), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n211), .A2(KEYINPUT17), .A3(G131), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n233), .A2(new_n237), .A3(KEYINPUT91), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n225), .A2(new_n226), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n227), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n233), .A2(new_n237), .A3(new_n238), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT91), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n217), .B(new_n220), .C1(new_n241), .C2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT93), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n242), .A2(new_n243), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n248), .A2(new_n239), .A3(new_n240), .A4(new_n227), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n249), .A2(KEYINPUT93), .A3(new_n220), .A4(new_n217), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n231), .B1(new_n221), .B2(new_n224), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT19), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n193), .A2(new_n195), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n253), .B2(new_n194), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n252), .B1(new_n255), .B2(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n217), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n220), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n251), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT20), .ZN(new_n261));
  NOR2_X1   g075(.A1(G475), .A2(G902), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n247), .A2(new_n250), .B1(new_n258), .B2(new_n257), .ZN(new_n264));
  INV_X1    g078(.A(new_n262), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT20), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n249), .A2(new_n217), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n247), .A2(new_n250), .B1(new_n258), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(G475), .B1(new_n269), .B2(G902), .ZN(new_n270));
  INV_X1    g084(.A(G902), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT96), .ZN(new_n272));
  XOR2_X1   g086(.A(G116), .B(G122), .Z(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(KEYINPUT14), .ZN(new_n274));
  INV_X1    g088(.A(G116), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT14), .A3(G122), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G107), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n272), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n276), .A2(G107), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(KEYINPUT96), .C1(new_n273), .C2(KEYINPUT14), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n205), .A2(G128), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT94), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n283), .A2(new_n205), .A3(G128), .ZN(new_n284));
  INV_X1    g098(.A(G128), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT94), .B1(new_n285), .B2(G143), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n282), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n287), .B(G134), .ZN(new_n288));
  XNOR2_X1  g102(.A(G116), .B(G122), .ZN(new_n289));
  INV_X1    g103(.A(G107), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(KEYINPUT95), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n281), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n282), .B(KEYINPUT13), .Z(new_n294));
  NOR2_X1   g108(.A1(new_n284), .A2(new_n286), .ZN(new_n295));
  OAI21_X1  g109(.A(G134), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n273), .A2(G107), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n291), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n296), .B(new_n298), .C1(G134), .C2(new_n287), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT9), .B(G234), .ZN(new_n300));
  INV_X1    g114(.A(G217), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n300), .A2(new_n301), .A3(G953), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n293), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n302), .B1(new_n293), .B2(new_n299), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n271), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT97), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G478), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(KEYINPUT15), .ZN(new_n310));
  OAI211_X1 g124(.A(KEYINPUT97), .B(new_n271), .C1(new_n304), .C2(new_n305), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n306), .A2(new_n310), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G952), .ZN(new_n316));
  AOI211_X1 g130(.A(G953), .B(new_n316), .C1(G234), .C2(G237), .ZN(new_n317));
  AOI211_X1 g131(.A(new_n271), .B(new_n203), .C1(G234), .C2(G237), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT21), .B(G898), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n267), .A2(new_n270), .A3(new_n315), .A4(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G472), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n271), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT11), .ZN(new_n326));
  INV_X1    g140(.A(G134), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(G137), .ZN(new_n328));
  INV_X1    g142(.A(G137), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT11), .A3(G134), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(G137), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G131), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n328), .A2(new_n330), .A3(new_n223), .A4(new_n331), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT68), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT0), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n285), .B1(new_n338), .B2(KEYINPUT64), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(KEYINPUT64), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(new_n285), .A3(KEYINPUT64), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n196), .A2(G143), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n205), .A2(KEYINPUT65), .A3(G146), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT65), .B1(new_n205), .B2(G146), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n205), .A2(G146), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n344), .A2(new_n348), .A3(KEYINPUT0), .A4(G128), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT66), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(G143), .B(G146), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n352), .A2(KEYINPUT66), .A3(KEYINPUT0), .A4(G128), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n343), .A2(new_n347), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n333), .A2(KEYINPUT68), .A3(new_n334), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n337), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT69), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n327), .A2(G137), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n329), .A2(G134), .ZN(new_n359));
  OAI21_X1  g173(.A(G131), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n334), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT1), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n344), .A2(new_n348), .A3(new_n362), .A4(G128), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n205), .A2(G146), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT65), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n365), .B1(new_n196), .B2(G143), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n205), .A2(KEYINPUT65), .A3(G146), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n285), .B1(new_n344), .B2(KEYINPUT1), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n363), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n357), .B1(new_n361), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n361), .A2(new_n370), .A3(new_n357), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n356), .A2(new_n372), .A3(KEYINPUT30), .A4(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT67), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT2), .B(G113), .Z(new_n376));
  XNOR2_X1  g190(.A(G116), .B(G119), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G119), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G116), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n275), .A2(G119), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT2), .B(G113), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n375), .B1(new_n378), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n376), .A2(new_n377), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(new_n383), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(KEYINPUT67), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n351), .A2(new_n353), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n347), .A2(new_n341), .A3(new_n342), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n335), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n361), .A2(new_n370), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT30), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n389), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n374), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT71), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G210), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n401), .A2(G237), .A3(G953), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n398), .B(KEYINPUT71), .ZN(new_n404));
  INV_X1    g218(.A(new_n402), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT26), .B(G101), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n403), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n407), .B1(new_n403), .B2(new_n406), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n356), .A2(new_n372), .A3(new_n373), .A4(new_n389), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT31), .B1(new_n397), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n410), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT73), .B(KEYINPUT28), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n385), .A2(new_n388), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n394), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n416), .B1(new_n411), .B2(new_n418), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n385), .A2(new_n388), .B1(new_n370), .B2(new_n361), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT28), .B1(new_n356), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n414), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n413), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n374), .A2(new_n396), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT31), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n411), .A4(new_n410), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT72), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n412), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n429), .A2(KEYINPUT72), .A3(new_n425), .A4(new_n424), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n325), .B1(new_n423), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT29), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n424), .A2(new_n414), .A3(new_n433), .A4(new_n411), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n434), .A2(new_n271), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n411), .A2(new_n418), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n415), .ZN(new_n437));
  INV_X1    g251(.A(new_n421), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n410), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n421), .B(KEYINPUT75), .ZN(new_n441));
  INV_X1    g255(.A(new_n411), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n361), .A2(new_n370), .A3(new_n357), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(new_n371), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n389), .B1(new_n444), .B2(new_n356), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT28), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n433), .B1(new_n441), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n435), .B1(new_n440), .B2(new_n447), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n432), .A2(KEYINPUT32), .B1(new_n448), .B2(G472), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT74), .B1(new_n432), .B2(KEYINPUT32), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT74), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT32), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n413), .A2(new_n422), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n428), .B2(new_n430), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n451), .B(new_n452), .C1(new_n454), .C2(new_n325), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n449), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n285), .A2(G119), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n379), .A2(G128), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT24), .B(G110), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT77), .B1(new_n379), .B2(G128), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT23), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT23), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n457), .A2(KEYINPUT77), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n463), .A2(new_n465), .A3(new_n458), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n461), .B1(new_n466), .B2(G110), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n236), .A3(new_n197), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT79), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(G110), .ZN(new_n471));
  OAI221_X1 g285(.A(new_n471), .B1(new_n459), .B2(new_n460), .C1(new_n231), .C2(new_n232), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n203), .A2(G221), .A3(G234), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT80), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT22), .B(G137), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n477), .B1(new_n470), .B2(new_n472), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n271), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT25), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g297(.A(KEYINPUT25), .B(new_n271), .C1(new_n479), .C2(new_n480), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(G217), .A2(G902), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n301), .B2(G234), .ZN(new_n487));
  XOR2_X1   g301(.A(new_n487), .B(KEYINPUT76), .Z(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n479), .A2(new_n480), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n488), .A2(G902), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G469), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT3), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n290), .A3(G104), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT82), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT82), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n499), .A2(new_n496), .A3(new_n290), .A4(G104), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n290), .A2(G104), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT3), .B1(new_n219), .B2(G107), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT81), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G101), .ZN(new_n506));
  OAI211_X1 g320(.A(KEYINPUT81), .B(KEYINPUT3), .C1(new_n219), .C2(G107), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n501), .A2(new_n505), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n219), .A2(G107), .ZN(new_n509));
  OAI21_X1  g323(.A(G101), .B1(new_n509), .B2(new_n502), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n363), .B1(new_n369), .B2(new_n352), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n370), .B1(new_n508), .B2(new_n510), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n335), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n514), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n512), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n333), .A2(KEYINPUT68), .A3(new_n334), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT68), .B1(new_n333), .B2(new_n334), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT12), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n515), .A2(KEYINPUT12), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n508), .A2(new_n510), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n370), .A2(KEYINPUT10), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT84), .B(KEYINPUT10), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n523), .A2(new_n524), .B1(new_n512), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(KEYINPUT83), .A2(G101), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n498), .A2(new_n500), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n503), .A2(new_n504), .ZN(new_n529));
  INV_X1    g343(.A(new_n502), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n507), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n527), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(KEYINPUT4), .A3(new_n508), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n501), .A2(new_n507), .A3(new_n505), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT4), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n534), .A2(KEYINPUT83), .A3(new_n535), .A4(G101), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n533), .A2(new_n354), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT85), .B1(new_n518), .B2(new_n519), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT85), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n337), .A2(new_n539), .A3(new_n355), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n526), .A2(new_n537), .A3(new_n538), .A4(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(G110), .B(G140), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n203), .A2(G227), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n521), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n518), .A2(new_n519), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n533), .A2(new_n354), .A3(new_n536), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n512), .A2(new_n525), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n508), .A2(KEYINPUT10), .A3(new_n370), .A4(new_n510), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n547), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n545), .B1(new_n552), .B2(new_n541), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n495), .B(new_n271), .C1(new_n546), .C2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n495), .A2(new_n271), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n538), .A2(new_n540), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n548), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n520), .B1(new_n513), .B2(new_n514), .ZN(new_n559));
  INV_X1    g373(.A(new_n335), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(new_n516), .B2(new_n512), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT12), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n544), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n552), .A2(new_n541), .A3(new_n545), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n554), .B(new_n556), .C1(new_n495), .C2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(G221), .B1(new_n300), .B2(G902), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G214), .B1(G237), .B2(G902), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n390), .A2(new_n391), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G125), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n368), .A2(new_n369), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n189), .A3(new_n363), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G224), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(G953), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT7), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT87), .B1(new_n575), .B2(new_n580), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT87), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n572), .A2(new_n583), .A3(new_n574), .A4(new_n579), .ZN(new_n584));
  XNOR2_X1  g398(.A(G110), .B(G122), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT8), .ZN(new_n586));
  INV_X1    g400(.A(G113), .ZN(new_n587));
  INV_X1    g401(.A(new_n380), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT5), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n377), .A2(KEYINPUT5), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n590), .A2(new_n591), .B1(new_n377), .B2(new_n376), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n508), .A2(new_n592), .A3(new_n510), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n508), .B2(new_n510), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n586), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AND4_X1   g410(.A1(new_n581), .A2(new_n582), .A3(new_n584), .A4(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n417), .A2(new_n533), .A3(new_n536), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT86), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n508), .A2(new_n592), .A3(KEYINPUT86), .A4(new_n510), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n598), .A2(new_n585), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(G902), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n585), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n417), .A2(new_n533), .A3(new_n536), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n600), .A2(new_n601), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(KEYINPUT6), .A3(new_n602), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n575), .B(new_n577), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT6), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n610), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(G210), .B1(G237), .B2(G902), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n603), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n613), .B1(new_n603), .B2(new_n612), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n570), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n569), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n323), .A2(new_n456), .A3(new_n494), .A4(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT98), .B(G101), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G3));
  OAI21_X1  g434(.A(G472), .B1(new_n454), .B2(G902), .ZN(new_n621));
  INV_X1    g435(.A(new_n432), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n623), .A2(new_n493), .A3(new_n569), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT99), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n268), .A2(new_n258), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n251), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n271), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n263), .A2(new_n266), .B1(new_n628), .B2(G475), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n570), .B(new_n321), .C1(new_n614), .C2(new_n615), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT33), .B1(new_n302), .B2(KEYINPUT100), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n304), .B2(new_n305), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n293), .A2(new_n299), .ZN(new_n633));
  INV_X1    g447(.A(new_n302), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n631), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n303), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n309), .A2(G902), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n632), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT101), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n632), .A2(new_n637), .A3(new_n642), .A4(new_n638), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n629), .A2(new_n630), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n625), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT102), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT34), .B(G104), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  NAND2_X1  g463(.A1(new_n270), .A2(KEYINPUT103), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n651), .B(G475), .C1(new_n269), .C2(G902), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n267), .A2(new_n650), .A3(new_n314), .A4(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n630), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n625), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT35), .B(G107), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  NOR2_X1   g471(.A1(new_n477), .A2(KEYINPUT36), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n473), .B(new_n658), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n485), .A2(new_n488), .B1(new_n491), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n623), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n323), .A3(new_n617), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  NAND2_X1  g478(.A1(new_n659), .A2(new_n491), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n489), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n456), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT104), .B(G900), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n317), .B1(new_n318), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n653), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n667), .A2(new_n668), .A3(new_n617), .A4(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n456), .A2(new_n617), .A3(new_n666), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n266), .A2(new_n263), .B1(new_n270), .B2(KEYINPUT103), .ZN(new_n674));
  INV_X1    g488(.A(new_n670), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n674), .A2(new_n314), .A3(new_n652), .A4(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT105), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  XOR2_X1   g493(.A(new_n670), .B(KEYINPUT39), .Z(new_n680));
  NAND3_X1  g494(.A1(new_n567), .A2(new_n568), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n681), .B(KEYINPUT40), .Z(new_n682));
  NAND2_X1  g496(.A1(new_n603), .A2(new_n612), .ZN(new_n683));
  INV_X1    g497(.A(new_n613), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n603), .A2(new_n612), .A3(new_n613), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(KEYINPUT38), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT38), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n688), .B1(new_n614), .B2(new_n615), .ZN(new_n689));
  AND4_X1   g503(.A1(new_n570), .A2(new_n660), .A3(new_n687), .A4(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n629), .A2(new_n315), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n442), .A2(new_n445), .ZN(new_n692));
  AOI21_X1  g506(.A(G902), .B1(new_n692), .B2(new_n414), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n410), .B1(new_n397), .B2(new_n442), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n324), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n432), .B2(KEYINPUT32), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n450), .A2(new_n696), .A3(new_n455), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n682), .A2(new_n690), .A3(new_n691), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  AOI211_X1 g513(.A(new_n670), .B(new_n644), .C1(new_n267), .C2(new_n270), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n456), .A3(new_n617), .A4(new_n666), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  NOR2_X1   g516(.A1(new_n546), .A2(new_n553), .ZN(new_n703));
  OAI21_X1  g517(.A(G469), .B1(new_n703), .B2(G902), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n554), .ZN(new_n705));
  INV_X1    g519(.A(new_n568), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n645), .A2(new_n456), .A3(new_n494), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT41), .B(G113), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G15));
  NAND4_X1  g524(.A1(new_n654), .A2(new_n456), .A3(new_n494), .A4(new_n707), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  NOR3_X1   g526(.A1(new_n616), .A2(new_n706), .A3(new_n705), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n323), .A2(new_n713), .A3(new_n456), .A4(new_n666), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT106), .B(G119), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G21));
  NAND2_X1  g530(.A1(new_n423), .A2(new_n431), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n324), .B1(new_n717), .B2(new_n271), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n410), .B1(new_n441), .B2(new_n446), .ZN(new_n719));
  INV_X1    g533(.A(new_n413), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n325), .B1(new_n721), .B2(new_n431), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n493), .A2(new_n718), .A3(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n629), .A2(new_n616), .A3(new_n315), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n723), .A2(new_n724), .A3(new_n321), .A4(new_n707), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NOR3_X1   g540(.A1(new_n660), .A2(new_n718), .A3(new_n722), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n700), .A2(new_n727), .A3(new_n713), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G125), .ZN(G27));
  INV_X1    g543(.A(KEYINPUT109), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n564), .B2(new_n565), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n565), .A2(new_n731), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n732), .A2(new_n734), .A3(new_n495), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n554), .A2(new_n556), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT108), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n547), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n526), .B2(new_n537), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n544), .B1(new_n558), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n521), .A2(new_n541), .A3(new_n545), .ZN(new_n741));
  AOI21_X1  g555(.A(G902), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n555), .B1(new_n742), .B2(new_n495), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n552), .A2(new_n541), .A3(new_n545), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n545), .B1(new_n521), .B2(new_n541), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT107), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(G469), .A3(new_n733), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n743), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n706), .B1(new_n737), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n570), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n614), .A2(new_n615), .A3(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n750), .A2(new_n456), .A3(new_n494), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n267), .A2(new_n270), .ZN(new_n754));
  INV_X1    g568(.A(new_n644), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n755), .A3(new_n675), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n730), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n456), .A2(new_n494), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n743), .A2(new_n747), .A3(new_n748), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n748), .B1(new_n743), .B2(new_n747), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n752), .B(new_n568), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n758), .A2(new_n762), .A3(KEYINPUT109), .A4(new_n700), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT42), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n757), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n432), .A2(KEYINPUT32), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT110), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n622), .A2(new_n452), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n448), .A2(G472), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n432), .A2(new_n770), .A3(KEYINPUT32), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n767), .A2(new_n768), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n494), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n773), .A2(new_n764), .A3(new_n761), .A4(new_n756), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n765), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G131), .ZN(G33));
  NOR2_X1   g591(.A1(new_n753), .A2(new_n676), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n327), .ZN(G36));
  NAND3_X1  g593(.A1(new_n685), .A2(new_n570), .A3(new_n686), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n623), .A2(new_n666), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(KEYINPUT112), .Z(new_n782));
  INV_X1    g596(.A(KEYINPUT43), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n754), .B2(new_n644), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n629), .A2(KEYINPUT43), .A3(new_n755), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n780), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n746), .A2(KEYINPUT45), .A3(new_n733), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n495), .B1(new_n566), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n555), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  OR3_X1    g607(.A1(new_n793), .A2(KEYINPUT111), .A3(KEYINPUT46), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT111), .B1(new_n793), .B2(KEYINPUT46), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(KEYINPUT46), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n794), .A2(new_n554), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n797), .A2(new_n568), .A3(new_n680), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n789), .B(new_n798), .C1(new_n788), .C2(new_n787), .ZN(new_n799));
  XOR2_X1   g613(.A(KEYINPUT113), .B(G137), .Z(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(G39));
  NOR2_X1   g615(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n797), .B2(new_n568), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n802), .ZN(new_n805));
  NAND2_X1  g619(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n797), .A2(new_n568), .A3(new_n807), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n756), .A2(new_n456), .A3(new_n494), .A4(new_n780), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n804), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  AND2_X1   g625(.A1(new_n705), .A2(KEYINPUT49), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n755), .A2(new_n570), .A3(new_n568), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n705), .A2(KEYINPUT49), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n812), .A2(new_n813), .A3(new_n814), .A4(new_n493), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n697), .B1(new_n687), .B2(new_n689), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n629), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n317), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n697), .A2(new_n493), .A3(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n780), .A2(new_n705), .A3(new_n706), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n821), .A2(new_n629), .A3(new_n644), .A4(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT119), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n820), .B1(new_n784), .B2(new_n785), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(new_n826), .A3(new_n822), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n826), .B1(new_n825), .B2(new_n822), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n727), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n707), .A2(new_n751), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n687), .B2(new_n689), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n825), .A2(new_n832), .A3(new_n723), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT50), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n825), .A2(new_n832), .A3(KEYINPUT50), .A4(new_n723), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n824), .A2(new_n830), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n705), .A2(new_n568), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n804), .B2(new_n808), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n825), .A2(new_n723), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n752), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n838), .A2(new_n839), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n824), .A2(new_n830), .A3(KEYINPUT120), .A4(new_n837), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n819), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n821), .A2(new_n754), .A3(new_n755), .A4(new_n822), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(G952), .A3(new_n203), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n713), .B2(new_n843), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT48), .ZN(new_n852));
  INV_X1    g666(.A(new_n829), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n827), .ZN(new_n854));
  INV_X1    g668(.A(new_n773), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI211_X1 g670(.A(KEYINPUT48), .B(new_n773), .C1(new_n853), .C2(new_n827), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT51), .B1(new_n841), .B2(new_n844), .ZN(new_n858));
  OAI221_X1 g672(.A(new_n851), .B1(new_n856), .B2(new_n857), .C1(new_n858), .C2(new_n838), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT121), .B1(new_n848), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n838), .A2(new_n839), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n842), .A2(new_n845), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n847), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n818), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n858), .A2(new_n838), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n851), .B1(new_n856), .B2(new_n857), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n860), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n666), .A2(new_n670), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n724), .A2(new_n750), .A3(new_n871), .A4(new_n697), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n872), .A2(new_n701), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n678), .A2(new_n728), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n872), .A2(new_n701), .A3(KEYINPUT52), .ZN(new_n877));
  AND4_X1   g691(.A1(KEYINPUT115), .A2(new_n678), .A3(new_n877), .A4(new_n728), .ZN(new_n878));
  INV_X1    g692(.A(new_n728), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n672), .B2(new_n677), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT115), .B1(new_n880), .B2(new_n877), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n876), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n711), .A2(new_n708), .A3(new_n618), .A4(new_n662), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n700), .A2(new_n727), .A3(new_n750), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n267), .A2(new_n650), .A3(new_n652), .ZN(new_n886));
  AND4_X1   g700(.A1(new_n568), .A2(new_n567), .A3(new_n315), .A4(new_n675), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n456), .A2(new_n886), .A3(new_n887), .A4(new_n666), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n780), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n778), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n629), .A2(new_n314), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n629), .B2(new_n644), .ZN(new_n892));
  INV_X1    g706(.A(new_n630), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n624), .A3(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n894), .A2(new_n714), .A3(new_n725), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n884), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n456), .A2(new_n494), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n897), .A2(new_n761), .A3(new_n756), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT42), .B1(new_n898), .B2(KEYINPUT109), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n774), .B1(new_n899), .B2(new_n757), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT53), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n896), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n882), .A2(new_n902), .ZN(new_n903));
  AOI22_X1  g717(.A1(new_n874), .A2(new_n875), .B1(new_n880), .B2(new_n877), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n894), .A2(new_n714), .A3(new_n725), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n883), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n776), .A2(new_n906), .A3(new_n890), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n901), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n903), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n896), .A2(new_n900), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT53), .B1(new_n882), .B2(new_n911), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n904), .A2(new_n907), .A3(new_n901), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(KEYINPUT116), .B(new_n910), .C1(new_n914), .C2(new_n909), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n910), .A2(KEYINPUT116), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n870), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(G952), .A2(G953), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n817), .B1(new_n917), .B2(new_n918), .ZN(G75));
  NOR2_X1   g733(.A1(new_n203), .A2(G952), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n903), .A2(new_n908), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(G210), .A3(G902), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n608), .A2(new_n611), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(new_n609), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT55), .Z(new_n927));
  OR2_X1    g741(.A1(new_n927), .A2(KEYINPUT56), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n921), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT56), .B1(new_n923), .B2(KEYINPUT122), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(KEYINPUT122), .B2(new_n923), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n929), .B1(new_n931), .B2(new_n927), .ZN(G51));
  NAND2_X1  g746(.A1(new_n790), .A2(new_n792), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT123), .ZN(new_n934));
  AOI211_X1 g748(.A(new_n271), .B(new_n934), .C1(new_n903), .C2(new_n908), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n555), .B(KEYINPUT57), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n903), .A2(new_n909), .A3(new_n908), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n909), .B1(new_n903), .B2(new_n908), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n703), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT124), .B1(new_n941), .B2(new_n920), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n776), .A2(new_n906), .A3(KEYINPUT53), .A4(new_n890), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n880), .A2(new_n877), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT115), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n880), .A2(KEYINPUT115), .A3(new_n877), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n944), .B1(new_n949), .B2(new_n876), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n876), .A2(new_n945), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT53), .B1(new_n951), .B2(new_n911), .ZN(new_n952));
  OAI21_X1  g766(.A(KEYINPUT54), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n910), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n703), .B1(new_n954), .B2(new_n936), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n943), .B(new_n921), .C1(new_n955), .C2(new_n935), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n942), .A2(new_n956), .ZN(G54));
  AND4_X1   g771(.A1(KEYINPUT58), .A2(new_n922), .A3(G475), .A4(G902), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n921), .B1(new_n958), .B2(new_n260), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n260), .B2(new_n958), .ZN(G60));
  INV_X1    g774(.A(new_n954), .ZN(new_n961));
  XNOR2_X1  g775(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n309), .A2(new_n271), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n632), .A2(new_n637), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n921), .B1(new_n961), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n915), .A2(new_n916), .A3(new_n964), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n632), .A2(new_n637), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(G63));
  XNOR2_X1  g783(.A(new_n486), .B(KEYINPUT60), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n903), .B2(new_n908), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n659), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n972), .B(new_n921), .C1(new_n490), .C2(new_n971), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(G66));
  OAI21_X1  g789(.A(G953), .B1(new_n319), .B2(new_n576), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n906), .B2(G953), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n925), .B1(G898), .B2(new_n203), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT126), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n977), .B(new_n979), .ZN(G69));
  INV_X1    g794(.A(new_n394), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n374), .B1(KEYINPUT30), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(new_n255), .ZN(new_n983));
  INV_X1    g797(.A(G900), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n983), .B1(new_n984), .B2(new_n203), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n855), .A2(new_n724), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n778), .B1(new_n798), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n799), .A2(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n880), .A2(new_n701), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n989), .A2(new_n810), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n988), .A2(new_n776), .A3(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n985), .B1(new_n992), .B2(new_n203), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n983), .B(KEYINPUT127), .Z(new_n994));
  NOR2_X1   g808(.A1(new_n681), .A2(new_n780), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n758), .A2(new_n892), .A3(new_n995), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n799), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n989), .A2(new_n698), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n997), .A2(new_n999), .A3(new_n810), .A4(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n994), .B1(new_n1001), .B2(new_n203), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n203), .B1(G227), .B2(G900), .ZN(new_n1003));
  OR3_X1    g817(.A1(new_n993), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1003), .B1(new_n993), .B2(new_n1002), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  INV_X1    g822(.A(new_n906), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1008), .B1(new_n991), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n397), .A2(new_n442), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n414), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n920), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1012), .A2(new_n694), .A3(new_n1008), .ZN(new_n1015));
  OR2_X1    g829(.A1(new_n914), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1008), .B1(new_n1001), .B2(new_n1009), .ZN(new_n1017));
  INV_X1    g831(.A(new_n694), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AND3_X1   g833(.A1(new_n1014), .A2(new_n1016), .A3(new_n1019), .ZN(G57));
endmodule


