//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G228gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n210));
  OR2_X1    g009(.A1(G197gat), .A2(G204gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G197gat), .A2(G204gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n209), .B1(new_n213), .B2(KEYINPUT72), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT72), .ZN(new_n215));
  XOR2_X1   g014(.A(G197gat), .B(G204gat), .Z(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(new_n210), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(KEYINPUT72), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n214), .B1(new_n219), .B2(new_n209), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n208), .B1(new_n220), .B2(KEYINPUT29), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n222));
  AND2_X1   g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT77), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT77), .ZN(new_n225));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT76), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(KEYINPUT2), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT2), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(KEYINPUT76), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n225), .B(new_n226), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G141gat), .B(G148gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n224), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G155gat), .ZN(new_n235));
  INV_X1    g034(.A(G162gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n226), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(G155gat), .A2(G162gat), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT80), .B1(new_n223), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n237), .A2(new_n242), .A3(new_n226), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n226), .A2(KEYINPUT2), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n241), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G141gat), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT79), .B1(new_n246), .B2(G148gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT79), .ZN(new_n248));
  INV_X1    g047(.A(G148gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n249), .A3(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT78), .B(G141gat), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n247), .B(new_n250), .C1(new_n251), .C2(new_n249), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n234), .A2(new_n239), .B1(new_n245), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n207), .B1(new_n221), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT29), .B1(new_n253), .B2(new_n208), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n220), .B1(new_n256), .B2(KEYINPUT85), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n229), .A2(KEYINPUT76), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n227), .A2(KEYINPUT2), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n223), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n233), .B1(new_n260), .B2(new_n225), .ZN(new_n261));
  NOR3_X1   g060(.A1(new_n222), .A2(KEYINPUT77), .A3(new_n223), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n239), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n252), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(new_n208), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT29), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n255), .B1(new_n257), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT86), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT86), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n255), .B(new_n272), .C1(new_n257), .C2(new_n269), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n207), .B(KEYINPUT84), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n221), .A2(new_n254), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n267), .A2(new_n220), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n206), .B1(new_n274), .B2(new_n280), .ZN(new_n281));
  AOI211_X1 g080(.A(G22gat), .B(new_n279), .C1(new_n271), .C2(new_n273), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n205), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n273), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n256), .A2(KEYINPUT85), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n268), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(new_n220), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n272), .B1(new_n287), .B2(new_n255), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n280), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G22gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n206), .A3(new_n280), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(new_n204), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n294));
  NAND2_X1  g093(.A1(G225gat), .A2(G233gat), .ZN(new_n295));
  INV_X1    g094(.A(G120gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G113gat), .ZN(new_n297));
  INV_X1    g096(.A(G113gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G120gat), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT1), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT67), .B(G134gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G127gat), .ZN(new_n303));
  INV_X1    g102(.A(G127gat), .ZN(new_n304));
  INV_X1    g103(.A(G134gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n308));
  XNOR2_X1  g107(.A(G127gat), .B(G134gat), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n300), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n308), .B1(new_n300), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n307), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n232), .B1(new_n313), .B2(KEYINPUT77), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n238), .B1(new_n314), .B2(new_n231), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n238), .A2(KEYINPUT80), .B1(KEYINPUT2), .B2(new_n226), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n252), .A2(new_n316), .A3(new_n243), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n312), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n297), .A2(new_n299), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n309), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT68), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n300), .A2(new_n308), .A3(new_n309), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n263), .A2(new_n324), .A3(new_n264), .A4(new_n307), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n295), .B1(new_n318), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n294), .B1(new_n326), .B2(KEYINPUT81), .ZN(new_n327));
  INV_X1    g126(.A(new_n295), .ZN(new_n328));
  AND4_X1   g127(.A1(new_n263), .A2(new_n324), .A3(new_n264), .A4(new_n307), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n263), .A2(new_n264), .B1(new_n324), .B2(new_n307), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT81), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT3), .B1(new_n315), .B2(new_n317), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(new_n265), .A3(new_n312), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n325), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n300), .B1(new_n304), .B2(new_n305), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n322), .A2(new_n323), .B1(new_n338), .B2(new_n303), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(new_n253), .A3(KEYINPUT4), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n335), .A2(new_n295), .A3(new_n337), .A4(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n327), .A2(new_n333), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G1gat), .B(G29gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n343), .B(KEYINPUT0), .ZN(new_n344));
  XNOR2_X1  g143(.A(G57gat), .B(G85gat), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n344), .B(new_n345), .Z(new_n346));
  AND2_X1   g145(.A1(new_n337), .A2(new_n340), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n347), .A2(new_n294), .A3(new_n295), .A4(new_n335), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n342), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT6), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n346), .B1(new_n342), .B2(new_n348), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT83), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n354), .A3(KEYINPUT6), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n342), .A2(new_n348), .ZN(new_n356));
  INV_X1    g155(.A(new_n346), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(KEYINPUT6), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT83), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n353), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n293), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT34), .ZN(new_n362));
  NAND2_X1  g161(.A1(G227gat), .A2(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT24), .ZN(new_n364));
  INV_X1    g163(.A(G183gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G190gat), .ZN(new_n366));
  INV_X1    g165(.A(G190gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G183gat), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n364), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(G183gat), .A3(G190gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT64), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G169gat), .ZN(new_n373));
  INV_X1    g172(.A(G176gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT23), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT65), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n379));
  INV_X1    g178(.A(new_n378), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT23), .B1(new_n373), .B2(new_n374), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n377), .A2(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT64), .ZN(new_n383));
  XNOR2_X1  g182(.A(G183gat), .B(G190gat), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n383), .B(new_n370), .C1(new_n384), .C2(new_n364), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n372), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n381), .A2(new_n380), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n389), .A2(KEYINPUT25), .A3(new_n375), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n370), .B1(new_n384), .B2(new_n364), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n378), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n378), .A2(KEYINPUT26), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n373), .A2(new_n374), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT28), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT27), .B(G183gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(KEYINPUT66), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT27), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT66), .B1(new_n402), .B2(G183gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n367), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n399), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n400), .A2(KEYINPUT28), .A3(new_n367), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n398), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n312), .B1(new_n394), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n392), .B1(new_n386), .B2(new_n387), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n410), .A2(new_n339), .A3(new_n407), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n362), .B(new_n363), .C1(new_n409), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT70), .ZN(new_n413));
  INV_X1    g212(.A(new_n363), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n394), .A2(new_n312), .A3(new_n408), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n339), .B1(new_n410), .B2(new_n407), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT70), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n418), .A3(new_n362), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n363), .B1(new_n409), .B2(new_n411), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT34), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n413), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n415), .A2(new_n414), .A3(new_n416), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424));
  XNOR2_X1  g223(.A(G15gat), .B(G43gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G71gat), .B(G99gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n423), .B(KEYINPUT32), .C1(new_n424), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n423), .A2(KEYINPUT32), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT69), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT69), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n423), .A2(new_n431), .A3(KEYINPUT32), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n427), .B1(new_n423), .B2(new_n424), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n422), .A2(new_n428), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n418), .B1(new_n417), .B2(new_n362), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n417), .A2(new_n362), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n434), .A2(new_n428), .B1(new_n438), .B2(new_n419), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n220), .ZN(new_n441));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n442), .B(KEYINPUT73), .Z(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n410), .B2(new_n407), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT74), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT74), .B(new_n443), .C1(new_n410), .C2(new_n407), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n266), .B1(new_n410), .B2(new_n407), .ZN(new_n449));
  INV_X1    g248(.A(new_n443), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n441), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n441), .A3(new_n444), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT75), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT75), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n446), .A2(new_n447), .B1(new_n450), .B2(new_n449), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n456), .B(new_n453), .C1(new_n457), .C2(new_n441), .ZN(new_n458));
  XNOR2_X1  g257(.A(G8gat), .B(G36gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(G64gat), .B(G92gat), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n459), .B(new_n460), .Z(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n455), .A2(new_n458), .A3(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n453), .B(new_n461), .C1(new_n457), .C2(new_n441), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n452), .A2(new_n454), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(KEYINPUT30), .A3(new_n461), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n463), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n440), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n361), .A2(new_n471), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n281), .A2(new_n282), .A3(new_n205), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n204), .B1(new_n290), .B2(new_n291), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n440), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n350), .B(new_n349), .C1(new_n352), .C2(KEYINPUT82), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n356), .A2(KEYINPUT82), .A3(new_n357), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n355), .B(new_n359), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n469), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT35), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n472), .B1(KEYINPUT89), .B2(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n293), .A2(new_n478), .A3(new_n469), .A4(new_n440), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT89), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT35), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n295), .B1(new_n347), .B2(new_n335), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT39), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n346), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n318), .A2(new_n295), .A3(new_n325), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT39), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT87), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n352), .B1(new_n492), .B2(KEYINPUT40), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n463), .A2(new_n466), .A3(new_n468), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n493), .B(new_n494), .C1(KEYINPUT40), .C2(new_n492), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT38), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT37), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n467), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n455), .A2(KEYINPUT37), .A3(new_n458), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n462), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT88), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n500), .A2(KEYINPUT88), .A3(new_n462), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n496), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n359), .A2(new_n355), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n461), .A2(KEYINPUT38), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n457), .A2(new_n220), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n451), .A2(new_n444), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n220), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT37), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n498), .B(new_n507), .C1(new_n508), .C2(new_n511), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n506), .A2(new_n353), .A3(new_n464), .A4(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n293), .B(new_n495), .C1(new_n505), .C2(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n473), .A2(new_n474), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n479), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT71), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n517), .B1(new_n440), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n434), .A2(new_n428), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n438), .A2(new_n419), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n522), .A2(KEYINPUT71), .A3(KEYINPUT36), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n516), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n481), .A2(new_n484), .B1(new_n514), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G43gat), .B(G50gat), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n527), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n528));
  NOR3_X1   g327(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT90), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  OAI221_X1 g331(.A(new_n528), .B1(KEYINPUT15), .B2(new_n527), .C1(new_n530), .C2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G29gat), .ZN(new_n534));
  INV_X1    g333(.A(G36gat), .ZN(new_n535));
  OAI22_X1  g334(.A1(new_n532), .A2(new_n529), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(KEYINPUT15), .A3(new_n527), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G85gat), .A2(G92gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542));
  INV_X1    g341(.A(G85gat), .ZN(new_n543));
  INV_X1    g342(.A(G92gat), .ZN(new_n544));
  AOI22_X1  g343(.A1(KEYINPUT8), .A2(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G99gat), .B(G106gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n526), .B1(new_n539), .B2(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT95), .Z(new_n551));
  XNOR2_X1  g350(.A(G190gat), .B(G218gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT17), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n548), .B(KEYINPUT94), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n551), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT93), .ZN(new_n559));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n559), .B(new_n560), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n553), .B1(new_n551), .B2(new_n556), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(KEYINPUT97), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(KEYINPUT97), .B2(new_n563), .ZN(new_n565));
  INV_X1    g364(.A(new_n561), .ZN(new_n566));
  INV_X1    g365(.A(new_n557), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n566), .B1(new_n567), .B2(new_n563), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n568), .A2(KEYINPUT96), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(KEYINPUT96), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n565), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G64gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(G57gat), .ZN(new_n574));
  INV_X1    g373(.A(G57gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(G64gat), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT9), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G71gat), .A2(G78gat), .ZN(new_n578));
  OR2_X1    g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT91), .B1(new_n573), .B2(G57gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT91), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n575), .A3(G64gat), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n581), .B(new_n583), .C1(new_n575), .C2(G64gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT9), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n578), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(KEYINPUT21), .ZN(new_n591));
  AND2_X1   g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(G127gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(G15gat), .B(G22gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT16), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n595), .B1(new_n596), .B2(G1gat), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(G1gat), .B2(new_n595), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G8gat), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n599), .B1(new_n590), .B2(KEYINPUT21), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n594), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G155gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n601), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n549), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n548), .A2(new_n588), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n613), .A2(KEYINPUT98), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(KEYINPUT98), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n549), .A2(new_n612), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n614), .A2(new_n615), .B1(new_n590), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G230gat), .A2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT99), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT100), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n590), .ZN(new_n621));
  INV_X1    g420(.A(new_n615), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n613), .A2(KEYINPUT98), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n625));
  INV_X1    g424(.A(new_n619), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n609), .A2(new_n610), .ZN(new_n628));
  INV_X1    g427(.A(new_n618), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n620), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n624), .A2(new_n618), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(new_n630), .A3(new_n634), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n572), .A2(new_n608), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n599), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n554), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n538), .A2(new_n599), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G229gat), .A2(G233gat), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(KEYINPUT18), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n538), .B(new_n599), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n646), .B(KEYINPUT13), .Z(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n643), .A2(new_n646), .A3(new_n644), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT18), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n647), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G113gat), .B(G141gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G197gat), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT11), .B(G169gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT12), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n654), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n525), .A2(new_n641), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n478), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT101), .B(G1gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1324gat));
  XOR2_X1   g465(.A(KEYINPUT16), .B(G8gat), .Z(new_n667));
  NAND3_X1  g466(.A1(new_n662), .A2(new_n494), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n662), .ZN(new_n669));
  OAI21_X1  g468(.A(G8gat), .B1(new_n669), .B2(new_n469), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n668), .ZN(new_n671));
  MUX2_X1   g470(.A(new_n668), .B(new_n671), .S(KEYINPUT42), .Z(G1325gat));
  AND2_X1   g471(.A1(new_n523), .A2(new_n519), .ZN(new_n673));
  OAI21_X1  g472(.A(G15gat), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n522), .A2(G15gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n669), .B2(new_n675), .ZN(G1326gat));
  NAND2_X1  g475(.A1(new_n662), .A2(new_n515), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT43), .B(G22gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NOR3_X1   g478(.A1(new_n608), .A2(new_n661), .A3(new_n639), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n525), .A2(new_n572), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n534), .A3(new_n663), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT45), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT35), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n483), .B1(new_n482), .B2(KEYINPUT35), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n687), .A2(new_n688), .A3(new_n472), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n516), .A2(new_n519), .A3(new_n523), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n503), .A2(new_n504), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT38), .ZN(new_n692));
  INV_X1    g491(.A(new_n513), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n495), .A2(new_n293), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n690), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n571), .B(new_n686), .C1(new_n689), .C2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n480), .A2(KEYINPUT89), .ZN(new_n701));
  INV_X1    g500(.A(new_n472), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n484), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n513), .B1(new_n691), .B2(KEYINPUT38), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n673), .B(new_n516), .C1(new_n704), .C2(new_n695), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n572), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(KEYINPUT104), .A3(new_n686), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n700), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n706), .B2(new_n710), .ZN(new_n711));
  OAI211_X1 g510(.A(KEYINPUT102), .B(KEYINPUT44), .C1(new_n525), .C2(new_n572), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(new_n478), .A3(new_n681), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n684), .B1(new_n715), .B2(new_n534), .ZN(G1328gat));
  NAND3_X1  g515(.A1(new_n682), .A2(new_n535), .A3(new_n494), .ZN(new_n717));
  AND2_X1   g516(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n718));
  NOR2_X1   g517(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n714), .A2(new_n469), .A3(new_n681), .ZN(new_n721));
  OAI221_X1 g520(.A(new_n720), .B1(new_n718), .B2(new_n717), .C1(new_n721), .C2(new_n535), .ZN(G1329gat));
  NOR3_X1   g521(.A1(new_n714), .A2(new_n673), .A3(new_n681), .ZN(new_n723));
  INV_X1    g522(.A(G43gat), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT106), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n682), .A2(new_n724), .A3(new_n440), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n723), .B2(new_n724), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n725), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n729), .A2(new_n730), .ZN(G1330gat));
  INV_X1    g530(.A(new_n525), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n608), .A2(new_n639), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n572), .A2(G50gat), .A3(new_n293), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n732), .A2(new_n660), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n714), .A2(new_n293), .A3(new_n681), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G50gat), .B1(new_n736), .B2(new_n737), .ZN(new_n739));
  OAI211_X1 g538(.A(KEYINPUT48), .B(new_n735), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(G50gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n735), .B1(new_n736), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n742), .A2(KEYINPUT107), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT107), .B1(new_n742), .B2(new_n743), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n740), .B1(new_n744), .B2(new_n745), .ZN(G1331gat));
  INV_X1    g545(.A(new_n608), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n747), .A2(new_n660), .A3(new_n571), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n639), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n478), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(new_n575), .ZN(G1332gat));
  XOR2_X1   g550(.A(new_n749), .B(KEYINPUT109), .Z(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n494), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n754));
  XOR2_X1   g553(.A(KEYINPUT49), .B(G64gat), .Z(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n753), .B2(new_n755), .ZN(G1333gat));
  NOR3_X1   g555(.A1(new_n749), .A2(G71gat), .A3(new_n522), .ZN(new_n757));
  INV_X1    g556(.A(new_n673), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n752), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n757), .B1(new_n759), .B2(G71gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n752), .A2(new_n515), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n608), .A2(new_n660), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n706), .A2(KEYINPUT51), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT51), .B1(new_n706), .B2(new_n764), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  MUX2_X1   g566(.A(new_n767), .B(new_n766), .S(KEYINPUT110), .Z(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n640), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n769), .A2(new_n543), .A3(new_n663), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n764), .A2(new_n639), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n708), .B2(new_n713), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773), .B2(new_n478), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n770), .A2(new_n774), .ZN(G1336gat));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n639), .A2(new_n544), .A3(new_n494), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n773), .A2(new_n469), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n779));
  OAI21_X1  g578(.A(G92gat), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n773), .A2(KEYINPUT111), .A3(new_n469), .ZN(new_n781));
  OAI221_X1 g580(.A(new_n776), .B1(new_n768), .B2(new_n777), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n778), .A2(new_n544), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n777), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT52), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(G1337gat));
  INV_X1    g585(.A(G99gat), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n769), .A2(new_n787), .A3(new_n440), .ZN(new_n788));
  OAI21_X1  g587(.A(G99gat), .B1(new_n773), .B2(new_n673), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1338gat));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  AOI211_X1 g590(.A(new_n293), .B(new_n771), .C1(new_n708), .C2(new_n713), .ZN(new_n792));
  INV_X1    g591(.A(G106gat), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n640), .A2(G106gat), .A3(new_n293), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI221_X1 g594(.A(new_n791), .B1(new_n792), .B2(new_n793), .C1(new_n768), .C2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n794), .B1(new_n765), .B2(new_n766), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n793), .B1(new_n772), .B2(new_n515), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n792), .A2(KEYINPUT112), .A3(new_n793), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n797), .B(KEYINPUT53), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT112), .B1(new_n792), .B2(new_n793), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n772), .A2(new_n515), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(new_n800), .A3(G106gat), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(new_n807), .A3(new_n798), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n797), .B1(new_n808), .B2(KEYINPUT53), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n796), .B1(new_n804), .B2(new_n809), .ZN(G1339gat));
  INV_X1    g609(.A(new_n638), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n619), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n637), .A2(KEYINPUT54), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n635), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT54), .B1(new_n620), .B2(new_n627), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n811), .B1(new_n816), .B2(KEYINPUT55), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n654), .A2(new_n659), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n645), .A2(new_n646), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n648), .A2(new_n649), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n818), .B1(new_n658), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n814), .B2(new_n815), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n817), .A2(new_n571), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n620), .A2(new_n627), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n827), .B1(new_n624), .B2(new_n618), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n634), .B1(new_n829), .B2(new_n812), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n661), .B1(new_n831), .B2(new_n823), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n832), .A2(new_n817), .B1(new_n639), .B2(new_n822), .ZN(new_n833));
  OAI211_X1 g632(.A(KEYINPUT114), .B(new_n825), .C1(new_n833), .C2(new_n571), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n828), .A2(KEYINPUT55), .A3(new_n830), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n836), .A2(new_n824), .A3(new_n660), .A4(new_n638), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n639), .A2(new_n822), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n571), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n571), .A2(new_n824), .A3(new_n822), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n836), .A2(new_n638), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n835), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n834), .A2(new_n843), .A3(new_n747), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n572), .A2(new_n661), .A3(new_n608), .A4(new_n640), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n293), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n522), .B1(new_n847), .B2(KEYINPUT115), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n478), .A2(new_n494), .ZN(new_n849));
  AOI211_X1 g648(.A(KEYINPUT115), .B(new_n515), .C1(new_n844), .C2(new_n845), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n852), .A2(new_n298), .A3(new_n661), .ZN(new_n853));
  INV_X1    g652(.A(new_n475), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n846), .A2(new_n663), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n855), .B(new_n856), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(new_n469), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n660), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n853), .B1(new_n859), .B2(new_n298), .ZN(G1340gat));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n296), .A3(new_n639), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n848), .A2(new_n639), .A3(new_n849), .A4(new_n851), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT117), .B1(new_n862), .B2(G120gat), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n862), .A2(KEYINPUT117), .A3(G120gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(G1341gat));
  NAND3_X1  g664(.A1(new_n858), .A2(new_n304), .A3(new_n608), .ZN(new_n866));
  OAI21_X1  g665(.A(G127gat), .B1(new_n852), .B2(new_n747), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1342gat));
  NOR2_X1   g667(.A1(new_n572), .A2(new_n302), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n857), .A2(new_n469), .A3(new_n869), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT56), .ZN(new_n871));
  OAI21_X1  g670(.A(G134gat), .B1(new_n852), .B2(new_n572), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(KEYINPUT56), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(G1343gat));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  INV_X1    g674(.A(new_n845), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n837), .A2(new_n877), .A3(new_n838), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n572), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n877), .B1(new_n837), .B2(new_n838), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n825), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n876), .B1(new_n881), .B2(new_n747), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT57), .B1(new_n882), .B2(new_n293), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n846), .A2(new_n884), .A3(new_n515), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n673), .A2(new_n849), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n883), .A2(new_n885), .A3(new_n660), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n251), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n846), .A2(KEYINPUT119), .A3(new_n663), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n758), .A2(new_n293), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n478), .B1(new_n844), .B2(new_n845), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(KEYINPUT119), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n889), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n846), .A2(new_n663), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n891), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n899), .B1(new_n893), .B2(KEYINPUT119), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n898), .A2(new_n900), .A3(KEYINPUT120), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n895), .A2(new_n469), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n660), .A2(new_n246), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n875), .B(new_n888), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n898), .A2(new_n900), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n660), .A2(new_n246), .A3(new_n469), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n888), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT58), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n904), .A2(new_n908), .ZN(G1344gat));
  NAND4_X1  g708(.A1(new_n895), .A2(new_n469), .A3(new_n639), .A4(new_n901), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT59), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n249), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n883), .A2(new_n885), .A3(new_n886), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n913), .A2(KEYINPUT59), .A3(new_n640), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n845), .B(KEYINPUT121), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n915), .B1(new_n881), .B2(new_n747), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n884), .B1(new_n916), .B2(new_n293), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g718(.A(KEYINPUT122), .B(new_n884), .C1(new_n916), .C2(new_n293), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n846), .A2(KEYINPUT57), .A3(new_n515), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n639), .A3(new_n886), .ZN(new_n923));
  AND2_X1   g722(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n914), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n912), .A2(new_n925), .ZN(G1345gat));
  OAI21_X1  g725(.A(G155gat), .B1(new_n913), .B2(new_n747), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n608), .A2(new_n235), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n902), .B2(new_n928), .ZN(G1346gat));
  OAI21_X1  g728(.A(G162gat), .B1(new_n913), .B2(new_n572), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n571), .A2(new_n236), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n902), .B2(new_n931), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n663), .A2(new_n469), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n848), .A2(new_n851), .A3(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(new_n373), .A3(new_n661), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n663), .B1(new_n844), .B2(new_n845), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n475), .A2(new_n469), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(G169gat), .B1(new_n938), .B2(new_n660), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n935), .A2(new_n939), .ZN(G1348gat));
  OAI21_X1  g739(.A(G176gat), .B1(new_n934), .B2(new_n640), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n374), .A3(new_n639), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT123), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n941), .A2(new_n945), .A3(new_n942), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(G1349gat));
  OAI21_X1  g746(.A(G183gat), .B1(new_n934), .B2(new_n747), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n938), .A2(new_n400), .A3(new_n608), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT60), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT60), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n948), .A2(new_n952), .A3(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1350gat));
  NAND4_X1  g753(.A1(new_n936), .A2(new_n367), .A3(new_n571), .A4(new_n937), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT124), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n848), .A2(new_n571), .A3(new_n851), .A4(new_n933), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(G190gat), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n515), .B1(new_n844), .B2(new_n845), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT115), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n440), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n933), .ZN(new_n965));
  NOR4_X1   g764(.A1(new_n964), .A2(new_n850), .A3(new_n572), .A4(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(KEYINPUT125), .B1(new_n966), .B2(new_n367), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n958), .A2(new_n957), .A3(G190gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(new_n968), .A3(KEYINPUT61), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n961), .A2(new_n969), .ZN(G1351gat));
  NOR2_X1   g769(.A1(new_n758), .A2(new_n965), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n922), .A2(new_n660), .A3(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n922), .A2(KEYINPUT126), .A3(new_n660), .A4(new_n971), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n974), .A2(G197gat), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n899), .A2(new_n469), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n936), .A2(new_n977), .ZN(new_n978));
  OR3_X1    g777(.A1(new_n978), .A2(G197gat), .A3(new_n661), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n976), .A2(new_n979), .ZN(G1352gat));
  NAND2_X1  g779(.A1(new_n922), .A2(new_n971), .ZN(new_n981));
  OAI21_X1  g780(.A(G204gat), .B1(new_n981), .B2(new_n640), .ZN(new_n982));
  INV_X1    g781(.A(new_n978), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n984));
  AOI21_X1  g783(.A(G204gat), .B1(new_n984), .B2(KEYINPUT62), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n983), .A2(new_n639), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n984), .A2(KEYINPUT62), .ZN(new_n987));
  XNOR2_X1  g786(.A(new_n986), .B(new_n987), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n982), .A2(new_n988), .ZN(G1353gat));
  OR3_X1    g788(.A1(new_n978), .A2(G211gat), .A3(new_n747), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n922), .A2(new_n608), .A3(new_n971), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n991), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n992));
  AOI21_X1  g791(.A(KEYINPUT63), .B1(new_n991), .B2(G211gat), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(G1354gat));
  OAI21_X1  g793(.A(G218gat), .B1(new_n981), .B2(new_n572), .ZN(new_n995));
  OR3_X1    g794(.A1(new_n978), .A2(G218gat), .A3(new_n572), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1355gat));
endmodule


