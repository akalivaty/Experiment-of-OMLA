//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(KEYINPUT15), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT87), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n208), .B1(new_n206), .B2(KEYINPUT15), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(new_n202), .A3(new_n203), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT88), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(KEYINPUT88), .A3(new_n213), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT15), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n210), .A2(new_n217), .A3(KEYINPUT89), .A4(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT89), .ZN(new_n220));
  INV_X1    g019(.A(G50gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G43gat), .ZN(new_n222));
  INV_X1    g021(.A(G43gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G50gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n204), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n222), .A2(new_n224), .A3(KEYINPUT15), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT87), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n229), .A3(new_n218), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n212), .A2(KEYINPUT88), .A3(new_n213), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(new_n214), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n220), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n219), .A2(new_n233), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n213), .A2(KEYINPUT86), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n213), .A2(KEYINPUT86), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n212), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n228), .B1(new_n237), .B2(new_n205), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G15gat), .B(G22gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT16), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(G1gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(G1gat), .B2(new_n241), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G8gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n246), .A2(KEYINPUT91), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT90), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n238), .B1(new_n219), .B2(new_n233), .ZN(new_n249));
  INV_X1    g048(.A(new_n245), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n240), .A2(KEYINPUT90), .A3(new_n245), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n246), .A2(KEYINPUT91), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n247), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G229gat), .A2(G233gat), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n256), .B(KEYINPUT13), .Z(new_n257));
  INV_X1    g056(.A(KEYINPUT18), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT17), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n259), .B1(new_n234), .B2(new_n239), .ZN(new_n260));
  AOI211_X1 g059(.A(KEYINPUT17), .B(new_n238), .C1(new_n219), .C2(new_n233), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n250), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n253), .A2(new_n262), .A3(new_n256), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n255), .A2(new_n257), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n253), .A2(new_n262), .A3(KEYINPUT18), .A4(new_n256), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT92), .B1(new_n263), .B2(new_n258), .ZN(new_n267));
  XNOR2_X1  g066(.A(G113gat), .B(G141gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(G197gat), .ZN(new_n269));
  XOR2_X1   g068(.A(KEYINPUT11), .B(G169gat), .Z(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n271), .B(KEYINPUT12), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n266), .A2(new_n274), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n264), .B(new_n265), .C1(new_n267), .C2(new_n273), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT80), .ZN(new_n279));
  OR2_X1    g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(KEYINPUT24), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G169gat), .ZN(new_n283));
  INV_X1    g082(.A(G176gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT23), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n281), .A2(KEYINPUT24), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n287), .A2(new_n288), .B1(G169gat), .B2(G176gat), .ZN(new_n289));
  AND4_X1   g088(.A1(new_n282), .A2(new_n285), .A3(new_n286), .A4(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(G169gat), .B2(G176gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT64), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n290), .A2(KEYINPUT65), .A3(KEYINPUT25), .A4(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n292), .B(KEYINPUT64), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n282), .A2(new_n285), .A3(new_n286), .A4(new_n289), .ZN(new_n297));
  OAI22_X1  g096(.A1(new_n296), .A2(new_n297), .B1(new_n287), .B2(new_n288), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT66), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n305), .A2(KEYINPUT26), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n305), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n306), .A2(new_n307), .B1(G183gat), .B2(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n299), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n310), .A2(new_n311), .A3(G226gat), .A4(G233gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(G226gat), .A2(G233gat), .ZN(new_n313));
  XOR2_X1   g112(.A(new_n313), .B(KEYINPUT76), .Z(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n295), .A2(new_n298), .B1(new_n304), .B2(new_n308), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n315), .B1(new_n316), .B2(KEYINPUT29), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT77), .B1(new_n316), .B2(new_n313), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n312), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT22), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n321), .A2(new_n322), .B1(G211gat), .B2(G218gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(new_n321), .B2(new_n322), .ZN(new_n324));
  XNOR2_X1  g123(.A(G211gat), .B(G218gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(G197gat), .B(G204gat), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n325), .B1(new_n324), .B2(new_n326), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n320), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n324), .A2(new_n326), .ZN(new_n330));
  INV_X1    g129(.A(new_n325), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(KEYINPUT75), .A3(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n313), .B1(new_n316), .B2(KEYINPUT29), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n310), .A2(new_n314), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n332), .A2(new_n333), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G8gat), .B(G36gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G64gat), .B(G92gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  NAND3_X1  g142(.A1(new_n336), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT78), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT30), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT30), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n344), .A2(KEYINPUT78), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n336), .A2(new_n340), .ZN(new_n349));
  INV_X1    g148(.A(new_n343), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT1), .ZN(new_n353));
  XNOR2_X1  g152(.A(G127gat), .B(G134gat), .ZN(new_n354));
  INV_X1    g153(.A(G113gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT67), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT67), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G113gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n358), .A3(G120gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT68), .ZN(new_n360));
  INV_X1    g159(.A(G120gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G113gat), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n359), .B2(new_n362), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n353), .B(new_n354), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n355), .A2(G120gat), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT1), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n367), .A2(new_n354), .ZN(new_n368));
  INV_X1    g167(.A(G155gat), .ZN(new_n369));
  INV_X1    g168(.A(G162gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT79), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n371), .A2(new_n375), .A3(new_n372), .ZN(new_n376));
  INV_X1    g175(.A(G141gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G148gat), .ZN(new_n378));
  INV_X1    g177(.A(G148gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(G141gat), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n378), .A2(new_n380), .B1(KEYINPUT2), .B2(new_n372), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n374), .A2(new_n376), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G141gat), .B(G148gat), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n372), .A2(KEYINPUT2), .ZN(new_n384));
  OAI211_X1 g183(.A(KEYINPUT79), .B(new_n373), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n365), .A2(new_n368), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT4), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n365), .A2(new_n389), .A3(new_n368), .A4(new_n386), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT3), .B1(new_n382), .B2(new_n385), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n365), .A2(new_n368), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n388), .A2(new_n390), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(KEYINPUT5), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT0), .ZN(new_n400));
  XNOR2_X1  g199(.A(G57gat), .B(G85gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n390), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n394), .A2(new_n395), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n404), .A2(new_n397), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT5), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n395), .A2(new_n385), .A3(new_n382), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n387), .ZN(new_n409));
  INV_X1    g208(.A(new_n397), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n398), .B(new_n403), .C1(new_n406), .C2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT6), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n412), .A2(new_n413), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n409), .A2(new_n410), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n416), .A2(KEYINPUT5), .B1(new_n396), .B2(new_n397), .ZN(new_n417));
  INV_X1    g216(.A(new_n398), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n402), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n279), .B1(new_n352), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n351), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n347), .B1(new_n344), .B2(KEYINPUT78), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n416), .A2(KEYINPUT5), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n396), .A2(new_n397), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n427), .A2(KEYINPUT6), .A3(new_n403), .A4(new_n398), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n403), .B1(new_n427), .B2(new_n398), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n424), .A2(new_n431), .A3(KEYINPUT80), .A4(new_n348), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT83), .ZN(new_n433));
  INV_X1    g232(.A(new_n393), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(KEYINPUT81), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT81), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(new_n393), .B2(KEYINPUT29), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n335), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n435), .B1(new_n327), .B2(new_n328), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n386), .B1(new_n440), .B2(new_n391), .ZN(new_n441));
  NAND2_X1  g240(.A1(G228gat), .A2(G233gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT82), .B(G22gat), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n339), .B1(new_n434), .B2(new_n435), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n442), .B1(new_n446), .B2(new_n441), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G78gat), .B(G106gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT31), .B(G50gat), .ZN(new_n450));
  XOR2_X1   g249(.A(new_n449), .B(new_n450), .Z(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G22gat), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(new_n444), .B2(new_n447), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n433), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n444), .A2(new_n447), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(G22gat), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n458), .A2(KEYINPUT83), .A3(new_n448), .A4(new_n452), .ZN(new_n459));
  INV_X1    g258(.A(new_n445), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n448), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n456), .A2(new_n459), .B1(new_n462), .B2(new_n451), .ZN(new_n463));
  INV_X1    g262(.A(new_n395), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n310), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n316), .A2(new_n395), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT32), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT33), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  XOR2_X1   g270(.A(G15gat), .B(G43gat), .Z(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT69), .ZN(new_n473));
  XNOR2_X1  g272(.A(G71gat), .B(G99gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n469), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT70), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(KEYINPUT33), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n468), .A2(KEYINPUT32), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT71), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n468), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n479), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT70), .A4(new_n475), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n478), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n466), .B1(new_n465), .B2(new_n467), .ZN(new_n487));
  OR3_X1    g286(.A1(new_n487), .A2(KEYINPUT72), .A3(KEYINPUT34), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT34), .B1(new_n487), .B2(KEYINPUT72), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n488), .A2(new_n489), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n492), .A2(new_n478), .A3(new_n484), .A4(new_n485), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n463), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n421), .A2(new_n432), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT85), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n491), .A2(new_n493), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n346), .A2(new_n348), .A3(new_n351), .ZN(new_n499));
  INV_X1    g298(.A(new_n463), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT35), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT84), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n419), .A2(new_n413), .A3(new_n412), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(new_n428), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n414), .A2(KEYINPUT84), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n497), .B1(new_n501), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n431), .A2(KEYINPUT84), .ZN(new_n509));
  INV_X1    g308(.A(new_n506), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT35), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n511), .A2(KEYINPUT85), .A3(new_n494), .A4(new_n499), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n421), .A2(new_n432), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n463), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT36), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n517), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n519), .A2(new_n517), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n518), .B1(new_n498), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n344), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n350), .B1(new_n349), .B2(KEYINPUT37), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n337), .A2(new_n338), .ZN(new_n525));
  OAI22_X1  g324(.A1(new_n339), .A2(new_n525), .B1(new_n319), .B2(new_n335), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT38), .B1(new_n526), .B2(KEYINPUT37), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n522), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT37), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n336), .B2(new_n340), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT38), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n509), .A2(new_n528), .A3(new_n510), .A4(new_n531), .ZN(new_n532));
  OR3_X1    g331(.A1(new_n396), .A2(KEYINPUT39), .A3(new_n397), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n408), .A2(new_n397), .A3(new_n387), .ZN(new_n534));
  OAI211_X1 g333(.A(KEYINPUT39), .B(new_n534), .C1(new_n396), .C2(new_n397), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n402), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT40), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n352), .A2(new_n412), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n532), .A2(new_n540), .A3(new_n500), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n515), .A2(new_n521), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n278), .B1(new_n513), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(KEYINPUT41), .ZN(new_n545));
  XNOR2_X1  g344(.A(G134gat), .B(G162gat), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n545), .B(new_n546), .Z(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G99gat), .B(G106gat), .Z(new_n549));
  NAND2_X1  g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT100), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT101), .ZN(new_n553));
  NAND3_X1  g352(.A1(KEYINPUT100), .A2(G85gat), .A3(G92gat), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT7), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  INV_X1    g355(.A(G85gat), .ZN(new_n557));
  INV_X1    g356(.A(G92gat), .ZN(new_n558));
  AOI22_X1  g357(.A1(KEYINPUT8), .A2(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT101), .B1(new_n550), .B2(KEYINPUT7), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT7), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(new_n550), .B2(new_n551), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n561), .B1(new_n554), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n549), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n552), .A2(KEYINPUT7), .A3(new_n554), .ZN(new_n566));
  INV_X1    g365(.A(new_n561), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n549), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n568), .A2(new_n569), .A3(new_n555), .A4(new_n559), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n565), .A2(new_n570), .A3(KEYINPUT102), .ZN(new_n571));
  INV_X1    g370(.A(new_n560), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT102), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n572), .A2(new_n573), .A3(new_n569), .A4(new_n568), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n576), .B1(new_n260), .B2(new_n261), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT103), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n240), .A2(new_n575), .B1(KEYINPUT41), .B2(new_n544), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n578), .B1(new_n577), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n301), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n240), .A2(KEYINPUT17), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n249), .A2(new_n259), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n575), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n544), .A2(KEYINPUT41), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(new_n576), .B2(new_n249), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT103), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(G190gat), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n582), .A2(G218gat), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT99), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(G218gat), .B1(new_n582), .B2(new_n590), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n548), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n582), .A2(new_n590), .ZN(new_n596));
  INV_X1    g395(.A(G218gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n598), .A2(new_n592), .A3(new_n591), .A4(new_n547), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n602));
  INV_X1    g401(.A(G57gat), .ZN(new_n603));
  OAI21_X1  g402(.A(G64gat), .B1(new_n603), .B2(KEYINPUT94), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT94), .ZN(new_n605));
  INV_X1    g404(.A(G64gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n606), .A3(G57gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(G71gat), .ZN(new_n609));
  INV_X1    g408(.A(G78gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT9), .ZN(new_n611));
  NAND2_X1  g410(.A1(G71gat), .A2(G78gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT93), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT93), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(G71gat), .B2(G78gat), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n618), .A3(new_n612), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT9), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n606), .A2(G57gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n603), .A2(G64gat), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n602), .B1(new_n615), .B2(new_n624), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n614), .B(KEYINPUT95), .C1(new_n623), .C2(new_n619), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n625), .A2(KEYINPUT97), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT97), .B1(new_n625), .B2(new_n626), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT21), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n250), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n630), .A2(KEYINPUT98), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(KEYINPUT98), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G231gat), .A2(G233gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT96), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n633), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n625), .A2(new_n626), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(KEYINPUT21), .ZN(new_n641));
  XOR2_X1   g440(.A(G127gat), .B(G155gat), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G183gat), .B(G211gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n639), .A2(new_n645), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n571), .A2(new_n625), .A3(new_n626), .A4(new_n574), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n615), .A2(new_n624), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n565), .A3(new_n570), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  OAI211_X1 g452(.A(KEYINPUT10), .B(new_n575), .C1(new_n627), .C2(new_n628), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G230gat), .A2(G233gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n649), .A2(new_n652), .ZN(new_n658));
  INV_X1    g457(.A(new_n656), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(new_n663), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n664), .B1(new_n657), .B2(new_n660), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n601), .A2(new_n648), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n543), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n420), .A2(KEYINPUT104), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n431), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  NAND3_X1  g478(.A1(new_n671), .A2(new_n352), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(G8gat), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(new_n671), .B2(new_n352), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT105), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n680), .A2(new_n681), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(G1325gat));
  INV_X1    g488(.A(new_n671), .ZN(new_n690));
  OAI21_X1  g489(.A(G15gat), .B1(new_n690), .B2(new_n521), .ZN(new_n691));
  INV_X1    g490(.A(new_n498), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n692), .A2(G15gat), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n690), .B2(new_n693), .ZN(G1326gat));
  AND2_X1   g493(.A1(new_n543), .A2(new_n463), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n670), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT43), .B(G22gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  INV_X1    g497(.A(new_n668), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n648), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n277), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT108), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n601), .B1(new_n513), .B2(new_n542), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n513), .A2(new_n542), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n706), .A2(new_n707), .A3(new_n600), .ZN(new_n708));
  AOI22_X1  g507(.A1(KEYINPUT109), .A2(new_n705), .B1(new_n708), .B2(KEYINPUT44), .ZN(new_n709));
  AOI211_X1 g508(.A(KEYINPUT110), .B(new_n601), .C1(new_n513), .C2(new_n542), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n710), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n676), .B(new_n702), .C1(new_n709), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT111), .ZN(new_n714));
  INV_X1    g513(.A(new_n702), .ZN(new_n715));
  AOI211_X1 g514(.A(KEYINPUT109), .B(new_n601), .C1(new_n513), .C2(new_n542), .ZN(new_n716));
  OAI22_X1  g515(.A1(new_n707), .A2(new_n710), .B1(new_n716), .B2(new_n711), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n705), .A2(KEYINPUT109), .A3(KEYINPUT44), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(new_n720), .A3(new_n676), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n714), .A2(new_n721), .A3(G29gat), .ZN(new_n722));
  AOI211_X1 g521(.A(new_n601), .B(new_n701), .C1(new_n513), .C2(new_n542), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n202), .A3(new_n676), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n724), .A2(KEYINPUT107), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(KEYINPUT107), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(KEYINPUT45), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n722), .A2(new_n727), .A3(new_n730), .ZN(G1328gat));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(KEYINPUT112), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT112), .B(KEYINPUT46), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n723), .A2(new_n203), .A3(new_n352), .ZN(new_n735));
  MUX2_X1   g534(.A(new_n733), .B(new_n734), .S(new_n735), .Z(new_n736));
  OAI211_X1 g535(.A(new_n352), .B(new_n702), .C1(new_n709), .C2(new_n712), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT113), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G36gat), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n737), .A2(new_n738), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n736), .B1(new_n740), .B2(new_n741), .ZN(G1329gat));
  NOR2_X1   g541(.A1(new_n521), .A2(new_n223), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n702), .B(new_n743), .C1(new_n709), .C2(new_n712), .ZN(new_n744));
  INV_X1    g543(.A(new_n723), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n223), .B1(new_n745), .B2(new_n692), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n221), .B1(new_n719), .B2(new_n463), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n700), .A2(new_n221), .A3(new_n600), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n695), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n749), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n702), .B1(new_n709), .B2(new_n712), .ZN(new_n755));
  OAI21_X1  g554(.A(G50gat), .B1(new_n755), .B2(new_n500), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(KEYINPUT48), .A3(new_n752), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(G1331gat));
  INV_X1    g557(.A(new_n648), .ZN(new_n759));
  NOR4_X1   g558(.A1(new_n759), .A2(new_n600), .A3(new_n277), .A4(new_n668), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n706), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n675), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(new_n603), .ZN(G1332gat));
  NOR2_X1   g562(.A1(new_n761), .A2(new_n499), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  AND2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n764), .B2(new_n765), .ZN(G1333gat));
  OAI21_X1  g567(.A(G71gat), .B1(new_n761), .B2(new_n521), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n498), .A2(new_n609), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n761), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g571(.A1(new_n761), .A2(new_n500), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(new_n610), .ZN(G1335gat));
  NOR2_X1   g573(.A1(new_n648), .A2(new_n277), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n699), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n776), .B(KEYINPUT114), .Z(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n709), .B2(new_n712), .ZN(new_n778));
  OAI21_X1  g577(.A(G85gat), .B1(new_n778), .B2(new_n675), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n703), .A2(KEYINPUT51), .A3(new_n775), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT51), .B1(new_n703), .B2(new_n775), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n699), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(new_n557), .A3(new_n676), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n779), .A2(new_n785), .ZN(G1336gat));
  INV_X1    g585(.A(new_n777), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n717), .B2(new_n718), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n558), .B1(new_n788), .B2(new_n352), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n352), .A2(new_n558), .A3(new_n699), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT115), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n781), .B2(new_n782), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT52), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G92gat), .B1(new_n778), .B2(new_n499), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n796), .A3(new_n792), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n797), .ZN(G1337gat));
  OAI21_X1  g597(.A(G99gat), .B1(new_n778), .B2(new_n521), .ZN(new_n799));
  OR3_X1    g598(.A1(new_n783), .A2(G99gat), .A3(new_n692), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(G1338gat));
  INV_X1    g600(.A(G106gat), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n783), .B2(new_n500), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n500), .A2(new_n802), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n777), .B(new_n804), .C1(new_n709), .C2(new_n712), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n803), .A2(KEYINPUT53), .A3(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(G1339gat));
  NOR2_X1   g609(.A1(new_n255), .A2(new_n257), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n256), .B1(new_n253), .B2(new_n262), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n271), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n266), .B2(new_n272), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n699), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n653), .A2(new_n654), .A3(new_n659), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n659), .B1(new_n653), .B2(new_n654), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT116), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n657), .A2(new_n821), .A3(KEYINPUT54), .A4(new_n817), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n664), .B1(new_n819), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT55), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n655), .A2(new_n824), .A3(new_n656), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(KEYINPUT55), .A3(new_n665), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n823), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n666), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT117), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n829), .B1(new_n820), .B2(new_n822), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n834), .A2(new_n835), .A3(new_n666), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n827), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n816), .B1(new_n837), .B2(new_n278), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n601), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n834), .A2(new_n666), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT117), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n835), .B1(new_n834), .B2(new_n666), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n826), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n600), .A2(new_n815), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n648), .B1(new_n839), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n669), .A2(new_n277), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n463), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n676), .A2(new_n499), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n692), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851), .B2(new_n278), .ZN(new_n852));
  INV_X1    g651(.A(new_n501), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n853), .B(new_n676), .C1(new_n845), .C2(new_n846), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n277), .A2(new_n356), .A3(new_n358), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(G1340gat));
  NOR3_X1   g655(.A1(new_n851), .A2(new_n361), .A3(new_n668), .ZN(new_n857));
  INV_X1    g656(.A(new_n854), .ZN(new_n858));
  AOI21_X1  g657(.A(G120gat), .B1(new_n858), .B2(new_n699), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n857), .A2(new_n859), .ZN(G1341gat));
  OR3_X1    g659(.A1(new_n854), .A2(KEYINPUT118), .A3(new_n759), .ZN(new_n861));
  INV_X1    g660(.A(G127gat), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT118), .B1(new_n854), .B2(new_n759), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n848), .A2(G127gat), .A3(new_n648), .A4(new_n850), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n864), .A2(KEYINPUT119), .A3(new_n865), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1342gat));
  OR3_X1    g669(.A1(new_n854), .A2(G134gat), .A3(new_n601), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n851), .B2(new_n601), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G1343gat));
  INV_X1    g674(.A(new_n521), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n849), .ZN(new_n877));
  XOR2_X1   g676(.A(new_n877), .B(KEYINPUT120), .Z(new_n878));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(new_n847), .B2(new_n500), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n500), .A2(new_n879), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n277), .A2(new_n827), .A3(new_n840), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n816), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n601), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n648), .B1(new_n884), .B2(new_n844), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n881), .B1(new_n885), .B2(new_n846), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n878), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n377), .B1(new_n887), .B2(new_n277), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n847), .A2(new_n675), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n876), .A2(new_n352), .A3(new_n500), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(G141gat), .A3(new_n278), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT58), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n891), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n377), .A3(new_n277), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  AOI211_X1 g695(.A(new_n278), .B(new_n878), .C1(new_n880), .C2(new_n886), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n895), .B(new_n896), .C1(new_n897), .C2(new_n377), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n893), .A2(new_n898), .ZN(G1344gat));
  NAND2_X1  g698(.A1(new_n699), .A2(new_n379), .ZN(new_n900));
  OR3_X1    g699(.A1(new_n891), .A2(KEYINPUT121), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT121), .B1(new_n891), .B2(new_n900), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n600), .A2(KEYINPUT122), .A3(new_n843), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n815), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT122), .B1(new_n600), .B2(new_n843), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n884), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n759), .ZN(new_n908));
  INV_X1    g707(.A(new_n846), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT57), .B1(new_n910), .B2(new_n463), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n847), .A2(new_n879), .A3(new_n500), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n878), .A2(new_n668), .ZN(new_n914));
  OAI211_X1 g713(.A(KEYINPUT59), .B(G148gat), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n379), .B1(new_n887), .B2(new_n699), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n903), .B(new_n915), .C1(KEYINPUT59), .C2(new_n916), .ZN(G1345gat));
  NAND3_X1  g716(.A1(new_n894), .A2(new_n369), .A3(new_n648), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n887), .A2(new_n648), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n369), .ZN(G1346gat));
  AOI21_X1  g719(.A(G162gat), .B1(new_n894), .B2(new_n600), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n601), .A2(new_n370), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n887), .B2(new_n922), .ZN(G1347gat));
  OR2_X1    g722(.A1(new_n845), .A2(new_n846), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n676), .A2(new_n499), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n498), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT123), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n924), .A2(new_n500), .A3(new_n927), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n928), .A2(new_n283), .A3(new_n278), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n494), .A2(new_n352), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n924), .A2(new_n675), .A3(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n277), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n929), .B1(new_n283), .B2(new_n933), .ZN(G1348gat));
  OAI21_X1  g733(.A(new_n284), .B1(new_n931), .B2(new_n668), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT124), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n928), .A2(new_n284), .A3(new_n668), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(G1349gat));
  OAI21_X1  g737(.A(G183gat), .B1(new_n928), .B2(new_n759), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT60), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n847), .A2(new_n676), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n942), .A2(new_n300), .A3(new_n648), .A4(new_n930), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n939), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n940), .A2(KEYINPUT60), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n944), .B(new_n945), .ZN(G1350gat));
  NAND3_X1  g745(.A1(new_n932), .A2(new_n301), .A3(new_n600), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n848), .A2(new_n600), .A3(new_n927), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(new_n949), .A3(G190gat), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n949), .B1(new_n948), .B2(G190gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(G1351gat));
  NAND2_X1  g752(.A1(new_n925), .A2(new_n521), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n846), .B1(new_n907), .B2(new_n759), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n879), .B1(new_n955), .B2(new_n500), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n924), .A2(new_n881), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n958), .A2(new_n277), .ZN(new_n959));
  XOR2_X1   g758(.A(KEYINPUT126), .B(G197gat), .Z(new_n960));
  NOR3_X1   g759(.A1(new_n876), .A2(new_n499), .A3(new_n500), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n961), .B(new_n675), .C1(new_n845), .C2(new_n846), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n277), .A2(new_n960), .ZN(new_n963));
  OAI22_X1  g762(.A1(new_n959), .A2(new_n960), .B1(new_n962), .B2(new_n963), .ZN(G1352gat));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n965));
  INV_X1    g764(.A(G204gat), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n966), .B1(new_n958), .B2(new_n699), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n668), .A2(G204gat), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  OR3_X1    g768(.A1(new_n962), .A2(KEYINPUT62), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT62), .B1(new_n962), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n965), .B1(new_n967), .B2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(new_n972), .ZN(new_n974));
  AOI211_X1 g773(.A(new_n668), .B(new_n954), .C1(new_n956), .C2(new_n957), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n974), .B(KEYINPUT127), .C1(new_n975), .C2(new_n966), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n973), .A2(new_n976), .ZN(G1353gat));
  INV_X1    g776(.A(G211gat), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n942), .A2(new_n978), .A3(new_n648), .A4(new_n961), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT63), .ZN(new_n980));
  AOI211_X1 g779(.A(new_n980), .B(new_n978), .C1(new_n958), .C2(new_n648), .ZN(new_n981));
  INV_X1    g780(.A(new_n954), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n648), .B(new_n982), .C1(new_n911), .C2(new_n912), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT63), .B1(new_n983), .B2(G211gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n979), .B1(new_n981), .B2(new_n984), .ZN(G1354gat));
  AND2_X1   g784(.A1(new_n958), .A2(new_n600), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n600), .A2(new_n597), .ZN(new_n987));
  OAI22_X1  g786(.A1(new_n986), .A2(new_n597), .B1(new_n962), .B2(new_n987), .ZN(G1355gat));
endmodule


