//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  AND2_X1   g003(.A1(new_n204), .A2(KEYINPUT83), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(KEYINPUT83), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  AND2_X1   g007(.A1(G211gat), .A2(G218gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(KEYINPUT22), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT72), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n215));
  AND2_X1   g014(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n216));
  AND2_X1   g015(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n218));
  OAI22_X1  g017(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT2), .ZN(new_n220));
  XOR2_X1   g019(.A(G155gat), .B(G162gat), .Z(new_n221));
  OR2_X1    g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT2), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n222), .A2(new_n226), .A3(new_n223), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n220), .A2(new_n225), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT3), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n214), .B1(KEYINPUT29), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n229), .B1(new_n212), .B2(KEYINPUT29), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n221), .A2(new_n227), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT75), .B(G155gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT76), .B(G162gat), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n226), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G155gat), .B(G162gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(new_n222), .A3(new_n223), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n234), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n233), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n232), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G22gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G228gat), .A2(G233gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n232), .A2(G22gat), .A3(new_n241), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n245), .B1(new_n244), .B2(new_n246), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n207), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n246), .ZN(new_n250));
  AOI21_X1  g049(.A(G22gat), .B1(new_n232), .B2(new_n241), .ZN(new_n251));
  OAI211_X1 g050(.A(G228gat), .B(G233gat), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n253), .A3(new_n205), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G1gat), .B(G29gat), .Z(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G57gat), .B(G85gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G127gat), .B(G134gat), .Z(new_n262));
  XNOR2_X1  g061(.A(G113gat), .B(G120gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n262), .B1(KEYINPUT1), .B2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G113gat), .B(G120gat), .Z(new_n265));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n266));
  XNOR2_X1  g065(.A(G127gat), .B(G134gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n240), .B(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G225gat), .A2(G233gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n271), .B(KEYINPUT77), .Z(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT5), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n264), .A2(new_n268), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n275), .B1(new_n228), .B2(new_n229), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n240), .A2(KEYINPUT3), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n272), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n228), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n281), .B1(new_n228), .B2(new_n275), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT79), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n281), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n283), .B(new_n285), .C1(new_n240), .C2(new_n269), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n278), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT80), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n240), .A2(new_n269), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT79), .B1(new_n290), .B2(new_n281), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(new_n286), .A3(new_n280), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT80), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(new_n293), .A3(new_n278), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n274), .B1(new_n289), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n278), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n290), .A2(new_n285), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(KEYINPUT4), .B2(new_n290), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n296), .A2(new_n298), .A3(KEYINPUT5), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n261), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n301));
  INV_X1    g100(.A(new_n274), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n292), .A2(new_n293), .A3(new_n278), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n293), .B1(new_n292), .B2(new_n278), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n299), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n260), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n300), .A2(new_n301), .A3(new_n307), .ZN(new_n308));
  OAI211_X1 g107(.A(KEYINPUT6), .B(new_n261), .C1(new_n295), .C2(new_n299), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G226gat), .A2(G233gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT24), .ZN(new_n313));
  INV_X1    g112(.A(G183gat), .ZN(new_n314));
  INV_X1    g113(.A(G190gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n316), .B(new_n317), .C1(G183gat), .C2(G190gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT23), .ZN(new_n320));
  NAND2_X1  g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n319), .A2(KEYINPUT23), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n318), .A2(new_n320), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT25), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AND4_X1   g124(.A1(KEYINPUT25), .A2(new_n322), .A3(new_n320), .A4(new_n321), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n317), .B(KEYINPUT65), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n314), .ZN(new_n329));
  NAND2_X1  g128(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n315), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n327), .A2(new_n316), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n325), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT67), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT27), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT27), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT67), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n338), .A3(G183gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n329), .A2(KEYINPUT27), .A3(new_n330), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n340), .A3(new_n315), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT68), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT28), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n342), .B1(new_n341), .B2(new_n343), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT27), .B(G183gat), .Z(new_n346));
  NOR3_X1   g145(.A1(new_n346), .A2(new_n343), .A3(G190gat), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n321), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n349), .A2(new_n319), .A3(KEYINPUT26), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n314), .A2(new_n315), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n319), .A2(KEYINPUT26), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n334), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n312), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n324), .A2(new_n323), .B1(new_n326), .B2(new_n332), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT68), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n361));
  INV_X1    g160(.A(new_n347), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n358), .B1(new_n363), .B2(new_n353), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(new_n311), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n214), .B1(new_n357), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  OAI21_X1  g168(.A(new_n311), .B1(new_n364), .B2(KEYINPUT29), .ZN(new_n370));
  INV_X1    g169(.A(new_n214), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n312), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n366), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT30), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT74), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(KEYINPUT74), .A3(new_n375), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n369), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n371), .B1(new_n370), .B2(new_n372), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n366), .A2(KEYINPUT30), .A3(new_n369), .A4(new_n373), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT73), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n382), .A2(new_n383), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT73), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT30), .A4(new_n369), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n310), .A2(new_n380), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT82), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n378), .A2(new_n379), .B1(new_n386), .B2(new_n389), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(new_n310), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n276), .A2(new_n277), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n397), .B(new_n297), .C1(KEYINPUT4), .C2(new_n290), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n272), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n399), .B(KEYINPUT39), .C1(new_n272), .C2(new_n270), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT39), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n398), .A2(new_n401), .A3(new_n272), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n260), .A3(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT40), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n404), .A2(new_n300), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n380), .A2(new_n406), .A3(new_n390), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(new_n380), .B2(new_n390), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT37), .B1(new_n382), .B2(new_n383), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT37), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n366), .A2(new_n411), .A3(new_n373), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n381), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT38), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n414), .B1(new_n413), .B2(KEYINPUT38), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT38), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n410), .A2(new_n412), .A3(new_n418), .A4(new_n381), .ZN(new_n419));
  AND4_X1   g218(.A1(new_n309), .A2(new_n308), .A3(new_n374), .A4(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n255), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n255), .A2(new_n396), .B1(new_n409), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n347), .B1(new_n359), .B2(KEYINPUT68), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n354), .B1(new_n423), .B2(new_n361), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n269), .B1(new_n424), .B2(new_n358), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n275), .B(new_n334), .C1(new_n348), .C2(new_n354), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G227gat), .A2(G233gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT34), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT70), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(KEYINPUT70), .B(KEYINPUT34), .C1(new_n427), .C2(new_n429), .ZN(new_n433));
  INV_X1    g232(.A(new_n427), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n428), .B(KEYINPUT64), .Z(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(KEYINPUT34), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n432), .A2(new_n433), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT69), .B1(new_n427), .B2(new_n435), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT69), .ZN(new_n439));
  INV_X1    g238(.A(new_n435), .ZN(new_n440));
  AOI211_X1 g239(.A(new_n439), .B(new_n440), .C1(new_n425), .C2(new_n426), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT32), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n438), .B2(new_n441), .ZN(new_n444));
  XOR2_X1   g243(.A(G15gat), .B(G43gat), .Z(new_n445));
  XNOR2_X1  g244(.A(G71gat), .B(G99gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n442), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n447), .ZN(new_n449));
  OAI221_X1 g248(.A(KEYINPUT32), .B1(new_n443), .B2(new_n449), .C1(new_n438), .C2(new_n441), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n437), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT71), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT36), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n453), .A2(KEYINPUT36), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n448), .A2(new_n437), .A3(new_n450), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n452), .A2(new_n454), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n448), .A2(new_n437), .A3(new_n450), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n453), .B(KEYINPUT36), .C1(new_n458), .C2(new_n451), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n458), .A2(new_n451), .A3(new_n255), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n392), .A2(new_n395), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n407), .A2(new_n408), .ZN(new_n464));
  INV_X1    g263(.A(new_n310), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(KEYINPUT35), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n422), .A2(new_n460), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(G29gat), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n470));
  XOR2_X1   g269(.A(KEYINPUT14), .B(G29gat), .Z(new_n471));
  OAI21_X1  g270(.A(new_n470), .B1(new_n471), .B2(G36gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(G43gat), .B(G50gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT15), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n473), .A2(KEYINPUT15), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n472), .A2(new_n474), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n472), .A2(new_n475), .A3(KEYINPUT87), .A4(new_n474), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT16), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n482), .B1(new_n483), .B2(G1gat), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(G1gat), .B2(new_n482), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n485), .B(G8gat), .Z(new_n486));
  OAI21_X1  g285(.A(KEYINPUT90), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT90), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n485), .B(G8gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n487), .A2(new_n491), .B1(new_n481), .B2(new_n486), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494));
  XOR2_X1   g293(.A(new_n494), .B(KEYINPUT13), .Z(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(KEYINPUT91), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT91), .ZN(new_n497));
  INV_X1    g296(.A(new_n495), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(new_n492), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT18), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT88), .B(KEYINPUT17), .Z(new_n502));
  NAND2_X1  g301(.A1(new_n488), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT89), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT89), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n505), .A3(new_n502), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n488), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(new_n490), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n507), .A2(new_n510), .B1(new_n487), .B2(new_n491), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n501), .B1(new_n511), .B2(new_n494), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n507), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n487), .A2(new_n491), .ZN(new_n514));
  AND4_X1   g313(.A1(new_n501), .A2(new_n513), .A3(new_n514), .A4(new_n494), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n500), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G113gat), .B(G141gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G169gat), .B(G197gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n521), .B(KEYINPUT12), .Z(new_n522));
  NAND2_X1  g321(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT92), .ZN(new_n524));
  INV_X1    g323(.A(new_n522), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n500), .B(new_n525), .C1(new_n512), .C2(new_n515), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n516), .A2(KEYINPUT92), .A3(new_n522), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n468), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G183gat), .B(G211gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(G71gat), .A2(G78gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(G71gat), .A2(G78gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n537), .B(KEYINPUT96), .Z(new_n538));
  INV_X1    g337(.A(new_n536), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(KEYINPUT9), .ZN(new_n540));
  XNOR2_X1  g339(.A(G57gat), .B(G64gat), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(G57gat), .B(G64gat), .Z(new_n543));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(KEYINPUT94), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n540), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT95), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT93), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n536), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n535), .ZN(new_n551));
  OR3_X1    g350(.A1(new_n547), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n548), .B1(new_n547), .B2(new_n551), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n542), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(KEYINPUT21), .ZN(new_n555));
  NAND2_X1  g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G127gat), .B(G155gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT20), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n557), .B(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n490), .B1(new_n554), .B2(KEYINPUT21), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(KEYINPUT98), .Z(new_n562));
  AND2_X1   g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n560), .A2(new_n562), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n534), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n560), .A2(new_n562), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n560), .A2(new_n562), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n533), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G85gat), .A2(G92gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT7), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(G99gat), .A2(G106gat), .ZN(new_n573));
  INV_X1    g372(.A(G85gat), .ZN(new_n574));
  INV_X1    g373(.A(G92gat), .ZN(new_n575));
  AOI22_X1  g374(.A1(KEYINPUT8), .A2(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(KEYINPUT100), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n571), .A2(new_n576), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(new_n572), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n578), .B1(new_n580), .B2(KEYINPUT100), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n581), .B1(new_n508), .B2(new_n488), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n582), .B1(new_n504), .B2(new_n506), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G190gat), .B(G218gat), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT41), .ZN(new_n587));
  NAND2_X1  g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588));
  OAI22_X1  g387(.A1(new_n481), .A2(new_n581), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n584), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n587), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT99), .ZN(new_n593));
  XOR2_X1   g392(.A(G134gat), .B(G162gat), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n585), .B1(new_n583), .B2(new_n589), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n595), .B1(new_n591), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n569), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n552), .A2(new_n553), .ZN(new_n602));
  INV_X1    g401(.A(new_n542), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n605), .A3(new_n581), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n580), .A2(KEYINPUT100), .ZN(new_n607));
  INV_X1    g406(.A(new_n578), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(KEYINPUT101), .B1(new_n554), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n554), .A2(new_n580), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT103), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n606), .A2(new_n610), .A3(new_n617), .A4(new_n611), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n554), .A2(new_n609), .A3(KEYINPUT10), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n616), .B1(new_n620), .B2(new_n613), .ZN(new_n621));
  AOI211_X1 g420(.A(KEYINPUT103), .B(new_n614), .C1(new_n618), .C2(new_n619), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n615), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(KEYINPUT102), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n620), .A2(new_n613), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n629), .A2(new_n626), .A3(new_n615), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n601), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n530), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n465), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G1gat), .ZN(G1324gat));
  INV_X1    g435(.A(new_n464), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n530), .A2(new_n637), .A3(new_n633), .ZN(new_n638));
  AND2_X1   g437(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(KEYINPUT42), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT104), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n641), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n638), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(G1325gat));
  INV_X1    g444(.A(G15gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n458), .A2(new_n451), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n634), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n460), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n634), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n650), .B2(new_n646), .ZN(G1326gat));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n255), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT43), .B(G22gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1327gat));
  INV_X1    g453(.A(new_n569), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n630), .B1(new_n623), .B2(new_n627), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR4_X1   g456(.A1(new_n468), .A2(new_n529), .A3(new_n600), .A4(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n658), .A2(new_n469), .A3(new_n465), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n659), .A2(KEYINPUT105), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(KEYINPUT105), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(KEYINPUT45), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n463), .A2(new_n467), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n409), .A2(new_n421), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n393), .A2(new_n394), .A3(new_n310), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n394), .B1(new_n393), .B2(new_n310), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n255), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n664), .A2(new_n667), .A3(new_n460), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT44), .B1(new_n669), .B2(new_n599), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  AOI211_X1 g470(.A(new_n671), .B(new_n600), .C1(new_n663), .C2(new_n668), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n529), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G29gat), .B1(new_n675), .B2(new_n310), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n662), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT45), .B1(new_n660), .B2(new_n661), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n677), .A2(new_n678), .ZN(G1328gat));
  INV_X1    g478(.A(G36gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n658), .A2(new_n680), .A3(new_n637), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT46), .Z(new_n682));
  OAI21_X1  g481(.A(G36gat), .B1(new_n675), .B2(new_n464), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(G1329gat));
  NAND3_X1  g483(.A1(new_n673), .A2(new_n649), .A3(new_n674), .ZN(new_n685));
  INV_X1    g484(.A(new_n647), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(G43gat), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n685), .A2(G43gat), .B1(new_n658), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n688), .B(new_n689), .Z(G1330gat));
  INV_X1    g489(.A(new_n255), .ZN(new_n691));
  OAI21_X1  g490(.A(G50gat), .B1(new_n675), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT48), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(G50gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n658), .A2(new_n695), .A3(new_n255), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n694), .B(new_n697), .ZN(G1331gat));
  AND2_X1   g497(.A1(new_n527), .A2(new_n528), .ZN(new_n699));
  NOR4_X1   g498(.A1(new_n468), .A2(new_n699), .A3(new_n601), .A4(new_n656), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n465), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT108), .B(G57gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1332gat));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n637), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT49), .B(G64gat), .Z(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n704), .B2(new_n706), .ZN(G1333gat));
  INV_X1    g506(.A(G71gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n700), .A2(new_n708), .A3(new_n647), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n700), .A2(new_n649), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n710), .B2(new_n708), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g511(.A1(new_n700), .A2(new_n255), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT109), .B(G78gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1335gat));
  NOR3_X1   g514(.A1(new_n656), .A2(G85gat), .A3(new_n310), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n699), .A2(new_n569), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n664), .A2(new_n460), .A3(new_n667), .ZN(new_n718));
  INV_X1    g517(.A(new_n408), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n393), .A2(new_n406), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n461), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n721), .A2(new_n466), .B1(new_n462), .B2(KEYINPUT35), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n599), .B(new_n717), .C1(new_n718), .C2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT51), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n669), .A2(KEYINPUT51), .A3(new_n599), .A4(new_n717), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n723), .A2(KEYINPUT111), .A3(new_n724), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n716), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n717), .B2(new_n632), .ZN(new_n735));
  NOR4_X1   g534(.A1(new_n699), .A2(new_n569), .A3(KEYINPUT110), .A4(new_n656), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n673), .A2(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n738), .A2(new_n465), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n733), .B1(new_n574), .B2(new_n739), .ZN(G1336gat));
  OAI21_X1  g539(.A(new_n671), .B1(new_n468), .B2(new_n600), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n669), .A2(KEYINPUT44), .A3(new_n599), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n741), .A2(new_n637), .A3(new_n742), .A4(new_n737), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G92gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT113), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n725), .A2(new_n727), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n464), .A2(G92gat), .A3(new_n656), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n744), .A2(KEYINPUT113), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT52), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT115), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n673), .A2(new_n753), .A3(new_n637), .A4(new_n737), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n743), .A2(KEYINPUT114), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n755), .A3(G92gat), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n728), .A2(new_n730), .A3(new_n747), .ZN(new_n758));
  AND4_X1   g557(.A1(new_n752), .A2(new_n756), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n758), .A2(new_n757), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n752), .B1(new_n760), .B2(new_n756), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n751), .B1(new_n759), .B2(new_n761), .ZN(G1337gat));
  NOR3_X1   g561(.A1(new_n686), .A2(G99gat), .A3(new_n656), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT116), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n731), .B2(new_n732), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n738), .A2(new_n649), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G99gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1338gat));
  NAND2_X1  g567(.A1(new_n738), .A2(new_n255), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G106gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n656), .A2(G106gat), .A3(new_n691), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n728), .A2(new_n730), .A3(new_n773), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n769), .A2(G106gat), .B1(new_n746), .B2(new_n773), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n772), .A2(new_n774), .B1(new_n775), .B2(new_n771), .ZN(G1339gat));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n620), .B2(new_n613), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n618), .A2(KEYINPUT117), .A3(new_n614), .A4(new_n619), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n620), .B2(new_n613), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n629), .A2(KEYINPUT103), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n620), .A2(new_n616), .A3(new_n613), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(new_n781), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n626), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n783), .A2(new_n786), .A3(KEYINPUT55), .A4(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n788), .A2(new_n631), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n783), .A2(new_n787), .A3(new_n786), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(new_n699), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n511), .A2(new_n494), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n493), .A2(new_n495), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n521), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n526), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n794), .B1(new_n632), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n656), .A2(KEYINPUT119), .A3(new_n798), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n599), .B1(new_n793), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n599), .A2(new_n526), .A3(new_n797), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n792), .A2(new_n631), .A3(new_n788), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT118), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n804), .B1(new_n790), .B2(new_n791), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n789), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n655), .B1(new_n803), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n633), .A2(new_n529), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n637), .A2(new_n310), .A3(new_n686), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n691), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(G113gat), .B1(new_n816), .B2(new_n529), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n310), .B1(new_n812), .B2(new_n813), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n721), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n529), .A2(G113gat), .ZN(new_n820));
  XOR2_X1   g619(.A(new_n820), .B(KEYINPUT120), .Z(new_n821));
  OAI21_X1  g620(.A(new_n817), .B1(new_n819), .B2(new_n821), .ZN(G1340gat));
  INV_X1    g621(.A(G120gat), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n816), .A2(new_n823), .A3(new_n656), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n818), .A2(new_n721), .A3(new_n632), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n823), .B2(new_n825), .ZN(G1341gat));
  INV_X1    g625(.A(G127gat), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n816), .A2(new_n827), .A3(new_n655), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n819), .A2(KEYINPUT121), .A3(new_n655), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(G127gat), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT121), .B1(new_n819), .B2(new_n655), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(G1342gat));
  OR2_X1    g631(.A1(new_n600), .A2(G134gat), .ZN(new_n833));
  OR3_X1    g632(.A1(new_n819), .A2(KEYINPUT56), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G134gat), .B1(new_n816), .B2(new_n600), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT56), .B1(new_n819), .B2(new_n833), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(G1343gat));
  INV_X1    g636(.A(G141gat), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n460), .A2(new_n255), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n839), .A2(new_n637), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n818), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n838), .B1(new_n841), .B2(new_n529), .ZN(new_n842));
  INV_X1    g641(.A(new_n813), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n789), .A2(new_n808), .A3(new_n809), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n808), .B1(new_n789), .B2(new_n809), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n788), .A2(new_n631), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n621), .A2(new_n622), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n626), .B1(new_n848), .B2(new_n781), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT55), .B1(new_n849), .B2(new_n783), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n847), .A2(new_n529), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n656), .A2(new_n798), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n600), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n843), .B1(new_n854), .B2(new_n655), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT57), .B1(new_n855), .B2(new_n691), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n691), .B1(new_n812), .B2(new_n813), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n649), .A2(new_n310), .A3(new_n637), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n529), .A2(new_n838), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n842), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n864), .B(new_n865), .ZN(G1344gat));
  NOR2_X1   g665(.A1(new_n841), .A2(new_n656), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n867), .A2(new_n868), .A3(G148gat), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n861), .B2(new_n656), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n691), .A2(KEYINPUT57), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n852), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n599), .B1(new_n793), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n806), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n655), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n872), .B1(new_n876), .B2(new_n813), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n632), .A2(new_n794), .A3(new_n799), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT119), .B1(new_n656), .B2(new_n798), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n600), .B1(new_n851), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n569), .B1(new_n846), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n255), .B1(new_n882), .B2(new_n843), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n877), .B1(new_n883), .B2(KEYINPUT57), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n860), .A2(KEYINPUT122), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n860), .A2(KEYINPUT122), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n656), .A2(new_n868), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n884), .A2(new_n885), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n870), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n869), .B1(new_n889), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g689(.A(new_n235), .B1(new_n861), .B2(new_n655), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n655), .A2(new_n235), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n841), .B2(new_n892), .ZN(G1346gat));
  INV_X1    g692(.A(new_n236), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n861), .A2(new_n894), .A3(new_n600), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n818), .A2(new_n599), .A3(new_n840), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n894), .B2(new_n896), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n464), .A2(new_n465), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n814), .A2(new_n647), .A3(new_n691), .A4(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(G169gat), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n899), .A2(new_n900), .A3(new_n529), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n814), .A2(new_n310), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT123), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n814), .A2(new_n904), .A3(new_n310), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n464), .A2(new_n686), .A3(new_n255), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n699), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n901), .B1(new_n908), .B2(new_n900), .ZN(G1348gat));
  NOR2_X1   g708(.A1(new_n656), .A2(G176gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n906), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G176gat), .B1(new_n899), .B2(new_n656), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n911), .A2(KEYINPUT124), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1349gat));
  NOR2_X1   g716(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n918));
  AND2_X1   g717(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n655), .A2(new_n346), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n904), .B1(new_n814), .B2(new_n310), .ZN(new_n921));
  AOI211_X1 g720(.A(KEYINPUT123), .B(new_n465), .C1(new_n812), .C2(new_n813), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n907), .B(new_n920), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n329), .A2(new_n330), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n924), .B1(new_n899), .B2(new_n655), .ZN(new_n925));
  AOI211_X1 g724(.A(new_n918), .B(new_n919), .C1(new_n923), .C2(new_n925), .ZN(new_n926));
  AND4_X1   g725(.A1(KEYINPUT125), .A2(new_n923), .A3(KEYINPUT60), .A4(new_n925), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(G1350gat));
  NAND4_X1  g727(.A1(new_n906), .A2(new_n315), .A3(new_n599), .A4(new_n907), .ZN(new_n929));
  OAI21_X1  g728(.A(G190gat), .B1(new_n899), .B2(new_n600), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(KEYINPUT61), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(KEYINPUT61), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1351gat));
  AOI21_X1  g732(.A(new_n569), .B1(new_n853), .B2(new_n806), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n871), .B1(new_n934), .B2(new_n843), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n898), .A2(new_n460), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n935), .B(new_n936), .C1(new_n857), .C2(new_n858), .ZN(new_n937));
  INV_X1    g736(.A(G197gat), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n937), .A2(new_n938), .A3(new_n529), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n839), .A2(new_n464), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n906), .A2(new_n699), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n941), .B2(new_n938), .ZN(G1352gat));
  NOR2_X1   g741(.A1(new_n656), .A2(G204gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n906), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT62), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n906), .A2(new_n946), .A3(new_n940), .A4(new_n943), .ZN(new_n947));
  OAI21_X1  g746(.A(G204gat), .B1(new_n937), .B2(new_n656), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(G1353gat));
  OAI21_X1  g748(.A(KEYINPUT127), .B1(new_n937), .B2(new_n655), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n884), .A2(new_n951), .A3(new_n569), .A4(new_n936), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n950), .A2(new_n952), .A3(G211gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT63), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT63), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n950), .A2(new_n952), .A3(new_n955), .A4(G211gat), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n655), .A2(G211gat), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n906), .A2(new_n957), .A3(new_n940), .A4(new_n958), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n940), .B(new_n958), .C1(new_n921), .C2(new_n922), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(KEYINPUT126), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n954), .A2(new_n956), .A3(new_n962), .ZN(G1354gat));
  OAI21_X1  g762(.A(G218gat), .B1(new_n937), .B2(new_n600), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n906), .A2(new_n940), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n600), .A2(G218gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(G1355gat));
endmodule


