//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n588, new_n589, new_n590, new_n591, new_n593, new_n594, new_n596,
    new_n597, new_n598, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901;
  XOR2_X1   g000(.A(G155gat), .B(G162gat), .Z(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT2), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT75), .ZN(new_n206));
  XOR2_X1   g005(.A(G141gat), .B(G148gat), .Z(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n205), .A2(KEYINPUT75), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n202), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n205), .A2(KEYINPUT76), .ZN(new_n211));
  INV_X1    g010(.A(new_n202), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n205), .A2(KEYINPUT76), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n207), .A4(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT29), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(KEYINPUT80), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT72), .B(G197gat), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n222), .A2(G204gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(G204gat), .ZN(new_n224));
  INV_X1    g023(.A(G211gat), .ZN(new_n225));
  INV_X1    g024(.A(G218gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI22_X1  g026(.A1(new_n223), .A2(new_n224), .B1(KEYINPUT22), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(KEYINPUT73), .ZN(new_n229));
  XOR2_X1   g028(.A(G211gat), .B(G218gat), .Z(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n231), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n220), .A2(KEYINPUT80), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n221), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n232), .A2(new_n233), .A3(new_n219), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n216), .B1(new_n237), .B2(new_n217), .ZN(new_n238));
  OAI211_X1 g037(.A(G228gat), .B(G233gat), .C1(new_n236), .C2(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n238), .A2(KEYINPUT79), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n234), .A2(new_n220), .B1(G228gat), .B2(G233gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n238), .B2(KEYINPUT79), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n239), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G22gat), .ZN(new_n244));
  INV_X1    g043(.A(G22gat), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n239), .B(new_n245), .C1(new_n240), .C2(new_n242), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G78gat), .B(G106gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT31), .B(G50gat), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n248), .B(new_n249), .Z(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT81), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT81), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n244), .A2(new_n253), .A3(new_n246), .A4(new_n250), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n250), .B1(new_n244), .B2(new_n246), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(KEYINPUT82), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n256), .A2(KEYINPUT82), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT83), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n256), .B(KEYINPUT82), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT83), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n261), .A2(new_n262), .A3(new_n255), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G1gat), .B(G29gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT0), .ZN(new_n266));
  XNOR2_X1  g065(.A(G57gat), .B(G85gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  XOR2_X1   g067(.A(G113gat), .B(G120gat), .Z(new_n269));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G127gat), .B(G134gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT1), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n273), .B(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n276), .A2(new_n215), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(KEYINPUT4), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(KEYINPUT77), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(KEYINPUT4), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n215), .A2(KEYINPUT3), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n218), .A2(new_n276), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G225gat), .A2(G233gat), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n280), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT78), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n276), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(new_n216), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n279), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n284), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n277), .A2(KEYINPUT4), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n294), .B(new_n285), .C1(new_n279), .C2(KEYINPUT4), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(KEYINPUT5), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n268), .B1(new_n288), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n268), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT39), .B1(new_n291), .B2(new_n292), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n284), .B1(new_n280), .B2(new_n283), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT39), .ZN(new_n302));
  AOI211_X1 g101(.A(new_n298), .B(new_n301), .C1(new_n302), .C2(new_n300), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n297), .B1(new_n303), .B2(KEYINPUT40), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(KEYINPUT40), .B2(new_n303), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n309), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n311), .A2(KEYINPUT64), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(KEYINPUT64), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(G183gat), .A2(G190gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(KEYINPUT65), .B2(KEYINPUT24), .ZN(new_n317));
  AND2_X1   g116(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n318));
  OAI221_X1 g117(.A(new_n315), .B1(G183gat), .B2(G190gat), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(KEYINPUT25), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n322), .B(new_n315), .C1(G183gat), .C2(G190gat), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n314), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n320), .B1(new_n324), .B2(KEYINPUT25), .ZN(new_n325));
  XOR2_X1   g124(.A(KEYINPUT27), .B(G183gat), .Z(new_n326));
  INV_X1    g125(.A(KEYINPUT66), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT28), .ZN(new_n328));
  AOI211_X1 g127(.A(G190gat), .B(new_n326), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n329), .B1(new_n327), .B2(new_n328), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT26), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n308), .A2(new_n331), .A3(new_n306), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n332), .B(new_n316), .C1(new_n331), .C2(new_n308), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n333), .A2(new_n334), .ZN(new_n336));
  OAI211_X1 g135(.A(KEYINPUT66), .B(KEYINPUT28), .C1(new_n326), .C2(G190gat), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n330), .A2(new_n335), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n325), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(KEYINPUT29), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n339), .B2(new_n340), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n344), .A2(new_n234), .ZN(new_n345));
  OR2_X1    g144(.A1(new_n345), .A2(KEYINPUT74), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n234), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n347), .A3(KEYINPUT74), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n346), .A2(new_n348), .A3(new_n353), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT30), .ZN(new_n356));
  OR2_X1    g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n356), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OR2_X1    g158(.A1(new_n305), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n288), .A2(new_n268), .A3(new_n296), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OR2_X1    g162(.A1(new_n363), .A2(new_n297), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n297), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT37), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n355), .B1(new_n368), .B2(new_n352), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n345), .A2(new_n347), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT38), .B1(new_n370), .B2(KEYINPUT37), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n354), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT38), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n349), .A2(KEYINPUT37), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n374), .B1(new_n369), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT84), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n264), .B(new_n360), .C1(new_n373), .C2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n359), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n260), .B(new_n263), .C1(new_n367), .C2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n339), .B1(KEYINPUT69), .B2(new_n276), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n276), .A2(KEYINPUT69), .ZN(new_n382));
  OR2_X1    g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n382), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G227gat), .A2(G233gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT34), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n387), .B1(new_n386), .B2(KEYINPUT71), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n389), .B1(new_n385), .B2(new_n386), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n393), .A2(KEYINPUT70), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n383), .A2(G227gat), .A3(G233gat), .A4(new_n384), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT32), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g197(.A(G15gat), .B(G43gat), .Z(new_n399));
  XNOR2_X1  g198(.A(G71gat), .B(G99gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n396), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n401), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n395), .B(KEYINPUT32), .C1(new_n397), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n394), .B(new_n405), .Z(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT36), .ZN(new_n407));
  OR2_X1    g206(.A1(new_n405), .A2(new_n393), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n405), .A2(new_n393), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n411), .A2(KEYINPUT36), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n378), .A2(new_n380), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT35), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n406), .B1(new_n260), .B2(new_n263), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n365), .A2(new_n364), .B1(new_n357), .B2(new_n358), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n261), .A2(new_n262), .A3(new_n255), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n262), .B1(new_n261), .B2(new_n255), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n417), .A2(new_n415), .A3(new_n410), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n414), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G43gat), .B(G50gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(KEYINPUT89), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT15), .ZN(new_n427));
  OR3_X1    g226(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT90), .ZN(new_n431));
  INV_X1    g230(.A(G29gat), .ZN(new_n432));
  INV_X1    g231(.A(G36gat), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n427), .B(new_n431), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT91), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT88), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n429), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n429), .A2(new_n436), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n428), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n439), .B1(new_n432), .B2(new_n433), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(KEYINPUT15), .A3(new_n425), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(G15gat), .B(G22gat), .Z(new_n444));
  INV_X1    g243(.A(G8gat), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n444), .A2(G1gat), .B1(KEYINPUT92), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(G1gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT16), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n445), .A2(KEYINPUT92), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n443), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT93), .B1(new_n442), .B2(new_n451), .ZN(new_n454));
  XOR2_X1   g253(.A(new_n453), .B(new_n454), .Z(new_n455));
  NAND2_X1  g254(.A1(G229gat), .A2(G233gat), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n456), .B(KEYINPUT13), .Z(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n442), .B(KEYINPUT17), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n452), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n451), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n456), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT18), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n460), .A2(KEYINPUT18), .A3(new_n456), .A4(new_n461), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n458), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G113gat), .B(G141gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(KEYINPUT86), .ZN(new_n468));
  XNOR2_X1  g267(.A(G169gat), .B(G197gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n466), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n474), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n458), .A2(new_n464), .A3(new_n476), .A4(new_n465), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n424), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT100), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(G85gat), .A3(G92gat), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT7), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G99gat), .A2(G106gat), .ZN(new_n484));
  INV_X1    g283(.A(G85gat), .ZN(new_n485));
  INV_X1    g284(.A(G92gat), .ZN(new_n486));
  AOI22_X1  g285(.A1(KEYINPUT8), .A2(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n480), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n483), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G99gat), .B(G106gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n483), .A2(new_n487), .A3(new_n490), .A4(new_n488), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n493), .A2(KEYINPUT101), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(KEYINPUT101), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT102), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT101), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n489), .A2(new_n498), .A3(new_n490), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n493), .A2(KEYINPUT101), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT102), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n492), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n459), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G190gat), .B(G218gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n443), .B2(new_n502), .ZN(new_n506));
  OR3_X1    g305(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT103), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT99), .ZN(new_n511));
  INV_X1    g310(.A(G134gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(new_n204), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n504), .B1(new_n503), .B2(new_n506), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n509), .A2(new_n514), .B1(new_n507), .B2(new_n515), .ZN(new_n516));
  AND4_X1   g315(.A1(KEYINPUT103), .A2(new_n507), .A3(new_n515), .A4(new_n514), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G57gat), .B(G64gat), .Z(new_n520));
  INV_X1    g319(.A(G71gat), .ZN(new_n521));
  INV_X1    g320(.A(G78gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n520), .B1(KEYINPUT9), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g323(.A1(KEYINPUT94), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(G71gat), .B2(G78gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n524), .B(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(KEYINPUT95), .B(KEYINPUT21), .Z(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G231gat), .A2(G233gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G127gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(new_n203), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n533), .B(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n451), .B1(KEYINPUT21), .B2(new_n527), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n536), .B(new_n537), .Z(new_n538));
  XNOR2_X1  g337(.A(G183gat), .B(G211gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT98), .ZN(new_n540));
  XOR2_X1   g339(.A(KEYINPUT96), .B(KEYINPUT97), .Z(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n538), .B(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n519), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT107), .ZN(new_n546));
  NAND2_X1  g345(.A1(G230gat), .A2(G233gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT10), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n489), .A2(KEYINPUT105), .ZN(new_n550));
  INV_X1    g349(.A(new_n490), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n489), .A2(KEYINPUT105), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n499), .A2(new_n500), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(new_n527), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n524), .B(new_n526), .Z(new_n556));
  AOI21_X1  g355(.A(KEYINPUT104), .B1(new_n502), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n496), .B1(new_n494), .B2(new_n495), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n499), .A2(KEYINPUT102), .A3(new_n500), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n491), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT104), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n560), .A2(new_n561), .A3(new_n527), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n549), .B(new_n555), .C1(new_n557), .C2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n556), .A2(new_n549), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT106), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT106), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n560), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n548), .B1(new_n563), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n561), .B1(new_n560), .B2(new_n527), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n502), .A2(KEYINPUT104), .A3(new_n556), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n547), .B1(new_n573), .B2(new_n555), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G120gat), .B(G148gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(G176gat), .B(G204gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  AOI21_X1  g377(.A(new_n546), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(new_n575), .B2(new_n578), .ZN(new_n580));
  OR3_X1    g379(.A1(new_n575), .A2(KEYINPUT107), .A3(new_n578), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n545), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n479), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n585), .A2(new_n366), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(new_n447), .ZN(G1324gat));
  NOR2_X1   g386(.A1(new_n585), .A2(new_n359), .ZN(new_n588));
  XOR2_X1   g387(.A(KEYINPUT16), .B(G8gat), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n590), .B1(new_n445), .B2(new_n588), .ZN(new_n591));
  MUX2_X1   g390(.A(new_n590), .B(new_n591), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g391(.A(G15gat), .B1(new_n585), .B2(new_n413), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n411), .A2(G15gat), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n593), .B1(new_n585), .B2(new_n594), .ZN(G1326gat));
  NAND3_X1  g394(.A1(new_n479), .A2(new_n421), .A3(new_n584), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT108), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT43), .B(G22gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(G1327gat));
  INV_X1    g398(.A(new_n543), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n600), .A2(new_n518), .A3(new_n583), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n424), .A2(new_n478), .A3(new_n601), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n602), .A2(G29gat), .A3(new_n366), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n603), .B(KEYINPUT45), .Z(new_n604));
  INV_X1    g403(.A(KEYINPUT44), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n378), .A2(new_n380), .A3(new_n413), .ZN(new_n606));
  INV_X1    g405(.A(new_n406), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n607), .B(new_n417), .C1(new_n419), .C2(new_n420), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT35), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n264), .A2(new_n415), .A3(new_n417), .A4(new_n410), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(KEYINPUT109), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT109), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n612), .B1(new_n418), .B2(new_n423), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n606), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n605), .B1(new_n614), .B2(new_n518), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n424), .A2(KEYINPUT44), .A3(new_n519), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n478), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n600), .A2(new_n618), .A3(new_n583), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n617), .A2(new_n367), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n604), .B1(new_n620), .B2(new_n432), .ZN(G1328gat));
  NOR2_X1   g420(.A1(new_n359), .A2(G36gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n602), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT46), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n615), .A2(new_n379), .A3(new_n616), .A4(new_n619), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(G36gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT110), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(G1329gat));
  NOR3_X1   g429(.A1(new_n602), .A2(G43gat), .A3(new_n411), .ZN(new_n631));
  INV_X1    g430(.A(new_n413), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n615), .A2(new_n632), .A3(new_n616), .A4(new_n619), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n631), .B1(new_n633), .B2(G43gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g434(.A1(new_n615), .A2(new_n421), .A3(new_n616), .A4(new_n619), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(G50gat), .ZN(new_n637));
  INV_X1    g436(.A(G50gat), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n479), .A2(new_n638), .A3(new_n421), .A4(new_n601), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT48), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(G1331gat));
  NOR3_X1   g441(.A1(new_n545), .A2(new_n478), .A3(new_n582), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT111), .B1(new_n614), .B2(new_n644), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n418), .A2(new_n423), .A3(new_n612), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT109), .B1(new_n609), .B2(new_n610), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n414), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT111), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(new_n649), .A3(new_n643), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(new_n366), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(G57gat), .Z(G1332gat));
  AOI21_X1  g452(.A(new_n359), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n645), .A2(new_n650), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT112), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT112), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n645), .A2(new_n657), .A3(new_n650), .A4(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1333gat));
  OAI21_X1  g460(.A(G71gat), .B1(new_n651), .B2(new_n413), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n645), .A2(new_n521), .A3(new_n650), .A4(new_n410), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT50), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1334gat));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n264), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(new_n522), .ZN(G1335gat));
  NOR3_X1   g467(.A1(new_n600), .A2(new_n478), .A3(new_n582), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n617), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(G85gat), .B1(new_n670), .B2(new_n366), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n600), .A2(new_n478), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n648), .A2(new_n519), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT113), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT51), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n677));
  NAND4_X1  g476(.A1(new_n648), .A2(new_n519), .A3(new_n672), .A4(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n582), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n485), .A3(new_n367), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n671), .A2(new_n680), .ZN(G1336gat));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n678), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n359), .A2(new_n582), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n486), .A3(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n615), .A2(new_n379), .A3(new_n616), .A4(new_n669), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G92gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT52), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT52), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n684), .A2(new_n689), .A3(new_n686), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(G1337gat));
  OAI21_X1  g490(.A(G99gat), .B1(new_n670), .B2(new_n413), .ZN(new_n692));
  INV_X1    g491(.A(G99gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n679), .A2(new_n693), .A3(new_n410), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(G1338gat));
  INV_X1    g494(.A(KEYINPUT53), .ZN(new_n696));
  AOI21_X1  g495(.A(G106gat), .B1(new_n679), .B2(new_n421), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n421), .A2(G106gat), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n617), .A2(new_n669), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n696), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n617), .A2(new_n669), .A3(new_n698), .ZN(new_n701));
  AOI211_X1 g500(.A(new_n264), .B(new_n582), .C1(new_n676), .C2(new_n678), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n701), .B(KEYINPUT53), .C1(new_n702), .C2(G106gat), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(G1339gat));
  NAND2_X1  g503(.A1(new_n584), .A2(new_n618), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT54), .ZN(new_n707));
  INV_X1    g506(.A(new_n555), .ZN(new_n708));
  AOI211_X1 g507(.A(KEYINPUT10), .B(new_n708), .C1(new_n571), .C2(new_n572), .ZN(new_n709));
  INV_X1    g508(.A(new_n569), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n707), .B(new_n547), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n578), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n568), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n567), .B1(new_n560), .B2(new_n564), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n548), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT54), .B1(new_n709), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT114), .B1(new_n717), .B2(new_n570), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n547), .B1(new_n709), .B2(new_n710), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT114), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n547), .B1(new_n566), .B2(new_n568), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n707), .B1(new_n563), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n713), .B1(new_n718), .B2(new_n723), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n724), .A2(KEYINPUT55), .B1(new_n575), .B2(new_n578), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT115), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n724), .B2(KEYINPUT55), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n578), .B1(new_n570), .B2(new_n707), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n717), .A2(new_n570), .A3(KEYINPUT114), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n720), .B1(new_n719), .B2(new_n722), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT55), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n731), .A2(KEYINPUT115), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n725), .A2(new_n727), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT116), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT116), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n725), .A2(new_n727), .A3(new_n733), .A4(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n735), .A2(new_n478), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n455), .A2(new_n457), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n472), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n583), .A2(new_n477), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT117), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n738), .A2(KEYINPUT117), .A3(new_n742), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n518), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n741), .A2(new_n477), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n518), .A2(new_n748), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n735), .A2(new_n737), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n600), .B1(new_n752), .B2(KEYINPUT118), .ZN(new_n753));
  INV_X1    g552(.A(new_n751), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n519), .B1(new_n743), .B2(new_n744), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n755), .B2(new_n746), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT118), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n706), .B1(new_n753), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n366), .ZN(new_n760));
  INV_X1    g559(.A(new_n416), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n379), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(G113gat), .B1(new_n763), .B2(new_n478), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT119), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n759), .B2(new_n421), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n543), .B1(new_n756), .B2(new_n757), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n747), .A2(new_n757), .A3(new_n751), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n705), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n769), .A2(KEYINPUT119), .A3(new_n264), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n379), .A2(new_n366), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n411), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n478), .A2(G113gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n764), .B1(new_n775), .B2(new_n776), .ZN(G1340gat));
  AOI21_X1  g576(.A(G120gat), .B1(new_n763), .B2(new_n583), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n583), .A2(G120gat), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n775), .B2(new_n779), .ZN(G1341gat));
  NAND3_X1  g579(.A1(new_n771), .A2(new_n600), .A3(new_n774), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G127gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n763), .A2(new_n532), .A3(new_n600), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1342gat));
  NAND4_X1  g583(.A1(new_n760), .A2(new_n512), .A3(new_n519), .A4(new_n762), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n770), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT119), .B1(new_n769), .B2(new_n264), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n519), .B(new_n774), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT120), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n790), .A2(new_n791), .A3(G134gat), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n790), .B2(G134gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n787), .B1(new_n792), .B2(new_n793), .ZN(G1343gat));
  NOR2_X1   g593(.A1(new_n632), .A2(new_n773), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT57), .B1(new_n769), .B2(new_n421), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n421), .A2(KEYINPUT57), .ZN(new_n797));
  XNOR2_X1  g596(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n478), .B(new_n725), .C1(new_n724), .C2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n519), .B1(new_n799), .B2(new_n742), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n543), .B1(new_n754), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n797), .B1(new_n705), .B2(new_n801), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n478), .B(new_n795), .C1(new_n796), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G141gat), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n632), .A2(new_n379), .A3(new_n264), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n618), .A2(G141gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n760), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT58), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n804), .A2(new_n810), .A3(new_n807), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1344gat));
  NOR2_X1   g611(.A1(new_n759), .A2(new_n797), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n518), .A2(new_n748), .A3(new_n734), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n543), .B1(new_n800), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n705), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT57), .B1(new_n816), .B2(new_n421), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n795), .A2(new_n583), .ZN(new_n819));
  OAI211_X1 g618(.A(KEYINPUT59), .B(G148gat), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n795), .B1(new_n796), .B2(new_n802), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT59), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n583), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n760), .A2(new_n805), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n822), .B1(new_n825), .B2(new_n583), .ZN(new_n826));
  OAI221_X1 g625(.A(new_n820), .B1(new_n821), .B2(new_n823), .C1(new_n826), .C2(G148gat), .ZN(G1345gat));
  NOR3_X1   g626(.A1(new_n824), .A2(KEYINPUT122), .A3(new_n543), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(G155gat), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT122), .B1(new_n824), .B2(new_n543), .ZN(new_n830));
  INV_X1    g629(.A(new_n821), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n543), .A2(new_n203), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n829), .A2(new_n830), .B1(new_n831), .B2(new_n832), .ZN(G1346gat));
  AOI21_X1  g632(.A(G162gat), .B1(new_n825), .B2(new_n519), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n518), .A2(new_n204), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n831), .B2(new_n835), .ZN(G1347gat));
  NOR2_X1   g635(.A1(new_n759), .A2(new_n367), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n761), .A2(new_n359), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n618), .A2(G169gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT123), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n379), .A2(new_n366), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n411), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n766), .B2(new_n770), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n478), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(G169gat), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n841), .A2(new_n847), .ZN(G1348gat));
  NAND4_X1  g647(.A1(new_n771), .A2(G176gat), .A3(new_n583), .A4(new_n843), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT124), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n845), .A2(KEYINPUT124), .A3(G176gat), .A4(new_n583), .ZN(new_n852));
  INV_X1    g651(.A(G176gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n582), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n851), .A2(new_n852), .A3(new_n855), .ZN(G1349gat));
  INV_X1    g655(.A(G183gat), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n845), .B2(new_n600), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n543), .A2(new_n326), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n837), .A2(new_n838), .A3(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT60), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n600), .B(new_n843), .C1(new_n788), .C2(new_n789), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(G183gat), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n865), .A3(new_n860), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n862), .A2(new_n866), .ZN(G1350gat));
  OR3_X1    g666(.A1(new_n854), .A2(G190gat), .A3(new_n518), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n519), .B(new_n843), .C1(new_n788), .C2(new_n789), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT61), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n869), .A2(new_n870), .A3(G190gat), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n869), .B2(G190gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(G1351gat));
  INV_X1    g672(.A(KEYINPUT126), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n632), .A2(new_n264), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n837), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  XOR2_X1   g676(.A(KEYINPUT125), .B(G197gat), .Z(new_n878));
  NOR2_X1   g677(.A1(new_n618), .A2(new_n878), .ZN(new_n879));
  AND4_X1   g678(.A1(new_n874), .A2(new_n877), .A3(new_n379), .A4(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n818), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n632), .A2(new_n842), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n478), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n878), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n876), .A2(new_n359), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n874), .B1(new_n885), .B2(new_n879), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n880), .B1(new_n884), .B2(new_n886), .ZN(G1352gat));
  NAND3_X1  g686(.A1(new_n881), .A2(new_n583), .A3(new_n882), .ZN(new_n888));
  XNOR2_X1  g687(.A(KEYINPUT127), .B(G204gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OR3_X1    g689(.A1(new_n359), .A2(new_n582), .A3(new_n889), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT62), .B1(new_n876), .B2(new_n891), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n876), .A2(KEYINPUT62), .A3(new_n891), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(G1353gat));
  NAND3_X1  g693(.A1(new_n885), .A2(new_n225), .A3(new_n600), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n600), .B(new_n882), .C1(new_n813), .C2(new_n817), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n896), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT63), .B1(new_n896), .B2(G211gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(G1354gat));
  NAND3_X1  g698(.A1(new_n885), .A2(new_n226), .A3(new_n519), .ZN(new_n900));
  NOR4_X1   g699(.A1(new_n818), .A2(new_n632), .A3(new_n518), .A4(new_n842), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n226), .ZN(G1355gat));
endmodule


