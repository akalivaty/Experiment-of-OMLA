//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT77), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT77), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  AOI21_X1  g004(.A(G107), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT79), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  OAI22_X1  g007(.A1(new_n191), .A2(new_n192), .B1(G104), .B2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n189), .A2(G104), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n187), .A2(KEYINPUT77), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n193), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT79), .ZN(new_n198));
  OAI21_X1  g012(.A(G101), .B1(new_n194), .B2(new_n198), .ZN(new_n199));
  XOR2_X1   g013(.A(G116), .B(G119), .Z(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT5), .ZN(new_n202));
  INV_X1    g016(.A(G113), .ZN(new_n203));
  INV_X1    g017(.A(G116), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT5), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT2), .A2(G113), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT2), .A2(G113), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n208), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n202), .A2(new_n207), .B1(new_n213), .B2(new_n201), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n187), .A2(KEYINPUT3), .A3(G107), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n215), .B1(new_n197), .B2(KEYINPUT3), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n188), .A2(new_n190), .A3(G107), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n199), .A2(new_n214), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n200), .A2(KEYINPUT69), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n221), .B(new_n213), .ZN(new_n222));
  INV_X1    g036(.A(new_n215), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n218), .B(new_n223), .C1(new_n191), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G101), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n223), .B1(new_n191), .B2(new_n224), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n218), .A2(new_n217), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT4), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n222), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT78), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n217), .A2(KEYINPUT4), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n225), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n232), .B1(new_n225), .B2(new_n233), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n220), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(G110), .B(G122), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n238), .B(new_n220), .C1(new_n231), .C2(new_n236), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(KEYINPUT6), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n243));
  INV_X1    g057(.A(G146), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(G143), .ZN(new_n245));
  INV_X1    g059(.A(G143), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT65), .A3(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(G143), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G128), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n249), .A2(KEYINPUT1), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n253), .B1(G143), .B2(new_n244), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(G128), .A3(new_n258), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n246), .A2(KEYINPUT64), .A3(G146), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT64), .B1(new_n246), .B2(G146), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n249), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n252), .A2(new_n253), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G125), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n245), .A2(new_n247), .B1(G143), .B2(new_n244), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT0), .A3(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT66), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT66), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n266), .A2(new_n269), .A3(KEYINPUT0), .A4(G128), .ZN(new_n270));
  XOR2_X1   g084(.A(KEYINPUT0), .B(G128), .Z(new_n271));
  AOI22_X1  g085(.A1(new_n268), .A2(new_n270), .B1(new_n262), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n265), .B1(new_n272), .B2(new_n264), .ZN(new_n273));
  INV_X1    g087(.A(G224), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G953), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT82), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n273), .B(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n237), .A2(new_n278), .A3(new_n239), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n242), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT83), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n242), .A2(new_n277), .A3(KEYINPUT83), .A4(new_n279), .ZN(new_n283));
  INV_X1    g097(.A(new_n241), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n199), .A2(new_n219), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n214), .ZN(new_n286));
  XOR2_X1   g100(.A(new_n238), .B(KEYINPUT8), .Z(new_n287));
  NAND2_X1  g101(.A1(new_n201), .A2(new_n213), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n202), .B(KEYINPUT84), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n207), .B(KEYINPUT85), .Z(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n199), .A2(new_n219), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n287), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n284), .B1(new_n286), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n275), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n273), .B(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n282), .A2(new_n283), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G210), .B1(G237), .B2(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n282), .A2(new_n298), .A3(new_n300), .A4(new_n283), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G214), .B1(G237), .B2(G902), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n299), .A2(KEYINPUT86), .A3(new_n301), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT87), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT87), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n305), .A2(new_n310), .A3(new_n306), .A4(new_n307), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT9), .B(G234), .ZN(new_n313));
  OAI21_X1  g127(.A(G221), .B1(new_n313), .B2(G902), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G469), .ZN(new_n316));
  INV_X1    g130(.A(G902), .ZN(new_n317));
  XNOR2_X1  g131(.A(G110), .B(G140), .ZN(new_n318));
  INV_X1    g132(.A(G953), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G227), .ZN(new_n320));
  XOR2_X1   g134(.A(new_n318), .B(new_n320), .Z(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n259), .A2(new_n262), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n266), .A2(new_n253), .A3(G128), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n292), .A2(KEYINPUT10), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n219), .A2(new_n226), .A3(KEYINPUT4), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n272), .B(new_n327), .C1(new_n234), .C2(new_n235), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n257), .A2(KEYINPUT80), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G128), .B1(new_n257), .B2(KEYINPUT80), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n250), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n324), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n199), .A3(new_n219), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT10), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n326), .A2(new_n328), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT81), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT11), .ZN(new_n339));
  INV_X1    g153(.A(G134), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(G137), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(G137), .ZN(new_n342));
  INV_X1    g156(.A(G137), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(KEYINPUT11), .A3(G134), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G131), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n326), .A2(new_n328), .A3(new_n349), .A4(new_n336), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n338), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n326), .A2(new_n328), .A3(new_n347), .A4(new_n336), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n322), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n285), .A2(new_n263), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n334), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT12), .B1(new_n355), .B2(new_n348), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT12), .ZN(new_n357));
  AOI211_X1 g171(.A(new_n357), .B(new_n347), .C1(new_n354), .C2(new_n334), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n352), .A2(new_n322), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n316), .B(new_n317), .C1(new_n353), .C2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n360), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n352), .B1(new_n356), .B2(new_n358), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n351), .A2(new_n363), .B1(new_n364), .B2(new_n321), .ZN(new_n365));
  OAI21_X1  g179(.A(G469), .B1(new_n365), .B2(G902), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n315), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G237), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n319), .A3(G214), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n246), .ZN(new_n370));
  NOR2_X1   g184(.A1(G237), .A2(G953), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(G143), .A3(G214), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n346), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT17), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT16), .ZN(new_n375));
  INV_X1    g189(.A(G140), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(G125), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(G125), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n264), .A2(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n377), .B1(new_n380), .B2(new_n375), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n244), .ZN(new_n382));
  OAI211_X1 g196(.A(G146), .B(new_n377), .C1(new_n380), .C2(new_n375), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n374), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n370), .A2(new_n346), .A3(new_n372), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n386), .A2(KEYINPUT17), .A3(new_n373), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G113), .B(G122), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(new_n187), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT89), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n380), .A2(KEYINPUT74), .A3(G146), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT74), .ZN(new_n394));
  XNOR2_X1  g208(.A(G125), .B(G140), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n394), .B1(new_n395), .B2(new_n244), .ZN(new_n396));
  OAI22_X1  g210(.A1(new_n393), .A2(new_n396), .B1(new_n244), .B2(new_n395), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n370), .A2(new_n372), .ZN(new_n398));
  AND2_X1   g212(.A1(KEYINPUT18), .A2(G131), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n399), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n388), .A2(new_n392), .A3(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n395), .A2(KEYINPUT19), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n395), .A2(KEYINPUT19), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n244), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n406), .B(new_n383), .C1(new_n373), .C2(new_n386), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n402), .ZN(new_n408));
  INV_X1    g222(.A(new_n390), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT88), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT88), .ZN(new_n411));
  AOI211_X1 g225(.A(new_n411), .B(new_n390), .C1(new_n407), .C2(new_n402), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n403), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(G475), .A2(G902), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT20), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n390), .B1(new_n388), .B2(new_n402), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n402), .B1(new_n387), .B2(new_n384), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(new_n391), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n317), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n415), .A2(new_n416), .B1(G475), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n413), .A2(KEYINPUT90), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT90), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n423), .B(new_n403), .C1(new_n410), .C2(new_n412), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n422), .A2(KEYINPUT20), .A3(new_n414), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n251), .A2(G143), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  XOR2_X1   g243(.A(G128), .B(G143), .Z(new_n430));
  OAI211_X1 g244(.A(new_n429), .B(G134), .C1(new_n427), .C2(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(G116), .B(G122), .Z(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G107), .ZN(new_n433));
  XNOR2_X1  g247(.A(G116), .B(G122), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n193), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G128), .B(G143), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n340), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n431), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n430), .A2(G134), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n438), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n204), .A2(KEYINPUT14), .A3(G122), .ZN(new_n442));
  OAI211_X1 g256(.A(G107), .B(new_n442), .C1(new_n432), .C2(KEYINPUT14), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n435), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G217), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n313), .A2(new_n445), .A3(G953), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n439), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n446), .B1(new_n439), .B2(new_n444), .ZN(new_n449));
  OAI211_X1 g263(.A(KEYINPUT93), .B(new_n317), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G478), .B1(KEYINPUT92), .B2(KEYINPUT15), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(KEYINPUT92), .B2(KEYINPUT15), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n439), .A2(new_n444), .ZN(new_n454));
  INV_X1    g268(.A(new_n446), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n447), .ZN(new_n457));
  INV_X1    g271(.A(new_n452), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n457), .A2(KEYINPUT93), .A3(new_n317), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT94), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n453), .A2(new_n459), .A3(KEYINPUT94), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(G234), .A2(G237), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(G952), .A3(new_n319), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(G902), .A3(G953), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(G898), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n426), .A2(new_n464), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n367), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n312), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT95), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n345), .A2(G131), .ZN(new_n478));
  INV_X1    g292(.A(new_n342), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n340), .A2(G137), .ZN(new_n480));
  OAI21_X1  g294(.A(G131), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT70), .B1(new_n263), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n482), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT70), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n325), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n268), .A2(new_n270), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n262), .A2(new_n271), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n348), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n222), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n483), .A2(new_n486), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT26), .B(G101), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n371), .A2(G210), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT72), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT72), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n491), .A2(new_n499), .A3(new_n496), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n484), .A2(new_n325), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n489), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n483), .A2(new_n486), .A3(new_n489), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n504), .B1(KEYINPUT30), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n498), .B(new_n500), .C1(new_n506), .C2(new_n490), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT31), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT28), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n489), .A2(new_n502), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n222), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n222), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n511), .B(new_n512), .C1(new_n509), .C2(new_n491), .ZN(new_n513));
  INV_X1    g327(.A(new_n496), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n505), .A2(KEYINPUT30), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n503), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n222), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT31), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n518), .A2(new_n519), .A3(new_n500), .A4(new_n498), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n508), .A2(new_n515), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(G472), .A2(G902), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(KEYINPUT32), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT73), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n522), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT32), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT73), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n521), .A2(new_n528), .A3(KEYINPUT32), .A4(new_n522), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n505), .A2(new_n222), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n509), .B1(new_n530), .B2(new_n491), .ZN(new_n531));
  INV_X1    g345(.A(new_n511), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(KEYINPUT29), .A3(new_n496), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n317), .ZN(new_n535));
  INV_X1    g349(.A(new_n491), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n517), .B2(new_n222), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(new_n496), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT29), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n513), .B2(new_n514), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G472), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n524), .A2(new_n527), .A3(new_n529), .A4(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n382), .A2(new_n383), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n206), .A2(G128), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n251), .A2(KEYINPUT23), .A3(G119), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n206), .A2(G128), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n546), .B(new_n547), .C1(new_n548), .C2(KEYINPUT23), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n251), .A2(G119), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n550), .A2(new_n546), .ZN(new_n551));
  XOR2_X1   g365(.A(KEYINPUT24), .B(G110), .Z(new_n552));
  AOI22_X1  g366(.A1(new_n549), .A2(G110), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n545), .A2(new_n553), .ZN(new_n554));
  OAI22_X1  g368(.A1(new_n549), .A2(G110), .B1(new_n551), .B2(new_n552), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n555), .B(new_n383), .C1(new_n393), .C2(new_n396), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT22), .B(G137), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT75), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n319), .A2(G221), .A3(G234), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n557), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n317), .ZN(new_n563));
  NOR2_X1   g377(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n567), .B1(new_n563), .B2(new_n564), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n445), .B1(G234), .B2(new_n317), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(G902), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n562), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n544), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n312), .A2(KEYINPUT95), .A3(new_n474), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n477), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(G101), .ZN(G3));
  INV_X1    g392(.A(G472), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n521), .B2(new_n317), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n525), .ZN(new_n582));
  INV_X1    g396(.A(new_n367), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n582), .A2(new_n574), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n302), .A2(new_n304), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n306), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(new_n471), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT96), .B(KEYINPUT33), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n455), .A2(KEYINPUT97), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n439), .A2(new_n444), .A3(new_n590), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n591), .A2(KEYINPUT33), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n454), .A2(KEYINPUT97), .A3(new_n455), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n457), .A2(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(G478), .A3(new_n317), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n456), .B2(new_n447), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n595), .B1(G478), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n426), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n588), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n585), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT34), .B(G104), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G6));
  NAND3_X1  g417(.A1(new_n422), .A2(new_n414), .A3(new_n424), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n416), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n605), .A2(new_n425), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n418), .A2(new_n409), .ZN(new_n607));
  AOI21_X1  g421(.A(G902), .B1(new_n403), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(G475), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT98), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n420), .A2(new_n611), .A3(G475), .ZN(new_n612));
  AND4_X1   g426(.A1(new_n462), .A2(new_n463), .A3(new_n610), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n588), .A2(new_n606), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n585), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT35), .B(G107), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT99), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n615), .B(new_n617), .ZN(G9));
  INV_X1    g432(.A(new_n570), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n565), .B2(new_n568), .ZN(new_n620));
  INV_X1    g434(.A(new_n561), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(KEYINPUT36), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(new_n557), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n572), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT100), .B1(new_n620), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n571), .A2(new_n627), .A3(new_n624), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n582), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n477), .A2(new_n576), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT37), .B(G110), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT101), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n630), .B(new_n632), .ZN(G12));
  NOR2_X1   g447(.A1(new_n583), .A2(new_n587), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT102), .B(G900), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n469), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n466), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n606), .A2(new_n635), .A3(new_n613), .A4(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n613), .A2(new_n425), .A3(new_n605), .A4(new_n638), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT103), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n628), .A2(new_n626), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n639), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n634), .A2(new_n643), .A3(new_n543), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G128), .ZN(G30));
  INV_X1    g459(.A(new_n507), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n496), .B1(new_n530), .B2(new_n491), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n317), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(G472), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n524), .A2(new_n527), .A3(new_n529), .A4(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n650), .B(KEYINPUT104), .Z(new_n651));
  NAND2_X1  g465(.A1(new_n305), .A2(new_n307), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(KEYINPUT38), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n638), .B(KEYINPUT39), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n367), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n655), .B(KEYINPUT40), .Z(new_n656));
  INV_X1    g470(.A(new_n306), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n426), .A2(new_n464), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n642), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n651), .A2(new_n653), .A3(new_n656), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT105), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G143), .ZN(G45));
  NAND3_X1  g476(.A1(new_n426), .A2(new_n597), .A3(new_n638), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n634), .A2(new_n543), .A3(new_n642), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G146), .ZN(G48));
  NOR2_X1   g480(.A1(new_n353), .A2(new_n361), .ZN(new_n667));
  OAI21_X1  g481(.A(G469), .B1(new_n667), .B2(G902), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n668), .A2(new_n314), .A3(new_n362), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT106), .ZN(new_n670));
  INV_X1    g484(.A(new_n574), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n668), .A2(new_n672), .A3(new_n314), .A4(new_n362), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n543), .A2(new_n670), .A3(new_n671), .A4(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n600), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT41), .B(G113), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  NOR2_X1   g491(.A1(new_n674), .A2(new_n614), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n204), .ZN(G18));
  NOR2_X1   g493(.A1(new_n587), .A2(new_n669), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n680), .A2(new_n543), .A3(new_n472), .A4(new_n642), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G119), .ZN(G21));
  NOR3_X1   g496(.A1(new_n587), .A2(new_n471), .A3(new_n658), .ZN(new_n683));
  INV_X1    g497(.A(new_n522), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n508), .A2(new_n520), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n496), .B1(new_n533), .B2(KEYINPUT107), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(KEYINPUT107), .B2(new_n533), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n684), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n688), .A2(new_n580), .A3(new_n574), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n683), .A2(new_n670), .A3(new_n673), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G122), .ZN(G24));
  NOR3_X1   g505(.A1(new_n688), .A2(new_n580), .A3(new_n663), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n680), .A2(new_n642), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n657), .B1(new_n305), .B2(new_n307), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n543), .A2(new_n671), .A3(new_n696), .A4(new_n367), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n695), .B1(new_n697), .B2(new_n663), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n527), .A2(new_n542), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n574), .B1(new_n699), .B2(new_n523), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n696), .A2(new_n367), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n700), .A2(new_n702), .A3(KEYINPUT42), .A4(new_n664), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G131), .ZN(G33));
  NAND2_X1  g519(.A1(new_n639), .A2(new_n641), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n697), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n340), .ZN(G36));
  OR2_X1    g522(.A1(new_n365), .A2(KEYINPUT45), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n365), .A2(KEYINPUT45), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(G469), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(G469), .A2(G902), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(KEYINPUT46), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n362), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n714), .A2(KEYINPUT108), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n711), .A2(new_n712), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n714), .A2(KEYINPUT108), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n719), .A2(new_n314), .A3(new_n654), .ZN(new_n720));
  INV_X1    g534(.A(new_n426), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n597), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n582), .A3(new_n642), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  INV_X1    g542(.A(new_n696), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n720), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G137), .ZN(G39));
  NOR4_X1   g546(.A1(new_n729), .A2(new_n543), .A3(new_n671), .A4(new_n663), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT109), .ZN(new_n734));
  INV_X1    g548(.A(new_n719), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT47), .B1(new_n735), .B2(new_n315), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n719), .A2(new_n737), .A3(new_n314), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n734), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G140), .ZN(G42));
  NAND2_X1  g554(.A1(new_n724), .A2(new_n467), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n743), .A2(new_n689), .ZN(new_n744));
  INV_X1    g558(.A(new_n653), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n669), .A2(new_n306), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(KEYINPUT50), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n743), .A2(new_n689), .A3(new_n746), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n748), .B1(new_n749), .B2(new_n653), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n729), .A2(new_n669), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n671), .A3(new_n467), .ZN(new_n754));
  OR4_X1    g568(.A1(new_n426), .A2(new_n754), .A3(new_n597), .A4(new_n651), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n743), .A2(new_n753), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n688), .A2(new_n580), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n642), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n751), .A2(new_n755), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n744), .A2(new_n696), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n736), .A2(new_n738), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n668), .A2(new_n315), .A3(new_n362), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n764));
  OR3_X1    g578(.A1(new_n759), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n764), .B1(new_n759), .B2(new_n763), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n756), .A2(new_n700), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n767), .B(KEYINPUT48), .Z(new_n768));
  INV_X1    g582(.A(G952), .ZN(new_n769));
  AOI211_X1 g583(.A(new_n769), .B(G953), .C1(new_n744), .C2(new_n680), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n754), .A2(new_n651), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n770), .B1(new_n598), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n765), .A2(new_n766), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n721), .A2(new_n460), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n471), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n312), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT112), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n312), .A2(new_n779), .A3(new_n776), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n778), .A2(new_n584), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n471), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n312), .A2(new_n584), .A3(new_n782), .A4(new_n599), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n577), .A2(new_n630), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT113), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT95), .B1(new_n312), .B2(new_n474), .ZN(new_n786));
  AOI211_X1 g600(.A(new_n476), .B(new_n473), .C1(new_n309), .C2(new_n311), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n585), .B1(new_n777), .B2(KEYINPUT112), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n788), .A2(new_n629), .B1(new_n789), .B2(new_n780), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n791));
  INV_X1    g605(.A(new_n783), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n788), .B2(new_n575), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n785), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n644), .A2(new_n693), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n587), .A2(new_n658), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n620), .A2(new_n625), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n367), .A2(new_n798), .A3(new_n638), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(new_n650), .A3(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n796), .A2(KEYINPUT52), .A3(new_n665), .A4(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n665), .A2(new_n644), .A3(new_n800), .A4(new_n693), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n690), .B(new_n681), .C1(new_n674), .C2(new_n600), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n460), .B1(new_n466), .B2(new_n637), .ZN(new_n807));
  AND4_X1   g621(.A1(new_n606), .A2(new_n610), .A3(new_n612), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n692), .B1(new_n543), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n696), .A2(new_n367), .A3(new_n642), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n806), .A2(new_n678), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n707), .B1(new_n698), .B2(new_n703), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n805), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT53), .B1(new_n795), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n817));
  AOI211_X1 g631(.A(new_n817), .B(new_n814), .C1(new_n785), .C2(new_n794), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT54), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n784), .A2(KEYINPUT113), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n791), .B1(new_n790), .B2(new_n793), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n815), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n817), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n795), .A2(KEYINPUT53), .A3(new_n815), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n774), .A2(new_n819), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT115), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n774), .A2(new_n829), .A3(new_n819), .A4(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n769), .A2(new_n319), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n574), .A2(new_n657), .A3(new_n315), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT110), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n668), .A2(new_n362), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n722), .B(new_n834), .C1(KEYINPUT49), .C2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(KEYINPUT49), .B2(new_n835), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n837), .A2(new_n651), .A3(new_n653), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n838), .B(KEYINPUT111), .Z(new_n839));
  NAND2_X1  g653(.A1(new_n832), .A2(new_n839), .ZN(G75));
  NOR2_X1   g654(.A1(new_n319), .A2(G952), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n317), .B1(new_n823), .B2(new_n825), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT56), .B1(new_n843), .B2(G210), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n242), .A2(new_n279), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(new_n277), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT55), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n842), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n823), .A2(new_n825), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(G210), .A3(G902), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT116), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n843), .A2(new_n852), .A3(G210), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT56), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n851), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n851), .A2(KEYINPUT117), .A3(new_n853), .A4(new_n855), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n848), .B1(new_n858), .B2(new_n859), .ZN(G51));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n711), .B(KEYINPUT120), .ZN(new_n862));
  OAI211_X1 g676(.A(G902), .B(new_n862), .C1(new_n816), .C2(new_n818), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n712), .B(KEYINPUT118), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT57), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n816), .A2(new_n818), .A3(KEYINPUT54), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n824), .B1(new_n823), .B2(new_n825), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n667), .B(KEYINPUT119), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n864), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n861), .B1(new_n871), .B2(new_n841), .ZN(new_n872));
  INV_X1    g686(.A(new_n870), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n819), .A2(new_n826), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n873), .B1(new_n874), .B2(new_n866), .ZN(new_n875));
  OAI211_X1 g689(.A(KEYINPUT121), .B(new_n842), .C1(new_n875), .C2(new_n864), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n872), .A2(new_n876), .ZN(G54));
  NAND2_X1  g691(.A1(KEYINPUT58), .A2(G475), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT122), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n843), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n422), .A2(new_n424), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n842), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n881), .B2(new_n880), .ZN(G60));
  NAND2_X1  g697(.A1(G478), .A2(G902), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT59), .Z(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(new_n819), .B2(new_n826), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n842), .B1(new_n886), .B2(new_n594), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n594), .B2(new_n886), .ZN(G63));
  NAND2_X1  g702(.A1(G217), .A2(G902), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT60), .Z(new_n890));
  NAND3_X1  g704(.A1(new_n849), .A2(new_n623), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n849), .A2(new_n890), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n842), .B(new_n891), .C1(new_n892), .C2(new_n562), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n893), .B(new_n894), .ZN(G66));
  NOR3_X1   g709(.A1(new_n470), .A2(new_n274), .A3(new_n319), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n806), .A2(new_n678), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n795), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n896), .B1(new_n899), .B2(new_n319), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n845), .B1(G898), .B2(new_n319), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n900), .B(new_n901), .ZN(G69));
  NOR2_X1   g716(.A1(new_n404), .A2(new_n405), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n506), .B(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n660), .A2(new_n665), .A3(new_n796), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT62), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT123), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n775), .A2(new_n598), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT124), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n575), .A2(new_n654), .A3(new_n702), .A4(new_n909), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n739), .A2(new_n731), .A3(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n907), .B(new_n911), .C1(KEYINPUT62), .C2(new_n905), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n904), .B1(new_n912), .B2(new_n319), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n731), .A2(new_n665), .A3(new_n796), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n720), .A2(new_n797), .A3(new_n700), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n914), .A2(new_n915), .A3(new_n739), .A4(new_n813), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(G953), .ZN(new_n917));
  NAND2_X1  g731(.A1(G900), .A2(G953), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n904), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n913), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n319), .B1(G227), .B2(G900), .ZN(new_n922));
  INV_X1    g736(.A(new_n920), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n922), .B1(new_n923), .B2(KEYINPUT125), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n921), .B(new_n924), .ZN(G72));
  XNOR2_X1  g739(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n579), .A2(new_n317), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n849), .B(new_n928), .C1(new_n646), .C2(new_n538), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT127), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n912), .B2(new_n898), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n537), .A2(new_n514), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n928), .B1(new_n898), .B2(new_n916), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n934), .A2(new_n514), .A3(new_n537), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n842), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n930), .A2(new_n936), .ZN(G57));
endmodule


