//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT80), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  INV_X1    g006(.A(G227), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G953), .ZN(new_n194));
  XOR2_X1   g008(.A(new_n192), .B(new_n194), .Z(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT79), .A2(KEYINPUT12), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT12), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n201), .A2(new_n203), .A3(new_n204), .A4(G128), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n206), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n207));
  XNOR2_X1  g021(.A(G143), .B(G146), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n205), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G104), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(G107), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n211), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(G104), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT77), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G101), .ZN(new_n221));
  XNOR2_X1  g035(.A(G104), .B(G107), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT77), .B1(new_n222), .B2(new_n215), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n209), .A2(new_n217), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n221), .A3(new_n217), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n201), .A2(new_n203), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n228), .B(KEYINPUT1), .C1(new_n202), .C2(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G128), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n228), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n227), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n205), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n224), .B1(new_n226), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G131), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(KEYINPUT66), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT11), .A2(G134), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT65), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G137), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n237), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(G137), .ZN(new_n243));
  OR2_X1    g057(.A1(KEYINPUT11), .A2(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n236), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT11), .A2(G134), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(G137), .B2(new_n237), .ZN(new_n248));
  INV_X1    g062(.A(new_n236), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT65), .B(G137), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n248), .B(new_n249), .C1(new_n237), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  AOI211_X1 g066(.A(new_n196), .B(new_n199), .C1(new_n234), .C2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n234), .A2(new_n197), .A3(new_n198), .A4(new_n252), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT10), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n224), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n211), .A2(new_n214), .A3(new_n216), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G101), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT0), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(new_n206), .ZN(new_n264));
  NOR3_X1   g078(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n227), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n208), .B1(new_n263), .B2(new_n206), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n259), .A2(new_n269), .A3(G101), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n261), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n258), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT78), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n225), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n223), .A2(new_n221), .A3(KEYINPUT78), .A4(new_n217), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT10), .A3(new_n233), .ZN(new_n278));
  INV_X1    g092(.A(new_n252), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n273), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n195), .B1(new_n256), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n280), .ZN(new_n282));
  INV_X1    g096(.A(new_n195), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n279), .B1(new_n273), .B2(new_n278), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n191), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n199), .B1(new_n234), .B2(new_n252), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(KEYINPUT79), .B2(KEYINPUT12), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n280), .A3(new_n254), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n283), .ZN(new_n290));
  INV_X1    g104(.A(new_n284), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(new_n280), .A3(new_n195), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(KEYINPUT80), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n286), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G469), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n256), .A2(new_n280), .A3(new_n195), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n283), .B1(new_n282), .B2(new_n284), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G469), .ZN(new_n300));
  OR2_X1    g114(.A1(new_n300), .A2(KEYINPUT81), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(KEYINPUT81), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n299), .A2(new_n294), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n190), .B1(new_n296), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT88), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT86), .ZN(new_n306));
  INV_X1    g120(.A(G237), .ZN(new_n307));
  INV_X1    g121(.A(G953), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(G214), .ZN(new_n309));
  NOR2_X1   g123(.A1(KEYINPUT85), .A2(G143), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(G237), .A2(G953), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n312), .B(G214), .C1(KEYINPUT85), .C2(G143), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n306), .B1(new_n314), .B2(G131), .ZN(new_n315));
  AOI211_X1 g129(.A(KEYINPUT86), .B(new_n235), .C1(new_n311), .C2(new_n313), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT17), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G125), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n319), .A2(KEYINPUT16), .A3(G140), .ZN(new_n320));
  XNOR2_X1  g134(.A(G125), .B(G140), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(KEYINPUT16), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(G146), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n305), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n314), .A2(G131), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT86), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n314), .A2(new_n306), .A3(G131), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n314), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n235), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n317), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n322), .B(new_n200), .ZN(new_n332));
  OAI211_X1 g146(.A(KEYINPUT88), .B(new_n332), .C1(new_n328), .C2(new_n317), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n324), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G113), .B(G122), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(new_n210), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT18), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n329), .B1(new_n337), .B2(new_n235), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n321), .B(new_n200), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n338), .B(new_n339), .C1(new_n337), .C2(new_n325), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n334), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n322), .A2(G146), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT19), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n321), .B(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n342), .B1(new_n344), .B2(G146), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT87), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(KEYINPUT87), .B(new_n342), .C1(new_n344), .C2(G146), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n328), .A2(new_n330), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n340), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n336), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n341), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT20), .ZN(new_n355));
  NOR2_X1   g169(.A1(G475), .A2(G902), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(KEYINPUT90), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT89), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n341), .A2(new_n360), .A3(new_n353), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n341), .B2(new_n353), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n357), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n359), .B1(new_n363), .B2(KEYINPUT20), .ZN(new_n364));
  INV_X1    g178(.A(new_n341), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n336), .B1(new_n334), .B2(new_n340), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n294), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G475), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n206), .A2(G143), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n206), .A2(G143), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G134), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G116), .B(G122), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(new_n213), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n370), .B1(new_n372), .B2(KEYINPUT13), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT91), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n372), .A2(KEYINPUT13), .ZN(new_n381));
  OAI211_X1 g195(.A(KEYINPUT91), .B(new_n370), .C1(new_n372), .C2(KEYINPUT13), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n375), .B(new_n377), .C1(new_n383), .C2(new_n374), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n373), .B(new_n374), .ZN(new_n385));
  INV_X1    g199(.A(G116), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT14), .A3(G122), .ZN(new_n387));
  INV_X1    g201(.A(new_n376), .ZN(new_n388));
  OAI211_X1 g202(.A(G107), .B(new_n387), .C1(new_n388), .C2(KEYINPUT14), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n385), .B(new_n389), .C1(G107), .C2(new_n388), .ZN(new_n390));
  XOR2_X1   g204(.A(KEYINPUT74), .B(G217), .Z(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n392), .A2(new_n188), .A3(G953), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n384), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n384), .B2(new_n390), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n294), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT15), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G478), .ZN(new_n398));
  INV_X1    g212(.A(G478), .ZN(new_n399));
  OAI221_X1 g213(.A(new_n294), .B1(KEYINPUT15), .B2(new_n399), .C1(new_n394), .C2(new_n395), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n398), .A2(KEYINPUT92), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT92), .B1(new_n398), .B2(new_n400), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n364), .A2(new_n369), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(G234), .A2(G237), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(G952), .A3(new_n308), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT93), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(KEYINPUT21), .B(G898), .Z(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n405), .A2(G902), .A3(G953), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n408), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G214), .B1(G237), .B2(G902), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(KEYINPUT68), .A2(G119), .ZN(new_n418));
  NOR2_X1   g232(.A1(KEYINPUT68), .A2(G119), .ZN(new_n419));
  OAI21_X1  g233(.A(G116), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n386), .A2(G119), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(KEYINPUT5), .A3(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n422), .B(G113), .C1(KEYINPUT5), .C2(new_n420), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT2), .B(G113), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n420), .A3(new_n421), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(new_n225), .ZN(new_n428));
  XOR2_X1   g242(.A(G110), .B(G122), .Z(new_n429));
  XOR2_X1   g243(.A(new_n429), .B(KEYINPUT8), .Z(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  MUX2_X1   g245(.A(new_n268), .B(new_n233), .S(new_n319), .Z(new_n432));
  INV_X1    g246(.A(G224), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(G953), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT7), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n432), .A2(new_n436), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n431), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT83), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n431), .A2(new_n441), .A3(new_n437), .A4(new_n438), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n277), .A2(new_n426), .A3(new_n423), .ZN(new_n443));
  OR2_X1    g257(.A1(KEYINPUT68), .A2(G119), .ZN(new_n444));
  NAND2_X1  g258(.A1(KEYINPUT68), .A2(G119), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n386), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n421), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n424), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n426), .A3(KEYINPUT69), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT69), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n450), .B(new_n424), .C1(new_n446), .C2(new_n447), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n449), .A2(new_n451), .A3(new_n270), .A4(new_n261), .ZN(new_n452));
  INV_X1    g266(.A(new_n429), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n443), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n440), .A2(new_n442), .A3(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(new_n432), .B(new_n434), .Z(new_n456));
  AOI21_X1  g270(.A(new_n427), .B1(new_n275), .B2(new_n276), .ZN(new_n457));
  INV_X1    g271(.A(new_n452), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n429), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n459), .A2(new_n454), .A3(KEYINPUT82), .A4(KEYINPUT6), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n459), .A2(new_n454), .A3(KEYINPUT6), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT82), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n453), .B1(new_n443), .B2(new_n452), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n456), .B(new_n460), .C1(new_n461), .C2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n455), .A2(new_n294), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G210), .B1(G237), .B2(G902), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT84), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n469), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n455), .A2(new_n466), .A3(new_n294), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n417), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n304), .A2(new_n404), .A3(new_n473), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n246), .A2(new_n251), .B1(new_n266), .B2(new_n267), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n449), .A2(new_n451), .ZN(new_n477));
  AOI21_X1  g291(.A(G134), .B1(new_n239), .B2(new_n241), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n374), .A2(new_n238), .ZN(new_n479));
  OAI21_X1  g293(.A(G131), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n235), .B1(new_n242), .B2(new_n245), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT70), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n233), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT70), .B1(new_n480), .B2(new_n481), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n476), .B(new_n477), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n486));
  NAND2_X1  g300(.A1(new_n312), .A2(G210), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT26), .B(G101), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n480), .A2(new_n481), .B1(new_n232), .B2(new_n205), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n491), .A2(new_n475), .A3(KEYINPUT30), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n476), .B1(new_n483), .B2(new_n484), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n492), .B1(KEYINPUT30), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n485), .B(new_n490), .C1(new_n494), .C2(new_n477), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT31), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n485), .A2(KEYINPUT28), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n480), .A2(new_n481), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT70), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n233), .A3(new_n482), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT28), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n501), .A2(new_n502), .A3(new_n476), .A4(new_n477), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n477), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n475), .B2(new_n491), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n490), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n501), .B2(new_n476), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n505), .B1(new_n511), .B2(new_n492), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT31), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n512), .A2(new_n513), .A3(new_n485), .A4(new_n490), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n496), .A2(new_n509), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT32), .ZN(new_n516));
  NOR2_X1   g330(.A1(G472), .A2(G902), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n516), .B1(new_n515), .B2(new_n517), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G472), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n512), .A2(new_n485), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT72), .B1(new_n522), .B2(new_n490), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n512), .A2(new_n485), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT72), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n508), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n504), .A2(new_n506), .A3(new_n490), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT29), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n523), .A2(new_n526), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n477), .B1(new_n501), .B2(new_n476), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n532), .B1(new_n497), .B2(new_n503), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n508), .A2(new_n528), .ZN(new_n534));
  AOI21_X1  g348(.A(G902), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n521), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT73), .B1(new_n520), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n515), .A2(new_n517), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT32), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT73), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n525), .B1(new_n524), .B2(new_n508), .ZN(new_n543));
  AOI211_X1 g357(.A(KEYINPUT72), .B(new_n490), .C1(new_n512), .C2(new_n485), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n543), .A2(new_n544), .A3(new_n529), .ZN(new_n545));
  INV_X1    g359(.A(new_n535), .ZN(new_n546));
  OAI21_X1  g360(.A(G472), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n541), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n537), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n321), .A2(new_n200), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n444), .A2(new_n445), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G128), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n206), .A2(KEYINPUT23), .A3(G119), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n551), .A2(G128), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n552), .B(new_n553), .C1(new_n554), .C2(KEYINPUT23), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(G110), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT24), .B(G110), .Z(new_n557));
  INV_X1    g371(.A(KEYINPUT75), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n552), .A2(new_n558), .B1(G119), .B2(new_n206), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n551), .A2(KEYINPUT75), .A3(G128), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n342), .B(new_n550), .C1(new_n556), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n555), .A2(G110), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n559), .A2(new_n557), .A3(new_n560), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n323), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT76), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n562), .A2(KEYINPUT76), .A3(new_n565), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n308), .A2(G221), .A3(G234), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT22), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(G137), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n568), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n566), .A2(new_n567), .A3(new_n572), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT25), .B1(new_n577), .B2(G902), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n392), .B1(G234), .B2(new_n294), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT25), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n576), .A2(new_n580), .A3(new_n294), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n579), .A2(G902), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n474), .A2(new_n549), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G101), .ZN(G3));
  NAND2_X1  g402(.A1(new_n515), .A2(new_n294), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G472), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n590), .A2(new_n538), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n304), .A2(new_n591), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n394), .A2(new_n395), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n593), .A2(KEYINPUT33), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(KEYINPUT33), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(G478), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n593), .A2(new_n399), .A3(new_n294), .ZN(new_n597));
  NAND2_X1  g411(.A1(G478), .A2(G902), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n364), .B2(new_n369), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n467), .A2(new_n468), .ZN(new_n602));
  INV_X1    g416(.A(new_n468), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n455), .A2(new_n466), .A3(new_n294), .A4(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n601), .A2(new_n417), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n592), .A2(new_n606), .A3(new_n586), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT34), .B(G104), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G6));
  NAND2_X1  g423(.A1(new_n363), .A2(KEYINPUT20), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n355), .B(new_n357), .C1(new_n361), .C2(new_n362), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n368), .ZN(new_n613));
  INV_X1    g427(.A(new_n403), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n613), .A2(new_n413), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n602), .A2(new_n414), .A3(new_n604), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n592), .A2(new_n615), .A3(new_n586), .A4(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT35), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n213), .ZN(G9));
  AND2_X1   g434(.A1(new_n304), .A2(new_n404), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n573), .A2(KEYINPUT36), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n566), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n583), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n582), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n621), .A2(new_n473), .A3(new_n591), .A4(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT37), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G110), .ZN(G12));
  INV_X1    g442(.A(G900), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n408), .B1(new_n629), .B2(new_n412), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n613), .A2(new_n614), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n582), .A2(new_n624), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n616), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n549), .A2(new_n304), .A3(new_n631), .A4(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G128), .ZN(G30));
  INV_X1    g449(.A(new_n485), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n508), .B1(new_n636), .B2(new_n532), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n637), .A2(KEYINPUT95), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n495), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(KEYINPUT95), .B2(new_n637), .ZN(new_n640));
  OAI21_X1  g454(.A(G472), .B1(new_n640), .B2(G902), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n625), .B1(new_n541), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n296), .A2(new_n303), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n189), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n630), .B(KEYINPUT96), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT39), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n414), .B(new_n642), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT38), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT94), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n470), .A2(new_n651), .A3(new_n472), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n651), .B1(new_n470), .B2(new_n472), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n654), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(KEYINPUT38), .A3(new_n652), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n649), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n364), .A2(new_n369), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n614), .ZN(new_n661));
  INV_X1    g475(.A(new_n647), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n659), .B(new_n661), .C1(KEYINPUT40), .C2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT97), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n202), .ZN(G45));
  INV_X1    g479(.A(new_n630), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n600), .B(new_n666), .C1(new_n364), .C2(new_n369), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n549), .A2(new_n304), .A3(new_n633), .A4(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT98), .B(G146), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G48));
  AOI21_X1  g485(.A(new_n585), .B1(new_n537), .B2(new_n548), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n299), .A2(new_n294), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G469), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n189), .A3(new_n303), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n672), .A2(new_n606), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT99), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT41), .B(G113), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G15));
  NOR2_X1   g494(.A1(new_n616), .A2(new_n675), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n549), .A2(new_n586), .A3(new_n615), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  NAND2_X1  g497(.A1(new_n660), .A2(new_n614), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n537), .B2(new_n548), .ZN(new_n685));
  INV_X1    g499(.A(new_n413), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n685), .A2(new_n686), .A3(new_n625), .A4(new_n681), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G119), .ZN(G21));
  OAI211_X1 g502(.A(new_n496), .B(new_n514), .C1(new_n490), .C2(new_n533), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n517), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n590), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n585), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n605), .A2(new_n417), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n692), .A2(new_n661), .A3(new_n693), .A4(new_n676), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G122), .ZN(G24));
  NOR2_X1   g509(.A1(new_n632), .A2(new_n691), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n668), .A3(new_n681), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G125), .ZN(G27));
  NAND3_X1  g512(.A1(new_n470), .A2(new_n472), .A3(new_n414), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n290), .A2(G469), .A3(new_n292), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n701), .A2(KEYINPUT100), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(KEYINPUT100), .ZN(new_n703));
  NAND2_X1  g517(.A1(G469), .A2(G902), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n702), .A2(new_n303), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n705), .A2(new_n189), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n672), .A2(new_n668), .A3(new_n700), .A4(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n518), .B2(new_n519), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n539), .A2(KEYINPUT101), .A3(new_n540), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n547), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(KEYINPUT42), .A3(new_n586), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n668), .A2(new_n700), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI22_X1  g529(.A1(new_n707), .A2(new_n708), .B1(new_n715), .B2(new_n706), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n235), .ZN(G33));
  NAND4_X1  g531(.A1(new_n672), .A2(new_n631), .A3(new_n700), .A4(new_n706), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G134), .ZN(G36));
  NAND2_X1  g533(.A1(new_n610), .A2(new_n358), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n720), .A2(new_n368), .A3(new_n600), .A4(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n364), .A2(new_n369), .A3(new_n599), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(KEYINPUT102), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n723), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n591), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n728), .A3(new_n625), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT104), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n290), .A2(KEYINPUT45), .A3(new_n292), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n286), .A2(new_n293), .ZN(new_n734));
  OAI211_X1 g548(.A(G469), .B(new_n733), .C1(new_n734), .C2(KEYINPUT45), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n735), .A2(new_n704), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n303), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n189), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n646), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n729), .A2(new_n730), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n699), .B(KEYINPUT103), .Z(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n732), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G137), .ZN(G39));
  NAND3_X1  g561(.A1(new_n739), .A2(KEYINPUT47), .A3(new_n189), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT47), .B1(new_n739), .B2(new_n189), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n537), .A2(new_n548), .A3(new_n585), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n751), .A2(new_n714), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n752), .A2(KEYINPUT105), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(KEYINPUT105), .ZN(new_n754));
  OAI22_X1  g568(.A1(new_n749), .A2(new_n750), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G140), .ZN(G42));
  NAND2_X1  g570(.A1(new_n674), .A2(new_n303), .ZN(new_n757));
  NOR2_X1   g571(.A1(KEYINPUT106), .A2(KEYINPUT49), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n415), .B1(KEYINPUT106), .B2(KEYINPUT49), .ZN(new_n760));
  AND4_X1   g574(.A1(new_n586), .A2(new_n759), .A3(new_n189), .A4(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n641), .A2(new_n541), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n658), .A4(new_n724), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n308), .A2(G952), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n414), .B1(new_n655), .B2(new_n657), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n692), .A2(new_n676), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n727), .A2(KEYINPUT111), .A3(new_n408), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT111), .B1(new_n727), .B2(new_n408), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n766), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n765), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n727), .A2(new_n408), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n727), .A2(KEYINPUT111), .A3(new_n408), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n767), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n774), .B1(new_n779), .B2(new_n766), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n773), .B1(new_n780), .B2(new_n772), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n771), .A2(KEYINPUT114), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(KEYINPUT115), .A3(new_n765), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n699), .A2(new_n675), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n762), .A2(new_n784), .A3(new_n586), .A4(new_n408), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n785), .A2(new_n369), .A3(new_n364), .A4(new_n600), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n696), .B(new_n784), .C1(new_n769), .C2(new_n770), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT116), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n777), .A2(new_n778), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(new_n790), .A3(new_n696), .A4(new_n784), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n786), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  AND4_X1   g606(.A1(KEYINPUT51), .A2(new_n781), .A3(new_n783), .A4(new_n792), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n789), .A2(new_n692), .A3(new_n743), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n749), .A2(new_n750), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n757), .B(KEYINPUT112), .Z(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n190), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n794), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n764), .B1(new_n793), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n712), .A2(new_n586), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n789), .A2(new_n801), .A3(new_n784), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT48), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n779), .A2(new_n617), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT117), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n797), .B(KEYINPUT113), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n794), .B1(new_n795), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n807), .A2(new_n783), .A3(new_n781), .A4(new_n792), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n800), .A2(new_n803), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n668), .A2(new_n706), .A3(new_n590), .A4(new_n690), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n520), .A2(new_n536), .A3(KEYINPUT73), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n542), .B1(new_n541), .B2(new_n547), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n304), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n398), .A2(new_n400), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT107), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n612), .A2(new_n368), .A3(new_n666), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT108), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n369), .B1(new_n610), .B2(new_n611), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT108), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n821), .A2(new_n822), .A3(new_n666), .A4(new_n818), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n812), .B1(new_n815), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n625), .A3(new_n700), .ZN(new_n826));
  INV_X1    g640(.A(new_n818), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n720), .A2(new_n827), .A3(new_n368), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n601), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n592), .A2(new_n586), .A3(new_n473), .A4(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n587), .A2(new_n626), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n826), .A2(new_n718), .A3(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n660), .A2(new_n616), .A3(new_n614), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n642), .A3(new_n666), .A4(new_n706), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n634), .A2(new_n669), .A3(new_n697), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n644), .B1(new_n537), .B2(new_n548), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n838), .B(new_n633), .C1(new_n631), .C2(new_n668), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(KEYINPUT52), .A3(new_n697), .A4(new_n834), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n832), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n687), .A2(new_n677), .A3(new_n682), .A4(new_n694), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n716), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n842), .B1(new_n844), .B2(KEYINPUT110), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT110), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n716), .B2(new_n843), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n841), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n826), .A2(new_n718), .A3(new_n831), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n837), .A2(new_n840), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n851), .A3(new_n844), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n842), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n848), .A2(new_n849), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT53), .A4(new_n844), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n854), .A2(KEYINPUT109), .B1(new_n856), .B2(KEYINPUT54), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n785), .A2(new_n601), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n856), .A2(KEYINPUT109), .A3(KEYINPUT54), .ZN(new_n859));
  NOR4_X1   g673(.A1(new_n811), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(G952), .A2(G953), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n763), .B1(new_n860), .B2(new_n861), .ZN(G75));
  NAND2_X1  g676(.A1(new_n848), .A2(new_n853), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(G210), .A3(G902), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n460), .B1(new_n461), .B2(new_n465), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(new_n456), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT55), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n868), .B1(new_n864), .B2(new_n865), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n308), .A2(G952), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT118), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(G51));
  XOR2_X1   g687(.A(new_n704), .B(KEYINPUT57), .Z(new_n874));
  AND3_X1   g688(.A1(new_n848), .A2(new_n849), .A3(new_n853), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n849), .B1(new_n848), .B2(new_n853), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(KEYINPUT119), .B(new_n874), .C1(new_n875), .C2(new_n876), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n299), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n863), .ZN(new_n882));
  OR3_X1    g696(.A1(new_n882), .A2(new_n294), .A3(new_n735), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n871), .B1(new_n881), .B2(new_n883), .ZN(G54));
  NOR2_X1   g698(.A1(new_n882), .A2(new_n294), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n361), .A2(new_n362), .ZN(new_n886));
  NAND2_X1  g700(.A1(KEYINPUT58), .A2(G475), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT120), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n886), .B1(new_n885), .B2(new_n888), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n889), .A2(new_n890), .A3(new_n871), .ZN(G60));
  XOR2_X1   g705(.A(new_n598), .B(KEYINPUT59), .Z(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n594), .A2(new_n595), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT121), .Z(new_n895));
  OAI211_X1 g709(.A(new_n893), .B(new_n895), .C1(new_n875), .C2(new_n876), .ZN(new_n896));
  INV_X1    g710(.A(new_n872), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n893), .B1(new_n857), .B2(new_n859), .ZN(new_n901));
  INV_X1    g715(.A(new_n895), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n896), .A2(KEYINPUT122), .A3(new_n897), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n900), .A2(new_n903), .A3(new_n904), .ZN(G63));
  NAND2_X1  g719(.A1(G217), .A2(G902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT60), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n848), .B2(new_n853), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n908), .A2(new_n623), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n897), .B1(new_n908), .B2(new_n576), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n912));
  OR2_X1    g726(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(KEYINPUT123), .B(KEYINPUT61), .C1(new_n909), .C2(new_n910), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(G66));
  INV_X1    g730(.A(new_n831), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(new_n843), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n308), .ZN(new_n919));
  OAI21_X1  g733(.A(G953), .B1(new_n410), .B2(new_n433), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n866), .B1(G898), .B2(new_n308), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(G69));
  INV_X1    g737(.A(new_n716), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n746), .A2(new_n755), .A3(new_n924), .A4(new_n718), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n839), .A2(new_n697), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n741), .A2(new_n801), .A3(new_n833), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n308), .B1(new_n925), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n629), .A2(G953), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(KEYINPUT125), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n931), .A2(new_n935), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n494), .B(new_n344), .Z(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  OAI221_X1 g754(.A(G953), .B1(new_n193), .B2(new_n629), .C1(new_n938), .C2(KEYINPUT126), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n928), .A2(new_n663), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n746), .A2(new_n755), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n672), .A2(new_n647), .A3(new_n700), .A4(new_n829), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n308), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n938), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n940), .A2(new_n941), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n941), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n938), .B1(new_n934), .B2(new_n936), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n939), .B1(new_n947), .B2(new_n308), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n950), .A2(new_n954), .ZN(G72));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT63), .Z(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n947), .B2(new_n918), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n958), .A2(new_n490), .A3(new_n524), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n523), .A2(new_n495), .A3(new_n526), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n957), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n961), .A2(KEYINPUT127), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n853), .B2(new_n855), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(KEYINPUT127), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n871), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n925), .A2(new_n918), .A3(new_n930), .ZN(new_n966));
  INV_X1    g780(.A(new_n957), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n508), .B(new_n522), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n959), .A2(new_n965), .A3(new_n968), .ZN(G57));
endmodule


