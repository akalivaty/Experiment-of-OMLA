//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901;
  XOR2_X1   g000(.A(KEYINPUT2), .B(G113), .Z(new_n187));
  XNOR2_X1  g001(.A(G116), .B(G119), .ZN(new_n188));
  OR2_X1    g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n187), .A2(new_n188), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT64), .B1(new_n192), .B2(G137), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n195));
  OAI211_X1 g009(.A(KEYINPUT64), .B(new_n195), .C1(new_n192), .C2(G137), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G131), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n194), .A2(new_n200), .A3(new_n196), .A4(new_n197), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(KEYINPUT65), .A3(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(G143), .B(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT0), .A3(G128), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT0), .B(G128), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n198), .A2(new_n208), .A3(G131), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n202), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n215), .A2(KEYINPUT1), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n216), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n213), .A2(KEYINPUT1), .A3(G146), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT66), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(G128), .B1(new_n212), .B2(new_n214), .ZN(new_n222));
  INV_X1    g036(.A(new_n220), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  NOR3_X1   g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n218), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n197), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n192), .A2(G137), .ZN(new_n228));
  OAI21_X1  g042(.A(G131), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n201), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT30), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n210), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(new_n210), .B2(new_n231), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n191), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n210), .A2(new_n231), .A3(new_n189), .A4(new_n190), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g051(.A(KEYINPUT67), .B(G237), .Z(new_n238));
  INV_X1    g052(.A(G953), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(G210), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n240), .B(KEYINPUT27), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(G101), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n241), .B(new_n242), .ZN(new_n243));
  OR2_X1    g057(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT29), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT28), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n210), .A2(new_n231), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n191), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n246), .B1(new_n248), .B2(new_n236), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n236), .A2(new_n246), .ZN(new_n250));
  INV_X1    g064(.A(new_n243), .ZN(new_n251));
  OR3_X1    g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n244), .A2(new_n245), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G902), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n253), .B(new_n254), .C1(new_n245), .C2(new_n252), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G472), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n235), .A2(new_n243), .A3(new_n236), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT31), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n235), .A2(KEYINPUT31), .A3(new_n243), .A4(new_n236), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n251), .B1(new_n249), .B2(new_n250), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT68), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n265), .B(new_n251), .C1(new_n249), .C2(new_n250), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT69), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(G472), .A2(G902), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n260), .A2(new_n261), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n270), .A2(new_n271), .A3(new_n264), .A4(new_n266), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n268), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT32), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n268), .A2(KEYINPUT32), .A3(new_n269), .A4(new_n272), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(KEYINPUT70), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n273), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT32), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n257), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n239), .A2(G221), .A3(G234), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n282), .B(KEYINPUT74), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT22), .B(G137), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(G125), .B(G140), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT73), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n211), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(KEYINPUT16), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT16), .ZN(new_n290));
  INV_X1    g104(.A(G140), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n291), .A3(G125), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n289), .A2(G146), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n216), .A2(KEYINPUT23), .A3(G119), .ZN(new_n294));
  INV_X1    g108(.A(G119), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G128), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(G128), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n294), .B(new_n296), .C1(new_n297), .C2(KEYINPUT23), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT72), .B(G110), .Z(new_n299));
  XOR2_X1   g113(.A(KEYINPUT24), .B(G110), .Z(new_n300));
  XNOR2_X1  g114(.A(G119), .B(G128), .ZN(new_n301));
  OAI22_X1  g115(.A1(new_n298), .A2(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n288), .A2(new_n293), .A3(new_n302), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n298), .A2(G110), .B1(new_n300), .B2(new_n301), .ZN(new_n304));
  INV_X1    g118(.A(new_n293), .ZN(new_n305));
  AOI21_X1  g119(.A(G146), .B1(new_n289), .B2(new_n292), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(KEYINPUT75), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n310), .B1(new_n303), .B2(new_n307), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n285), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n285), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n313), .B1(new_n308), .B2(KEYINPUT75), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n254), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n312), .A2(new_n314), .A3(new_n254), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n316), .ZN(new_n320));
  NAND2_X1  g134(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G217), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n323), .B1(G234), .B2(new_n254), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT71), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n324), .A2(G902), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n315), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n322), .A2(new_n325), .B1(new_n315), .B2(new_n327), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT77), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n220), .B1(new_n203), .B2(G128), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n224), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n219), .A2(KEYINPUT66), .A3(new_n220), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n217), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT10), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G104), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT3), .B1(new_n341), .B2(G107), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n343));
  INV_X1    g157(.A(G107), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(G104), .ZN(new_n345));
  INV_X1    g159(.A(G101), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n341), .A2(G107), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n342), .A2(new_n345), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n341), .A2(G107), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n344), .A2(G104), .ZN(new_n350));
  OAI21_X1  g164(.A(G101), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT79), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n352), .B1(new_n217), .B2(new_n335), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n340), .A2(new_n353), .B1(new_n354), .B2(new_n339), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n202), .A2(new_n209), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n342), .A2(new_n345), .A3(new_n347), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G101), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(KEYINPUT4), .A3(new_n348), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n360), .A3(G101), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n207), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n207), .A2(KEYINPUT78), .A3(new_n359), .A4(new_n361), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n355), .A2(new_n356), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G110), .B(G140), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n239), .A2(G227), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT80), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT79), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n352), .B(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n338), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n356), .B1(new_n375), .B2(new_n354), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n372), .B1(new_n376), .B2(KEYINPUT12), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n354), .B1(new_n353), .B2(new_n226), .ZN(new_n378));
  INV_X1    g192(.A(new_n356), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n378), .A2(new_n372), .A3(KEYINPUT12), .A4(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(KEYINPUT12), .B2(new_n376), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n371), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n356), .B1(new_n355), .B2(new_n366), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n370), .B1(new_n367), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT82), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT82), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n386), .B(new_n370), .C1(new_n367), .C2(new_n383), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n382), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G469), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(new_n254), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n383), .B1(new_n371), .B2(KEYINPUT81), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n367), .B2(new_n370), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n381), .A2(new_n377), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n370), .B1(new_n395), .B2(new_n367), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n396), .A3(G469), .ZN(new_n397));
  NAND2_X1  g211(.A1(G469), .A2(G902), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n390), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT9), .B(G234), .ZN(new_n400));
  OAI21_X1  g214(.A(G221), .B1(new_n400), .B2(G902), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G113), .B(G122), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(new_n341), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n238), .A2(G214), .A3(new_n239), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT87), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n238), .A2(new_n408), .A3(G214), .A4(new_n239), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n406), .A2(new_n407), .A3(new_n213), .A4(new_n409), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n405), .A2(new_n213), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(G143), .B1(new_n405), .B2(KEYINPUT87), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n407), .B1(new_n413), .B2(new_n409), .ZN(new_n414));
  OAI21_X1  g228(.A(G131), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n409), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT88), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n417), .A2(new_n200), .A3(new_n410), .A4(new_n411), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT17), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n415), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n305), .A2(new_n306), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT89), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n420), .B(new_n422), .C1(new_n419), .C2(new_n415), .ZN(new_n423));
  OAI211_X1 g237(.A(KEYINPUT18), .B(G131), .C1(new_n412), .C2(new_n414), .ZN(new_n424));
  NAND2_X1  g238(.A1(KEYINPUT18), .A2(G131), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n417), .A2(new_n410), .A3(new_n411), .A4(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n288), .B1(new_n211), .B2(new_n286), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n404), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n415), .A2(new_n418), .A3(new_n419), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n422), .B1(new_n415), .B2(new_n419), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n404), .B(new_n428), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n254), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G475), .ZN(new_n435));
  INV_X1    g249(.A(new_n428), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n287), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n437), .B2(new_n286), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n293), .B1(new_n439), .B2(G146), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n415), .B2(new_n418), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n432), .B1(new_n442), .B2(new_n404), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n444));
  NOR2_X1   g258(.A1(G475), .A2(G902), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n444), .B1(new_n443), .B2(new_n445), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n435), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G128), .B(G143), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(new_n192), .ZN(new_n451));
  INV_X1    g265(.A(G116), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT14), .A3(G122), .ZN(new_n453));
  XOR2_X1   g267(.A(G116), .B(G122), .Z(new_n454));
  OAI211_X1 g268(.A(G107), .B(new_n453), .C1(new_n454), .C2(KEYINPUT14), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n451), .B(new_n455), .C1(G107), .C2(new_n454), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n454), .B(G107), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n450), .A2(KEYINPUT13), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n213), .A2(G128), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n458), .B(G134), .C1(KEYINPUT13), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n450), .A2(new_n192), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT90), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n456), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n400), .A2(new_n323), .A3(G953), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n464), .A2(new_n466), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n254), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT15), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(G478), .ZN(new_n471));
  INV_X1    g285(.A(G478), .ZN(new_n472));
  OAI221_X1 g286(.A(new_n254), .B1(KEYINPUT15), .B2(new_n472), .C1(new_n467), .C2(new_n468), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT91), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n471), .A2(KEYINPUT91), .A3(new_n473), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G952), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n479), .A2(KEYINPUT92), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(KEYINPUT92), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n239), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(G234), .B2(G237), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  XOR2_X1   g298(.A(KEYINPUT21), .B(G898), .Z(new_n485));
  AOI211_X1 g299(.A(new_n254), .B(new_n239), .C1(G234), .C2(G237), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n484), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n478), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n449), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G214), .B1(G237), .B2(G902), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G210), .B1(G237), .B2(G902), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n207), .A2(G125), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n495), .B1(new_n338), .B2(G125), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n239), .A2(G224), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT86), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n496), .B(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n295), .A2(G116), .ZN(new_n500));
  OAI21_X1  g314(.A(G113), .B1(new_n500), .B2(KEYINPUT5), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(KEYINPUT5), .B2(new_n188), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(new_n188), .B2(new_n187), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n353), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT84), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n191), .A2(new_n359), .A3(new_n361), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT83), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n353), .A2(new_n503), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT84), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(G110), .B(G122), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n505), .A2(new_n507), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n505), .A2(new_n507), .A3(new_n510), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n511), .B(KEYINPUT85), .Z(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(KEYINPUT6), .A3(new_n515), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n499), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT7), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n498), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n496), .B(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n508), .B1(new_n503), .B2(new_n352), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n511), .B(KEYINPUT8), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(G902), .B1(new_n525), .B2(new_n512), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n494), .B1(new_n519), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n499), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n512), .A2(KEYINPUT6), .B1(new_n514), .B2(new_n515), .ZN(new_n530));
  INV_X1    g344(.A(new_n518), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n493), .A3(new_n526), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n492), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n402), .A2(new_n490), .A3(new_n534), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n281), .A2(new_n334), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(new_n346), .ZN(G3));
  NAND3_X1  g351(.A1(new_n268), .A2(new_n254), .A3(new_n272), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G472), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n273), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n399), .A2(new_n401), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n540), .A2(new_n334), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n534), .A2(new_n488), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n467), .A2(new_n468), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(KEYINPUT33), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G478), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n469), .A2(G478), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n472), .A2(new_n254), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n449), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n543), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n542), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g368(.A(KEYINPUT34), .B(G104), .Z(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(G6));
  NAND2_X1  g370(.A1(new_n443), .A2(new_n445), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT20), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT93), .A3(new_n446), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n478), .B1(G475), .B2(new_n434), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT93), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n448), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(new_n543), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n542), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT35), .B(G107), .Z(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(G9));
  INV_X1    g382(.A(new_n535), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n313), .A2(KEYINPUT36), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(new_n308), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n327), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n326), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(new_n540), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT37), .B(G110), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(G12));
  INV_X1    g391(.A(G900), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n483), .B1(new_n578), .B2(new_n486), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n559), .A2(new_n560), .A3(new_n562), .A4(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(KEYINPUT94), .A3(new_n534), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n584));
  INV_X1    g398(.A(new_n534), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n584), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n277), .A2(new_n280), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n256), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n587), .A2(new_n589), .A3(new_n402), .A4(new_n573), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT95), .B(G128), .Z(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G30));
  XOR2_X1   g406(.A(new_n579), .B(KEYINPUT39), .Z(new_n593));
  NAND2_X1  g407(.A1(new_n402), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n594), .A2(KEYINPUT40), .ZN(new_n595));
  INV_X1    g409(.A(new_n478), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n449), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n528), .A2(new_n533), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n573), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n491), .ZN(new_n602));
  NOR4_X1   g416(.A1(new_n595), .A2(new_n597), .A3(new_n600), .A4(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n237), .A2(new_n251), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n248), .A2(new_n236), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n254), .B1(new_n606), .B2(new_n243), .ZN(new_n607));
  OAI21_X1  g421(.A(G472), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n588), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n603), .B(new_n609), .C1(KEYINPUT40), .C2(new_n594), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT97), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G143), .ZN(G45));
  AOI22_X1  g426(.A1(new_n558), .A2(new_n446), .B1(new_n434), .B2(G475), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(new_n550), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n580), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n615), .A2(new_n585), .A3(new_n541), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n589), .A2(new_n616), .A3(new_n573), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G146), .ZN(G48));
  INV_X1    g432(.A(new_n334), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n388), .A2(new_n254), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G469), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n621), .A2(new_n390), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n401), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n589), .A2(new_n619), .A3(new_n553), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT41), .B(G113), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G15));
  NAND4_X1  g441(.A1(new_n589), .A2(new_n619), .A3(new_n565), .A4(new_n624), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G116), .ZN(G18));
  AND4_X1   g443(.A1(new_n534), .A2(new_n401), .A3(new_n390), .A4(new_n621), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n630), .A2(new_n490), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n589), .A2(new_n631), .A3(new_n573), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G119), .ZN(G21));
  NOR2_X1   g447(.A1(new_n623), .A2(new_n543), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT98), .B(G472), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n270), .A2(new_n263), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n538), .A2(new_n635), .B1(new_n269), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n637), .A2(new_n332), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n597), .A2(KEYINPUT99), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n449), .A2(new_n640), .A3(new_n596), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n634), .A2(new_n638), .A3(new_n639), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G122), .ZN(G24));
  AND2_X1   g457(.A1(new_n637), .A2(new_n573), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n552), .A2(new_n579), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n645), .A3(new_n630), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G125), .ZN(G27));
  NOR2_X1   g461(.A1(new_n598), .A2(new_n492), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n541), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n541), .A2(new_n649), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n645), .B(new_n648), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n275), .A2(new_n256), .A3(new_n276), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n332), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT42), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n648), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n402), .A2(KEYINPUT100), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n657), .B1(new_n658), .B2(new_n650), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n615), .A2(KEYINPUT42), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n589), .A2(new_n659), .A3(new_n660), .A4(new_n619), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(new_n200), .ZN(G33));
  AND4_X1   g477(.A1(new_n589), .A2(new_n659), .A3(new_n619), .A4(new_n582), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n192), .ZN(G36));
  AOI21_X1  g479(.A(KEYINPUT45), .B1(new_n394), .B2(new_n396), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n389), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n394), .A2(KEYINPUT45), .A3(new_n396), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n398), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n672), .B(KEYINPUT102), .Z(new_n673));
  OAI21_X1  g487(.A(new_n390), .B1(new_n670), .B2(new_n671), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT101), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n674), .A2(KEYINPUT101), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n677), .A2(new_n401), .A3(new_n593), .ZN(new_n678));
  AOI21_X1  g492(.A(KEYINPUT43), .B1(new_n613), .B2(new_n551), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT103), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n613), .A2(KEYINPUT104), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n613), .A2(KEYINPUT104), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n551), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n680), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n540), .A3(new_n573), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n657), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n678), .B(new_n688), .C1(new_n687), .C2(new_n686), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G137), .ZN(G39));
  NAND2_X1  g504(.A1(new_n677), .A2(new_n401), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n677), .A2(KEYINPUT47), .A3(new_n401), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n615), .A2(new_n619), .A3(new_n657), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n281), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G140), .ZN(G42));
  INV_X1    g512(.A(new_n622), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n699), .A2(KEYINPUT49), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(KEYINPUT49), .ZN(new_n701));
  INV_X1    g515(.A(new_n401), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n329), .A2(new_n492), .A3(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n700), .A2(new_n600), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  OR3_X1    g518(.A1(new_n704), .A2(new_n609), .A3(new_n684), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n625), .A2(new_n628), .A3(new_n632), .A4(new_n642), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n662), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n474), .B(KEYINPUT106), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n449), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n543), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n542), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n711), .B1(new_n574), .B2(new_n540), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n542), .A2(new_n553), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n713), .B1(new_n536), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n589), .A2(new_n619), .A3(new_n569), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(KEYINPUT105), .A3(new_n554), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n712), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n708), .A2(new_n580), .ZN(new_n719));
  AND4_X1   g533(.A1(new_n435), .A2(new_n719), .A3(new_n559), .A4(new_n562), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n589), .A2(new_n402), .A3(new_n573), .A4(new_n720), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n644), .B(new_n645), .C1(new_n651), .C2(new_n652), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n664), .B1(new_n723), .B2(new_n648), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n707), .A2(new_n718), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT107), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n707), .A2(new_n718), .A3(new_n724), .A4(new_n727), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n639), .A2(new_n641), .A3(new_n534), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n573), .A2(new_n579), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT108), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n609), .A2(new_n731), .A3(new_n402), .A4(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n590), .A2(new_n734), .A3(new_n617), .A4(new_n646), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n644), .A2(new_n645), .A3(new_n630), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n281), .A2(new_n601), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n738), .B1(new_n739), .B2(new_n616), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(KEYINPUT52), .A3(new_n590), .A4(new_n734), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n737), .A2(new_n741), .A3(KEYINPUT110), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT110), .B1(new_n737), .B2(new_n741), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n729), .A2(KEYINPUT53), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n737), .A2(new_n741), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n735), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n736), .B2(new_n752), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n729), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n748), .A2(new_n749), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n759), .A3(KEYINPUT54), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n726), .A2(new_n728), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n756), .B1(new_n761), .B2(new_n744), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n718), .A2(new_n724), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n707), .A2(KEYINPUT53), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n766), .B1(new_n763), .B2(new_n764), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(new_n754), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n769), .A2(KEYINPUT54), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n760), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n759), .B1(new_n758), .B2(KEYINPUT54), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n685), .A2(new_n483), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n775), .A2(new_n638), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n630), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n623), .A2(new_n657), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n619), .A3(new_n483), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n609), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n482), .B1(new_n780), .B2(new_n614), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n775), .A2(new_n778), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n783), .B(KEYINPUT118), .Z(new_n784));
  INV_X1    g598(.A(new_n655), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT48), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT48), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n784), .A2(new_n788), .A3(new_n785), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n782), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n784), .A2(new_n644), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n624), .A2(new_n492), .A3(new_n600), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT117), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n776), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n776), .A2(new_n648), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n695), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n622), .B(KEYINPUT116), .Z(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n702), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n797), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n780), .A2(new_n613), .A3(new_n550), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n791), .A2(new_n796), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n802), .B1(new_n800), .B2(KEYINPUT115), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n695), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n799), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n810), .A2(new_n791), .A3(new_n796), .A4(new_n805), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n790), .B(new_n806), .C1(new_n811), .C2(KEYINPUT51), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n771), .A2(new_n772), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(G952), .A2(G953), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n705), .B1(new_n813), .B2(new_n814), .ZN(G75));
  NOR2_X1   g629(.A1(new_n239), .A2(G952), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n254), .B1(new_n762), .B2(new_n768), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT56), .B1(new_n817), .B2(G210), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n816), .B1(new_n818), .B2(KEYINPUT119), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n530), .A2(new_n531), .A3(new_n529), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n519), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT55), .Z(new_n822));
  AOI211_X1 g636(.A(KEYINPUT119), .B(new_n822), .C1(new_n818), .C2(KEYINPUT120), .ZN(new_n823));
  INV_X1    g637(.A(new_n822), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n769), .A2(G210), .A3(G902), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT56), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(KEYINPUT120), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n824), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n819), .B1(new_n823), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT121), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n832), .B(new_n819), .C1(new_n823), .C2(new_n829), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(G51));
  NAND2_X1  g648(.A1(new_n769), .A2(KEYINPUT54), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n770), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n398), .B(KEYINPUT57), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n388), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n669), .B(KEYINPUT122), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n817), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n816), .B1(new_n838), .B2(new_n840), .ZN(G54));
  NAND2_X1  g655(.A1(KEYINPUT58), .A2(G475), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT123), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n817), .A2(new_n843), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n844), .A2(new_n443), .ZN(new_n845));
  INV_X1    g659(.A(new_n816), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n443), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT124), .ZN(G60));
  XNOR2_X1  g663(.A(new_n548), .B(KEYINPUT59), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n545), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n846), .B1(new_n836), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n850), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n771), .B2(new_n772), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n852), .B1(new_n854), .B2(new_n545), .ZN(G63));
  NAND2_X1  g669(.A1(G217), .A2(G902), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT60), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n762), .B2(new_n768), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n571), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT125), .Z(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n846), .B1(new_n858), .B2(new_n315), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(KEYINPUT61), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n865), .B1(new_n860), .B2(new_n862), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n864), .A2(new_n866), .ZN(G66));
  AOI21_X1  g681(.A(new_n239), .B1(new_n485), .B2(G224), .ZN(new_n868));
  INV_X1    g682(.A(new_n718), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n869), .A2(new_n706), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n868), .B1(new_n870), .B2(new_n239), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n517), .B(new_n518), .C1(G898), .C2(new_n239), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n871), .B(new_n872), .Z(G69));
  INV_X1    g687(.A(new_n662), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n697), .A2(new_n689), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n740), .A2(new_n590), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT126), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n730), .A2(new_n655), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n664), .B1(new_n678), .B2(new_n878), .ZN(new_n879));
  AND4_X1   g693(.A1(new_n874), .A2(new_n875), .A3(new_n877), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n239), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n233), .A2(new_n234), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(new_n439), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n881), .B(new_n883), .C1(new_n578), .C2(new_n239), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n611), .A2(new_n877), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT62), .Z(new_n886));
  AOI211_X1 g700(.A(new_n657), .B(new_n594), .C1(new_n552), .C2(new_n709), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n887), .A2(new_n589), .A3(new_n619), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n886), .A2(new_n888), .A3(new_n875), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(G953), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n884), .B1(new_n890), .B2(new_n883), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n239), .B1(G227), .B2(G900), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n891), .B(new_n892), .ZN(G72));
  AND2_X1   g707(.A1(new_n244), .A2(new_n258), .ZN(new_n894));
  NAND2_X1  g708(.A1(G472), .A2(G902), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT63), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n816), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n237), .A2(new_n251), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n889), .A2(new_n604), .B1(new_n880), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n897), .B1(new_n899), .B2(new_n870), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n894), .A2(new_n896), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n758), .B2(new_n901), .ZN(G57));
endmodule


