//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n204));
  XOR2_X1   g003(.A(G211gat), .B(G218gat), .Z(new_n205));
  INV_X1    g004(.A(KEYINPUT72), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  INV_X1    g007(.A(G211gat), .ZN(new_n209));
  INV_X1    g008(.A(G218gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n208), .B1(KEYINPUT22), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n207), .B(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n204), .B1(new_n213), .B2(KEYINPUT29), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT75), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT75), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G141gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT76), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n216), .A2(new_n218), .A3(new_n219), .A4(G148gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  INV_X1    g020(.A(G155gat), .ZN(new_n222));
  INV_X1    g021(.A(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n221), .B1(new_n224), .B2(KEYINPUT2), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT76), .B1(new_n215), .B2(G148gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT75), .B(G141gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(G148gat), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT77), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n216), .A2(new_n218), .A3(G148gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n227), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT77), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n233), .A2(new_n234), .A3(new_n220), .A4(new_n225), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G148gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G141gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n215), .A2(G148gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT74), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n238), .A2(new_n239), .B1(new_n240), .B2(KEYINPUT2), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n221), .A2(KEYINPUT74), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(G155gat), .A3(G162gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n243), .A3(new_n224), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n236), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n203), .B1(new_n214), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n245), .B1(new_n230), .B2(new_n235), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n204), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT29), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT86), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n213), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n252), .A2(KEYINPUT86), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n248), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT87), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT87), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n258), .B(new_n248), .C1(new_n254), .C2(new_n255), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT85), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n205), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n205), .A2(new_n261), .ZN(new_n263));
  OR3_X1    g062(.A1(new_n262), .A2(new_n263), .A3(new_n212), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT29), .B1(new_n263), .B2(new_n212), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n249), .B1(new_n204), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n267), .B1(new_n252), .B2(new_n213), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n268), .B1(G228gat), .B2(G233gat), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n260), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(KEYINPUT31), .B(G50gat), .Z(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n272), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n260), .A2(new_n270), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G78gat), .B(G106gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(G22gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT25), .ZN(new_n281));
  NOR2_X1   g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n282), .B1(KEYINPUT23), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G176gat), .ZN(new_n285));
  INV_X1    g084(.A(G169gat), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n286), .A2(KEYINPUT23), .ZN(new_n287));
  AOI211_X1 g086(.A(new_n281), .B(new_n284), .C1(new_n285), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT24), .B1(new_n289), .B2(KEYINPUT65), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(KEYINPUT65), .B2(new_n289), .ZN(new_n291));
  AND3_X1   g090(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n292));
  INV_X1    g091(.A(G183gat), .ZN(new_n293));
  INV_X1    g092(.A(G190gat), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n289), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n295), .B1(KEYINPUT24), .B2(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(KEYINPUT64), .B(G176gat), .Z(new_n300));
  AOI21_X1  g099(.A(new_n284), .B1(new_n300), .B2(new_n287), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n281), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT27), .B(G183gat), .Z(new_n305));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n305), .A2(new_n306), .A3(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(KEYINPUT66), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(new_n293), .B2(KEYINPUT27), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n294), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n307), .B1(new_n311), .B2(new_n306), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n286), .A2(new_n285), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT26), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(new_n314), .A3(new_n283), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n315), .B(new_n289), .C1(new_n314), .C2(new_n313), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT67), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n304), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n320));
  OAI21_X1  g119(.A(G120gat), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G113gat), .ZN(new_n322));
  INV_X1    g121(.A(G120gat), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT1), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G134gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G127gat), .ZN(new_n326));
  INV_X1    g125(.A(G127gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G134gat), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n321), .A2(new_n324), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n326), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n322), .A2(new_n323), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT1), .ZN(new_n333));
  NAND2_X1  g132(.A1(G113gat), .A2(G120gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n327), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT70), .ZN(new_n339));
  OR2_X1    g138(.A1(new_n318), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n318), .A2(new_n339), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G227gat), .A2(G233gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT34), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT34), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n340), .A2(new_n341), .A3(new_n346), .A4(new_n343), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G15gat), .B(G43gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(G71gat), .B(G99gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n342), .A2(new_n344), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT33), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n352), .A2(KEYINPUT32), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT33), .B1(new_n342), .B2(new_n344), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n345), .B(new_n347), .C1(new_n357), .C2(new_n351), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n356), .B1(new_n355), .B2(new_n358), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n273), .A2(new_n278), .A3(new_n275), .ZN(new_n362));
  AND4_X1   g161(.A1(new_n202), .A2(new_n280), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  AOI211_X1 g162(.A(new_n245), .B(new_n338), .C1(new_n230), .C2(new_n235), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n339), .A2(new_n247), .ZN(new_n367));
  XOR2_X1   g166(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(new_n338), .A3(new_n250), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n247), .A2(new_n338), .ZN(new_n374));
  INV_X1    g173(.A(new_n338), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n249), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n370), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n370), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n249), .A2(new_n375), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n382), .B2(new_n364), .ZN(new_n383));
  INV_X1    g182(.A(new_n379), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT80), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n373), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT81), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n373), .B(new_n388), .C1(new_n380), .C2(new_n385), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n367), .A2(new_n368), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT82), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n367), .A2(KEYINPUT82), .A3(new_n368), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n393), .B(new_n394), .C1(new_n365), .C2(new_n364), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n395), .A2(new_n370), .A3(new_n372), .A4(new_n379), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G1gat), .B(G29gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(KEYINPUT0), .ZN(new_n399));
  XNOR2_X1  g198(.A(G57gat), .B(G85gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n397), .A2(KEYINPUT6), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n390), .B2(new_n396), .ZN(new_n404));
  INV_X1    g203(.A(new_n389), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n378), .B1(new_n377), .B2(new_n379), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n383), .A2(KEYINPUT80), .A3(new_n384), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n388), .B1(new_n408), .B2(new_n373), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n396), .B(new_n401), .C1(new_n405), .C2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n403), .B1(new_n404), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n213), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n318), .A2(G226gat), .A3(G233gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n318), .A2(new_n251), .B1(G226gat), .B2(G233gat), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT73), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n417), .A2(KEYINPUT73), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n417), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n415), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(new_n213), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  NAND2_X1  g226(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n427), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n420), .B2(new_n423), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(KEYINPUT30), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT30), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n424), .A2(new_n432), .A3(new_n427), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n413), .A2(KEYINPUT88), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT88), .B1(new_n413), .B2(new_n434), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n363), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT89), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n363), .B(KEYINPUT89), .C1(new_n435), .C2(new_n436), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT84), .ZN(new_n442));
  INV_X1    g241(.A(new_n403), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n404), .B1(new_n412), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n410), .A2(KEYINPUT83), .A3(new_n411), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n434), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n442), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n410), .A2(KEYINPUT83), .A3(new_n411), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT83), .B1(new_n410), .B2(new_n411), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n450), .A2(new_n451), .A3(new_n404), .ZN(new_n452));
  OAI211_X1 g251(.A(KEYINPUT84), .B(new_n434), .C1(new_n452), .C2(new_n443), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n280), .A2(new_n362), .ZN(new_n454));
  INV_X1    g253(.A(new_n361), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n449), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT35), .ZN(new_n458));
  INV_X1    g257(.A(new_n454), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n449), .B2(new_n453), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT36), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n361), .A2(KEYINPUT71), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(KEYINPUT71), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n462), .A2(KEYINPUT71), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n464), .B(new_n465), .C1(new_n359), .C2(new_n360), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n427), .B1(new_n424), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT38), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n213), .B1(new_n418), .B2(new_n419), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT37), .B1(new_n422), .B2(new_n414), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n428), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n424), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT37), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n471), .B1(new_n477), .B2(new_n469), .ZN(new_n478));
  OR3_X1    g277(.A1(new_n475), .A2(new_n413), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n434), .A2(new_n404), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n370), .B1(new_n395), .B2(new_n372), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT39), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n402), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n374), .A2(new_n376), .A3(new_n370), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT39), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT40), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n454), .B1(new_n480), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n467), .B1(new_n479), .B2(new_n488), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n441), .A2(new_n458), .B1(new_n461), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT16), .ZN(new_n492));
  INV_X1    g291(.A(G1gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT94), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT94), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G1gat), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n492), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT95), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n491), .B1(new_n497), .B2(new_n498), .ZN(new_n500));
  OAI221_X1 g299(.A(KEYINPUT96), .B1(G1gat), .B2(new_n491), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(G8gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT97), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT15), .ZN(new_n504));
  INV_X1    g303(.A(G43gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(G50gat), .ZN(new_n506));
  INV_X1    g305(.A(G50gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(G43gat), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n504), .B1(new_n509), .B2(KEYINPUT92), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT92), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n506), .B2(new_n508), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G29gat), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n514), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT14), .B(G29gat), .ZN(new_n516));
  INV_X1    g315(.A(G36gat), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n507), .A2(G43gat), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n508), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(new_n521), .B2(new_n522), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n518), .B1(new_n524), .B2(new_n504), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n520), .B1(new_n513), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n503), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n512), .ZN(new_n530));
  MUX2_X1   g329(.A(new_n518), .B(new_n525), .S(new_n530), .Z(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n531), .A2(new_n532), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n534), .A2(new_n502), .A3(new_n535), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n527), .A2(new_n529), .A3(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n537), .A2(KEYINPUT18), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(KEYINPUT18), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n503), .B(new_n526), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n528), .B(KEYINPUT13), .Z(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT91), .ZN(new_n545));
  XOR2_X1   g344(.A(G169gat), .B(G197gat), .Z(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n549), .B(KEYINPUT12), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n550), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n538), .A2(new_n552), .A3(new_n539), .A4(new_n542), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT7), .ZN(new_n556));
  INV_X1    g355(.A(G85gat), .ZN(new_n557));
  OAI21_X1  g356(.A(G92gat), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G92gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n558), .A2(new_n560), .B1(new_n556), .B2(new_n557), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(new_n563), .B2(KEYINPUT103), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(KEYINPUT103), .B2(new_n563), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G99gat), .B(G106gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n526), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G232gat), .ZN(new_n570));
  INV_X1    g369(.A(G233gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n533), .A2(new_n568), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n574), .B1(new_n575), .B2(new_n535), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(G190gat), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n577), .A2(new_n210), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT102), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n210), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n582), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n578), .A2(new_n579), .A3(new_n584), .A4(new_n580), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G134gat), .B(G162gat), .Z(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n583), .A2(new_n585), .A3(new_n587), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT21), .ZN(new_n593));
  NAND2_X1  g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  OR3_X1    g394(.A1(new_n595), .A2(KEYINPUT100), .A3(KEYINPUT9), .ZN(new_n596));
  INV_X1    g395(.A(G64gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(KEYINPUT99), .A3(G57gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n596), .B(new_n598), .C1(new_n595), .C2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT100), .B1(new_n595), .B2(KEYINPUT9), .ZN(new_n601));
  XOR2_X1   g400(.A(G57gat), .B(G64gat), .Z(new_n602));
  OAI21_X1  g401(.A(new_n601), .B1(new_n602), .B2(KEYINPUT99), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n602), .A2(KEYINPUT9), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n599), .A2(KEYINPUT98), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(KEYINPUT98), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n594), .A3(new_n606), .ZN(new_n607));
  OAI22_X1  g406(.A1(new_n600), .A2(new_n603), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n503), .B1(new_n593), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n593), .ZN(new_n610));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n609), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT101), .ZN(new_n616));
  XOR2_X1   g415(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n614), .A2(new_n620), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n568), .A2(new_n608), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT105), .Z(new_n628));
  AOI21_X1  g427(.A(KEYINPUT104), .B1(new_n568), .B2(new_n608), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n625), .B(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n630), .A2(new_n626), .ZN(new_n631));
  INV_X1    g430(.A(G230gat), .ZN(new_n632));
  OAI22_X1  g431(.A1(new_n628), .A2(new_n631), .B1(new_n632), .B2(new_n571), .ZN(new_n633));
  OR3_X1    g432(.A1(new_n630), .A2(new_n632), .A3(new_n571), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n633), .A2(new_n634), .A3(new_n638), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n592), .A2(new_n624), .A3(new_n643), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n490), .A2(new_n555), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n447), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n448), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n648), .A2(G8gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT16), .B(G8gat), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT42), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(KEYINPUT42), .B2(new_n651), .ZN(G1325gat));
  INV_X1    g452(.A(new_n645), .ZN(new_n654));
  INV_X1    g453(.A(new_n467), .ZN(new_n655));
  OAI21_X1  g454(.A(G15gat), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n455), .A2(G15gat), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n656), .B1(new_n654), .B2(new_n657), .ZN(G1326gat));
  NAND2_X1  g457(.A1(new_n645), .A2(new_n454), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT43), .B(G22gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  INV_X1    g460(.A(KEYINPUT45), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n624), .A2(new_n555), .A3(new_n642), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OR3_X1    g463(.A1(new_n490), .A2(new_n592), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n447), .A2(new_n514), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n662), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n665), .A2(new_n662), .A3(new_n666), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n592), .A2(KEYINPUT44), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n489), .B1(new_n460), .B2(KEYINPUT106), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672));
  AOI211_X1 g471(.A(new_n672), .B(new_n459), .C1(new_n449), .C2(new_n453), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n439), .A2(new_n440), .B1(new_n457), .B2(KEYINPUT35), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n669), .B(new_n670), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT44), .B1(new_n490), .B2(new_n592), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n441), .A2(new_n458), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n679), .B1(new_n673), .B2(new_n671), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n669), .B1(new_n680), .B2(new_n670), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n664), .B1(new_n678), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(new_n447), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n667), .B(new_n668), .C1(new_n684), .C2(new_n514), .ZN(G1328gat));
  NAND2_X1  g484(.A1(new_n448), .A2(new_n517), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n665), .A2(KEYINPUT46), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT46), .B1(new_n665), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n683), .A2(new_n448), .ZN(new_n691));
  OAI211_X1 g490(.A(KEYINPUT108), .B(new_n690), .C1(new_n691), .C2(new_n517), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n517), .B1(new_n683), .B2(new_n448), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(new_n689), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n695), .ZN(G1329gat));
  NAND3_X1  g495(.A1(new_n683), .A2(G43gat), .A3(new_n467), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n505), .B1(new_n665), .B2(new_n455), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT47), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n697), .A2(new_n701), .A3(new_n698), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(G1330gat));
  NAND2_X1  g502(.A1(new_n676), .A2(new_n677), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n454), .B(new_n663), .C1(new_n704), .C2(new_n681), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT109), .B1(new_n705), .B2(G50gat), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n665), .A2(G50gat), .A3(new_n459), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n705), .B2(G50gat), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI221_X4 g509(.A(new_n707), .B1(KEYINPUT109), .B2(KEYINPUT48), .C1(new_n705), .C2(G50gat), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(G1331gat));
  NOR2_X1   g511(.A1(new_n674), .A2(new_n675), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n592), .A2(new_n555), .A3(new_n624), .A4(new_n642), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n447), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g516(.A(new_n434), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT110), .B(KEYINPUT111), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1333gat));
  XOR2_X1   g522(.A(new_n361), .B(KEYINPUT112), .Z(new_n724));
  AOI21_X1  g523(.A(G71gat), .B1(new_n715), .B2(new_n724), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n467), .A2(G71gat), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n715), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1334gat));
  NAND2_X1  g528(.A1(new_n715), .A2(new_n454), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G78gat), .ZN(G1335gat));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n624), .A2(new_n554), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n591), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n713), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n680), .A2(KEYINPUT51), .A3(new_n591), .A4(new_n733), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n737), .A2(new_n557), .A3(new_n447), .A4(new_n642), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n733), .A2(new_n642), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n678), .B2(new_n682), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n740), .A2(new_n447), .ZN(new_n741));
  OAI211_X1 g540(.A(KEYINPUT114), .B(new_n738), .C1(new_n741), .C2(new_n557), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT114), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n557), .B1(new_n740), .B2(new_n447), .ZN(new_n744));
  INV_X1    g543(.A(new_n738), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n742), .A2(new_n746), .ZN(G1336gat));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n643), .A2(new_n434), .A3(G92gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n737), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n740), .A2(new_n448), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n748), .B(new_n750), .C1(new_n751), .C2(new_n559), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n559), .B1(new_n740), .B2(new_n448), .ZN(new_n753));
  INV_X1    g552(.A(new_n750), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT52), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(G1337gat));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n467), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G99gat), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n455), .A2(new_n643), .A3(G99gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n737), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1338gat));
  NOR3_X1   g560(.A1(new_n459), .A2(G106gat), .A3(new_n643), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n735), .B2(new_n736), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT53), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n764), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n740), .A2(new_n454), .ZN(new_n768));
  INV_X1    g567(.A(G106gat), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n766), .B(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(KEYINPUT115), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n769), .B1(new_n740), .B2(new_n454), .ZN(new_n772));
  OAI211_X1 g571(.A(KEYINPUT53), .B(new_n771), .C1(new_n772), .C2(new_n764), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(G1339gat));
  INV_X1    g573(.A(new_n447), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n775), .A2(new_n448), .A3(new_n455), .ZN(new_n776));
  OR4_X1    g575(.A1(new_n632), .A2(new_n628), .A3(new_n631), .A4(new_n571), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(KEYINPUT54), .A3(new_n633), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779));
  OAI221_X1 g578(.A(new_n779), .B1(new_n632), .B2(new_n571), .C1(new_n628), .C2(new_n631), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n780), .A2(new_n781), .A3(new_n639), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n781), .B1(new_n780), .B2(new_n639), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n778), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n529), .B1(new_n527), .B2(new_n536), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n787), .A2(KEYINPUT117), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(KEYINPUT117), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n788), .B(new_n789), .C1(new_n540), .C2(new_n541), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n549), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n786), .A2(new_n553), .A3(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n778), .B(KEYINPUT55), .C1(new_n782), .C2(new_n783), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n793), .A2(new_n641), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n792), .A2(new_n591), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n791), .A2(new_n642), .A3(new_n553), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n786), .A2(new_n554), .A3(new_n641), .A4(new_n793), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n591), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT118), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n792), .A2(new_n591), .A3(new_n794), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n797), .A2(new_n796), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n800), .B(new_n801), .C1(new_n802), .C2(new_n591), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n799), .A2(new_n803), .A3(new_n623), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n644), .A2(new_n554), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT119), .B1(new_n807), .B2(new_n459), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809));
  AOI211_X1 g608(.A(new_n809), .B(new_n454), .C1(new_n804), .C2(new_n806), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n776), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(KEYINPUT120), .B(new_n776), .C1(new_n808), .C2(new_n810), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n554), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(G113gat), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n807), .A2(new_n456), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n817), .A2(new_n447), .A3(new_n434), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n319), .A2(new_n320), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n819), .A3(new_n554), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n820), .ZN(G1340gat));
  AOI21_X1  g620(.A(G120gat), .B1(new_n818), .B2(new_n642), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n813), .A2(new_n814), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n643), .A2(new_n323), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(G1341gat));
  NAND3_X1  g624(.A1(new_n813), .A2(new_n624), .A3(new_n814), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G127gat), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n818), .A2(new_n327), .A3(new_n624), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(G1342gat));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n591), .A3(new_n814), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G134gat), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n592), .A2(new_n448), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n817), .A2(new_n325), .A3(new_n447), .A4(new_n832), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT56), .Z(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n834), .ZN(G1343gat));
  NOR2_X1   g634(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT122), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n775), .A2(new_n467), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n434), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n801), .B1(new_n802), .B2(new_n591), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n624), .B1(new_n842), .B2(KEYINPUT118), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n805), .B1(new_n843), .B2(new_n803), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n841), .B1(new_n844), .B2(new_n459), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n623), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n806), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n459), .A2(new_n841), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n840), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n228), .B1(new_n850), .B2(new_n554), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n844), .A2(new_n459), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n555), .A2(G141gat), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n852), .A2(new_n434), .A3(new_n839), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n838), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n228), .ZN(new_n858));
  INV_X1    g657(.A(new_n840), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT57), .B1(new_n807), .B2(new_n454), .ZN(new_n860));
  INV_X1    g659(.A(new_n849), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n858), .B1(new_n862), .B2(new_n555), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n863), .A2(new_n855), .A3(new_n854), .A4(new_n837), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n857), .A2(new_n864), .ZN(G1344gat));
  AND2_X1   g664(.A1(new_n852), .A2(new_n839), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n866), .A2(new_n434), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n237), .A3(new_n642), .ZN(new_n868));
  AOI211_X1 g667(.A(KEYINPUT59), .B(new_n237), .C1(new_n850), .C2(new_n642), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n807), .A2(new_n848), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT57), .B1(new_n847), .B2(new_n454), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n642), .B(new_n859), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n870), .B1(new_n873), .B2(G148gat), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n868), .B1(new_n869), .B2(new_n874), .ZN(G1345gat));
  NAND3_X1  g674(.A1(new_n867), .A2(new_n222), .A3(new_n624), .ZN(new_n876));
  OAI21_X1  g675(.A(G155gat), .B1(new_n862), .B2(new_n623), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1346gat));
  OAI21_X1  g677(.A(G162gat), .B1(new_n862), .B2(new_n592), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n866), .A2(new_n223), .A3(new_n832), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1347gat));
  NOR2_X1   g680(.A1(new_n447), .A2(new_n434), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n817), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(G169gat), .B1(new_n883), .B2(new_n554), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n882), .B(KEYINPUT123), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n724), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n809), .B1(new_n844), .B2(new_n454), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n807), .A2(KEYINPUT119), .A3(new_n459), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n555), .A2(new_n286), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n884), .B1(new_n889), .B2(new_n890), .ZN(G1348gat));
  AOI21_X1  g690(.A(G176gat), .B1(new_n883), .B2(new_n642), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n643), .A2(new_n300), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n889), .B2(new_n893), .ZN(G1349gat));
  AOI21_X1  g693(.A(new_n293), .B1(new_n889), .B2(new_n624), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n623), .A2(new_n305), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n807), .A2(new_n456), .A3(new_n882), .A4(new_n896), .ZN(new_n897));
  XOR2_X1   g696(.A(new_n897), .B(KEYINPUT124), .Z(new_n898));
  OAI21_X1  g697(.A(KEYINPUT60), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT60), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n897), .B(KEYINPUT124), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n623), .B(new_n886), .C1(new_n887), .C2(new_n888), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n900), .B(new_n901), .C1(new_n902), .C2(new_n293), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n899), .A2(new_n903), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n883), .A2(new_n294), .A3(new_n591), .ZN(new_n905));
  INV_X1    g704(.A(new_n886), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n591), .B(new_n906), .C1(new_n808), .C2(new_n810), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n907), .A2(new_n908), .A3(G190gat), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n907), .B2(G190gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(G1351gat));
  INV_X1    g710(.A(G197gat), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n885), .A2(new_n655), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n554), .B(new_n913), .C1(new_n871), .C2(new_n872), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n914), .B2(KEYINPUT125), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(KEYINPUT125), .B2(new_n914), .ZN(new_n916));
  NOR4_X1   g715(.A1(new_n467), .A2(new_n459), .A3(new_n447), .A4(new_n434), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n807), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n912), .A3(new_n554), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n916), .A2(new_n920), .ZN(G1352gat));
  NOR3_X1   g720(.A1(new_n918), .A2(G204gat), .A3(new_n643), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT62), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n642), .B(new_n913), .C1(new_n871), .C2(new_n872), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G204gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1353gat));
  NAND3_X1  g725(.A1(new_n919), .A2(new_n209), .A3(new_n624), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n624), .B(new_n913), .C1(new_n871), .C2(new_n872), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT63), .B1(new_n928), .B2(G211gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(G1354gat));
  NOR2_X1   g730(.A1(new_n592), .A2(new_n210), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n913), .B(new_n932), .C1(new_n871), .C2(new_n872), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n807), .A2(new_n591), .A3(new_n917), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n934), .A2(new_n935), .A3(new_n210), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n934), .B2(new_n210), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


