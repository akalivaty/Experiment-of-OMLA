//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n797, new_n798, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(G22gat), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  AND2_X1   g005(.A1(G211gat), .A2(G218gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(KEYINPUT22), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n205), .B1(new_n210), .B2(KEYINPUT29), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n212));
  INV_X1    g011(.A(G141gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G148gat), .ZN(new_n214));
  INV_X1    g013(.A(G148gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(G141gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(G141gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(G148gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT79), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n217), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT78), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT78), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(G155gat), .A3(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n222), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT80), .B(G155gat), .ZN(new_n232));
  INV_X1    g031(.A(G162gat), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT2), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n219), .A2(new_n220), .B1(new_n228), .B2(new_n223), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n211), .A2(new_n237), .ZN(new_n238));
  AOI221_X4 g037(.A(KEYINPUT3), .B1(new_n234), .B2(new_n235), .C1(new_n222), .C2(new_n230), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(KEYINPUT29), .ZN(new_n240));
  INV_X1    g039(.A(new_n210), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n238), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G228gat), .A2(G233gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT88), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(KEYINPUT88), .A3(new_n243), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT31), .B(G50gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n243), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n210), .B(KEYINPUT75), .Z(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n238), .B(new_n251), .C1(new_n253), .C2(new_n240), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n248), .A2(new_n250), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n250), .B1(new_n248), .B2(new_n254), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n204), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n257), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n259), .A2(new_n203), .A3(new_n255), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n263));
  AOI21_X1  g062(.A(G190gat), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT66), .B1(new_n264), .B2(new_n267), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(KEYINPUT28), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G183gat), .ZN(new_n273));
  INV_X1    g072(.A(G190gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G169gat), .ZN(new_n277));
  INV_X1    g076(.A(G176gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT26), .ZN(new_n280));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT26), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n272), .A2(new_n276), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT23), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT23), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n286), .A2(new_n287), .A3(new_n281), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT24), .ZN(new_n289));
  NOR2_X1   g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290));
  OR3_X1    g089(.A1(new_n275), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(G183gat), .A3(G190gat), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n288), .A2(KEYINPUT25), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT64), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT25), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n286), .A2(new_n292), .A3(new_n287), .A4(new_n281), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n275), .A2(new_n289), .A3(new_n290), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n293), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n294), .B1(new_n293), .B2(new_n298), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n284), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n302));
  INV_X1    g101(.A(G120gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G113gat), .ZN(new_n304));
  INV_X1    g103(.A(G113gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G120gat), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n302), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G127gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G134gat), .ZN(new_n310));
  INV_X1    g109(.A(G134gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G127gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n304), .A2(new_n306), .A3(new_n302), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n308), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT67), .B(G134gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n310), .B1(new_n318), .B2(new_n309), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT1), .B1(new_n304), .B2(new_n306), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n301), .A2(new_n323), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n304), .A2(new_n306), .A3(new_n302), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n325), .A2(new_n307), .A3(new_n314), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT67), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(G134gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n311), .A2(KEYINPUT67), .ZN(new_n329));
  OAI21_X1  g128(.A(G127gat), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n320), .B1(new_n330), .B2(new_n310), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n284), .B(new_n332), .C1(new_n299), .C2(new_n300), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n324), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G227gat), .A2(G233gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n337), .A2(KEYINPUT34), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(KEYINPUT34), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(KEYINPUT74), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT32), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT33), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT69), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n334), .B2(new_n336), .ZN(new_n344));
  AOI211_X1 g143(.A(KEYINPUT69), .B(new_n335), .C1(new_n324), .C2(new_n333), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G15gat), .B(G43gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(G71gat), .B(G99gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n341), .B1(new_n351), .B2(KEYINPUT33), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(new_n344), .B2(new_n345), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT72), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n356), .B(new_n353), .C1(new_n344), .C2(new_n345), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n340), .A2(new_n352), .A3(new_n355), .A4(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT74), .B1(new_n338), .B2(new_n339), .ZN(new_n359));
  OR2_X1    g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n359), .ZN(new_n361));
  AOI211_X1 g160(.A(KEYINPUT35), .B(new_n261), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT87), .B(KEYINPUT6), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(KEYINPUT86), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n222), .A2(new_n230), .B1(new_n234), .B2(new_n235), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n332), .A2(new_n365), .A3(KEYINPUT4), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT4), .B1(new_n365), .B2(new_n332), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n367), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n205), .B1(new_n231), .B2(new_n236), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n239), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT81), .B1(new_n326), .B2(new_n331), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n317), .A2(new_n322), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n372), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT79), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT79), .B1(new_n219), .B2(new_n220), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n229), .B1(new_n382), .B2(new_n218), .ZN(new_n383));
  INV_X1    g182(.A(new_n236), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT3), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n365), .A2(new_n205), .ZN(new_n386));
  AND4_X1   g185(.A1(new_n372), .A2(new_n378), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n371), .B1(new_n379), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT83), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT5), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n378), .A2(new_n237), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n323), .B2(new_n237), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n391), .B1(new_n393), .B2(new_n370), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n371), .B(KEYINPUT83), .C1(new_n379), .C2(new_n387), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n379), .A2(new_n387), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT85), .ZN(new_n398));
  INV_X1    g197(.A(new_n368), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n399), .B2(new_n366), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT85), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n397), .A2(new_n402), .A3(new_n391), .A4(new_n369), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(G1gat), .B(G29gat), .Z(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G57gat), .B(G85gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n364), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n403), .A3(new_n409), .ZN(new_n412));
  INV_X1    g211(.A(new_n363), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n409), .B1(new_n396), .B2(new_n403), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n412), .B(new_n413), .C1(new_n416), .C2(new_n364), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G226gat), .A2(G233gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n293), .A2(new_n298), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n284), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n419), .B1(new_n421), .B2(KEYINPUT29), .ZN(new_n422));
  INV_X1    g221(.A(new_n419), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n301), .A2(KEYINPUT76), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT76), .B1(new_n301), .B2(new_n423), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n241), .B(new_n422), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT29), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n301), .A2(new_n427), .A3(new_n419), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n284), .A2(new_n423), .A3(new_n420), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n252), .A3(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G8gat), .B(G36gat), .ZN(new_n431));
  INV_X1    g230(.A(G64gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G92gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n426), .A2(new_n430), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n426), .A2(new_n430), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n439), .B1(new_n440), .B2(new_n435), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT77), .ZN(new_n442));
  INV_X1    g241(.A(new_n437), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n442), .B1(new_n443), .B2(KEYINPUT30), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n437), .A2(KEYINPUT77), .A3(new_n438), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n418), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n362), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n352), .A2(new_n355), .A3(new_n357), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n338), .A2(new_n339), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(KEYINPUT73), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n449), .A2(new_n451), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n452), .A2(new_n453), .A3(new_n261), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n447), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n448), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n393), .A2(new_n370), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT89), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT89), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n397), .A2(new_n402), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n461), .B2(new_n370), .ZN(new_n462));
  OAI211_X1 g261(.A(KEYINPUT39), .B(new_n459), .C1(new_n462), .C2(new_n458), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT39), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n461), .A2(new_n464), .A3(new_n370), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n409), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT40), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n416), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n463), .A2(KEYINPUT40), .A3(new_n409), .A4(new_n465), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n468), .A2(new_n446), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n261), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT90), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n475), .A2(new_n210), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n252), .B1(new_n428), .B2(new_n429), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT37), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n440), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT37), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT38), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n478), .A2(new_n481), .A3(new_n482), .A4(new_n435), .ZN(new_n483));
  AND4_X1   g282(.A1(new_n474), .A2(new_n418), .A3(new_n437), .A4(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n443), .B1(new_n415), .B2(new_n417), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n474), .B1(new_n485), .B2(new_n483), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n481), .A2(new_n435), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n479), .A2(new_n480), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT38), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n473), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT36), .ZN(new_n492));
  INV_X1    g291(.A(new_n361), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n358), .A2(new_n359), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n261), .B1(new_n418), .B2(new_n446), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT36), .B1(new_n452), .B2(new_n453), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n457), .B1(new_n491), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G29gat), .A2(G36gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT91), .ZN(new_n501));
  OR3_X1    g300(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G43gat), .B(G50gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(KEYINPUT15), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n506), .B(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT92), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n509), .B(new_n501), .C1(new_n510), .C2(new_n502), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n504), .A2(KEYINPUT92), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT16), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(G1gat), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(G1gat), .B2(new_n514), .ZN(new_n517));
  INV_X1    g316(.A(G8gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n513), .B(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G229gat), .A2(G233gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT13), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT93), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n517), .B(G8gat), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n513), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n513), .B(KEYINPUT17), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(new_n519), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n521), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT18), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n528), .A2(KEYINPUT18), .A3(new_n521), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n524), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT11), .B(G169gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(G197gat), .ZN(new_n536));
  XOR2_X1   g335(.A(G113gat), .B(G141gat), .Z(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT12), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n539), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n533), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G71gat), .B(G78gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT94), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT9), .ZN(new_n547));
  INV_X1    g346(.A(G71gat), .ZN(new_n548));
  INV_X1    g347(.A(G78gat), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n432), .A2(G57gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n432), .A2(G57gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(KEYINPUT95), .B(G57gat), .Z(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(new_n432), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n550), .B1(new_n556), .B2(new_n551), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n544), .B(KEYINPUT96), .Z(new_n558));
  OAI21_X1  g357(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT21), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n519), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G183gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(G231gat), .A2(G233gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G211gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n564), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n559), .A2(new_n560), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n568), .B(new_n569), .Z(new_n570));
  OR2_X1    g369(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n570), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G85gat), .A2(G92gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT7), .ZN(new_n575));
  INV_X1    g374(.A(G99gat), .ZN(new_n576));
  INV_X1    g375(.A(G106gat), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT8), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n575), .B(new_n578), .C1(G85gat), .C2(G92gat), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT98), .Z(new_n580));
  XOR2_X1   g379(.A(G99gat), .B(G106gat), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n579), .B(KEYINPUT98), .ZN(new_n583));
  INV_X1    g382(.A(new_n581), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n527), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n585), .ZN(new_n587));
  AND2_X1   g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n587), .A2(new_n513), .B1(KEYINPUT41), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G134gat), .B(G162gat), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT97), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n590), .B(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n588), .A2(KEYINPUT41), .ZN(new_n594));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n593), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n573), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G230gat), .ZN(new_n599));
  INV_X1    g398(.A(G233gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n559), .ZN(new_n602));
  INV_X1    g401(.A(new_n585), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n583), .A2(new_n584), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT10), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n582), .A2(new_n585), .A3(new_n559), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n587), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n601), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI211_X1 g409(.A(new_n599), .B(new_n600), .C1(new_n605), .C2(new_n607), .ZN(new_n611));
  XNOR2_X1  g410(.A(G120gat), .B(G148gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G176gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G204gat), .ZN(new_n614));
  OR3_X1    g413(.A1(new_n610), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n614), .B1(new_n610), .B2(new_n611), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(KEYINPUT99), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT99), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n618), .B(new_n614), .C1(new_n610), .C2(new_n611), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n598), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n499), .A2(new_n543), .A3(new_n622), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n623), .A2(KEYINPUT100), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(KEYINPUT100), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n418), .B(KEYINPUT101), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT102), .B(G1gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(G1324gat));
  INV_X1    g429(.A(new_n446), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(new_n624), .B2(new_n625), .ZN(new_n632));
  NAND2_X1  g431(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n515), .A2(new_n518), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT42), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n632), .A2(KEYINPUT42), .A3(new_n633), .A4(new_n634), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n637), .B(new_n638), .C1(new_n518), .C2(new_n632), .ZN(G1325gat));
  NOR2_X1   g438(.A1(new_n493), .A2(new_n494), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(G15gat), .B1(new_n626), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n495), .ZN(new_n643));
  INV_X1    g442(.A(new_n497), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n646), .A2(KEYINPUT103), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(KEYINPUT103), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n624), .B2(new_n625), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n642), .B1(G15gat), .B2(new_n651), .ZN(G1326gat));
  NAND2_X1  g451(.A1(new_n626), .A2(new_n261), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT43), .B(G22gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  INV_X1    g454(.A(new_n597), .ZN(new_n656));
  INV_X1    g455(.A(new_n543), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n573), .A2(new_n657), .A3(new_n621), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n499), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n627), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n659), .A2(G29gat), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(KEYINPUT45), .Z(new_n662));
  NAND4_X1  g461(.A1(new_n499), .A2(KEYINPUT104), .A3(KEYINPUT44), .A4(new_n656), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n418), .A2(new_n437), .A3(new_n483), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT90), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n485), .A2(new_n474), .A3(new_n483), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n490), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n473), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n498), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n447), .A2(new_n362), .B1(new_n455), .B2(KEYINPUT35), .ZN(new_n670));
  OAI211_X1 g469(.A(KEYINPUT104), .B(new_n656), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n663), .A2(new_n673), .A3(new_n658), .ZN(new_n674));
  OAI21_X1  g473(.A(G29gat), .B1(new_n674), .B2(new_n660), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n662), .A2(new_n675), .ZN(G1328gat));
  NOR3_X1   g475(.A1(new_n659), .A2(G36gat), .A3(new_n631), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT46), .ZN(new_n678));
  OAI21_X1  g477(.A(G36gat), .B1(new_n674), .B2(new_n631), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(G1329gat));
  OAI21_X1  g479(.A(G43gat), .B1(new_n674), .B2(new_n645), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n659), .A2(G43gat), .A3(new_n640), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n681), .A2(new_n683), .A3(KEYINPUT47), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n663), .A2(new_n673), .A3(new_n649), .A4(new_n658), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n685), .A2(KEYINPUT105), .A3(G43gat), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT105), .B1(new_n685), .B2(G43gat), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n686), .A2(new_n687), .A3(new_n682), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n684), .B1(new_n688), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g488(.A(G50gat), .B1(new_n674), .B2(new_n472), .ZN(new_n690));
  OR3_X1    g489(.A1(new_n659), .A2(G50gat), .A3(new_n472), .ZN(new_n691));
  OR2_X1    g490(.A1(KEYINPUT106), .A2(KEYINPUT48), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(KEYINPUT106), .A2(KEYINPUT48), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1331gat));
  NOR2_X1   g494(.A1(new_n669), .A2(new_n670), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n543), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n598), .A2(new_n620), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n627), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(new_n555), .ZN(G1332gat));
  INV_X1    g501(.A(KEYINPUT49), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n432), .ZN(new_n704));
  NAND2_X1  g503(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n700), .A2(new_n446), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n703), .B(new_n432), .C1(new_n699), .C2(new_n631), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT107), .B(KEYINPUT108), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1333gat));
  NAND3_X1  g509(.A1(new_n700), .A2(new_n548), .A3(new_n641), .ZN(new_n711));
  OAI21_X1  g510(.A(G71gat), .B1(new_n699), .B2(new_n650), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n472), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT109), .B(G78gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1335gat));
  NOR2_X1   g516(.A1(new_n573), .A2(new_n543), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n656), .B(new_n718), .C1(new_n669), .C2(new_n670), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT51), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n660), .A2(G85gat), .A3(new_n620), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n663), .A2(new_n673), .A3(new_n621), .A4(new_n718), .ZN(new_n726));
  OAI21_X1  g525(.A(G85gat), .B1(new_n726), .B2(new_n660), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(G1336gat));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729));
  OR3_X1    g528(.A1(new_n726), .A2(new_n729), .A3(new_n631), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n726), .B2(new_n631), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(G92gat), .A3(new_n731), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n721), .A2(new_n434), .A3(new_n446), .A4(new_n621), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n734));
  AND2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G92gat), .B1(new_n726), .B2(new_n631), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n733), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT52), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n739), .ZN(G1337gat));
  NAND4_X1  g539(.A1(new_n723), .A2(new_n576), .A3(new_n641), .A4(new_n621), .ZN(new_n741));
  OAI21_X1  g540(.A(G99gat), .B1(new_n726), .B2(new_n650), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1338gat));
  OAI21_X1  g542(.A(G106gat), .B1(new_n726), .B2(new_n472), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT113), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n472), .A2(G106gat), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n721), .A2(new_n621), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n745), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n744), .B(new_n747), .C1(KEYINPUT113), .C2(KEYINPUT53), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(G1339gat));
  NAND2_X1  g551(.A1(new_n622), .A2(new_n657), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n608), .A2(new_n609), .A3(new_n601), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT54), .ZN(new_n755));
  OR3_X1    g554(.A1(new_n754), .A2(new_n610), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n610), .A2(new_n755), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n757), .A2(KEYINPUT114), .A3(new_n614), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT114), .B1(new_n757), .B2(new_n614), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OR3_X1    g561(.A1(new_n528), .A2(KEYINPUT115), .A3(new_n521), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n520), .A2(new_n522), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT116), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT115), .B1(new_n528), .B2(new_n521), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n763), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n534), .A2(new_n539), .B1(new_n767), .B2(new_n538), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT55), .B(new_n756), .C1(new_n758), .C2(new_n759), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n762), .A2(new_n768), .A3(new_n615), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n597), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n762), .A2(new_n543), .A3(new_n615), .A4(new_n769), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n621), .A2(new_n773), .A3(new_n768), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n767), .A2(new_n538), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n540), .A2(new_n617), .A3(new_n619), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT117), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n772), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n771), .B1(new_n597), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n753), .B1(new_n779), .B2(new_n573), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT118), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n782), .B(new_n753), .C1(new_n779), .C2(new_n573), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n781), .A2(new_n627), .A3(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n784), .A2(new_n454), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(new_n631), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n543), .A2(new_n305), .ZN(new_n787));
  XOR2_X1   g586(.A(new_n787), .B(KEYINPUT119), .Z(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n640), .A2(new_n261), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n784), .A2(new_n631), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G113gat), .B1(new_n791), .B2(new_n657), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(G1340gat));
  NAND3_X1  g592(.A1(new_n786), .A2(new_n303), .A3(new_n621), .ZN(new_n794));
  OAI21_X1  g593(.A(G120gat), .B1(new_n791), .B2(new_n620), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(G1341gat));
  INV_X1    g595(.A(new_n573), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n791), .A2(new_n309), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n785), .A2(new_n631), .A3(new_n573), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n798), .B1(new_n799), .B2(new_n309), .ZN(G1342gat));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n597), .A2(new_n318), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n784), .A2(new_n631), .A3(new_n454), .A4(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n801), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  OAI21_X1  g606(.A(G134gat), .B1(new_n791), .B2(new_n597), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n803), .A2(KEYINPUT120), .A3(KEYINPUT56), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n806), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(G1343gat));
  NOR2_X1   g609(.A1(new_n657), .A2(G141gat), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n647), .A2(new_n261), .A3(new_n648), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT121), .B1(new_n784), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n781), .A2(new_n627), .A3(new_n783), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n815), .A2(new_n816), .A3(new_n812), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n631), .B(new_n811), .C1(new_n814), .C2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n781), .A2(new_n820), .A3(new_n261), .A4(new_n783), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n645), .A2(new_n631), .A3(new_n627), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n656), .B1(new_n772), .B2(new_n776), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n797), .B1(new_n823), .B2(new_n771), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n753), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n261), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n822), .B1(new_n826), .B2(KEYINPUT57), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n821), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(G141gat), .B1(new_n828), .B2(new_n657), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n818), .A2(new_n819), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n784), .A2(new_n631), .A3(new_n811), .A4(new_n813), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT58), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(G1344gat));
  NOR2_X1   g633(.A1(new_n620), .A2(G148gat), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n631), .B(new_n835), .C1(new_n814), .C2(new_n817), .ZN(new_n836));
  INV_X1    g635(.A(new_n828), .ZN(new_n837));
  AOI211_X1 g636(.A(KEYINPUT59), .B(new_n215), .C1(new_n837), .C2(new_n621), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n781), .A2(new_n783), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT57), .B1(new_n840), .B2(new_n472), .ZN(new_n841));
  INV_X1    g640(.A(new_n822), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n820), .A3(new_n261), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n841), .A2(new_n621), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n839), .B1(new_n844), .B2(G148gat), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n836), .B1(new_n838), .B2(new_n845), .ZN(G1345gat));
  OAI211_X1 g645(.A(new_n631), .B(new_n573), .C1(new_n814), .C2(new_n817), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n797), .A2(new_n232), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT122), .Z(new_n849));
  AOI22_X1  g648(.A1(new_n847), .A2(new_n232), .B1(new_n837), .B2(new_n849), .ZN(G1346gat));
  NOR3_X1   g649(.A1(new_n828), .A2(new_n233), .A3(new_n597), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n631), .B(new_n656), .C1(new_n814), .C2(new_n817), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n233), .ZN(G1347gat));
  NAND4_X1  g652(.A1(new_n781), .A2(new_n446), .A3(new_n660), .A4(new_n783), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n454), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n277), .A3(new_n543), .ZN(new_n858));
  INV_X1    g657(.A(new_n790), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n543), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n861), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT123), .B1(new_n861), .B2(G169gat), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(G1348gat));
  NOR4_X1   g663(.A1(new_n854), .A2(new_n278), .A3(new_n859), .A4(new_n620), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n857), .A2(new_n621), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(new_n278), .ZN(G1349gat));
  NAND2_X1  g666(.A1(new_n262), .A2(new_n263), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n573), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n854), .A2(new_n859), .A3(new_n797), .ZN(new_n870));
  OAI22_X1  g669(.A1(new_n856), .A2(new_n869), .B1(new_n870), .B2(new_n273), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT60), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n873));
  OAI221_X1 g672(.A(new_n873), .B1(new_n870), .B2(new_n273), .C1(new_n856), .C2(new_n869), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(G1350gat));
  NOR3_X1   g674(.A1(new_n854), .A2(new_n859), .A3(new_n597), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n274), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT61), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n877), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n857), .A2(new_n274), .A3(new_n656), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n878), .B(new_n879), .C1(new_n876), .C2(new_n274), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G1351gat));
  NOR3_X1   g684(.A1(new_n649), .A2(new_n631), .A3(new_n627), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n841), .A2(new_n843), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(G197gat), .B1(new_n887), .B2(new_n657), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n854), .A2(G197gat), .A3(new_n812), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n889), .A2(KEYINPUT125), .A3(new_n543), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT125), .B1(new_n889), .B2(new_n543), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(G1352gat));
  NOR3_X1   g691(.A1(new_n854), .A2(G204gat), .A3(new_n812), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n621), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT126), .B1(new_n894), .B2(KEYINPUT62), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(KEYINPUT62), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n841), .A2(new_n621), .A3(new_n843), .A4(new_n886), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G204gat), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n893), .A2(new_n899), .A3(new_n900), .A4(new_n621), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n895), .A2(new_n896), .A3(new_n898), .A4(new_n901), .ZN(G1353gat));
  NOR2_X1   g701(.A1(new_n854), .A2(new_n812), .ZN(new_n903));
  INV_X1    g702(.A(G211gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n904), .A3(new_n573), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n841), .A2(new_n573), .A3(new_n843), .A4(new_n886), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n906), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT63), .B1(new_n906), .B2(G211gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(G1354gat));
  AOI21_X1  g708(.A(G218gat), .B1(new_n903), .B2(new_n656), .ZN(new_n910));
  INV_X1    g709(.A(new_n887), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n656), .A2(G218gat), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT127), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n910), .B1(new_n911), .B2(new_n913), .ZN(G1355gat));
endmodule


