//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1236, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  INV_X1    g0006(.A(G244), .ZN(new_n207));
  INV_X1    g0007(.A(G116), .ZN(new_n208));
  INV_X1    g0008(.A(G270), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n210), .B(new_n215), .C1(G68), .C2(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n201), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n228), .A2(new_n229), .A3(G50), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n222), .A2(G13), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n231), .B(G250), .C1(G257), .C2(G264), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT0), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n225), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT66), .Z(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n217), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n209), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(new_n208), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NAND2_X1  g0051(.A1(new_n203), .A2(G20), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G150), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n252), .B(new_n254), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n226), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n202), .ZN(new_n266));
  INV_X1    g0066(.A(new_n261), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n263), .A2(G20), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n262), .B(new_n266), .C1(new_n202), .C2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT70), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(G222), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G223), .ZN(new_n280));
  OAI221_X1 g0080(.A(new_n278), .B1(new_n206), .B2(new_n276), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n226), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n263), .A2(G274), .ZN(new_n287));
  AND2_X1   g0087(.A1(KEYINPUT67), .A2(G41), .ZN(new_n288));
  NOR2_X1   g0088(.A1(KEYINPUT67), .A2(G41), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n287), .B1(new_n290), .B2(G45), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT68), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(new_n282), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G226), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n286), .A2(new_n291), .A3(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n272), .A2(KEYINPUT9), .B1(G200), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n300), .B(new_n302), .C1(KEYINPUT9), .C2(new_n272), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT13), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n276), .A2(G226), .A3(new_n277), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n276), .A2(G232), .A3(G1698), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G97), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n285), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n297), .A2(G238), .ZN(new_n313));
  AND4_X1   g0113(.A1(new_n307), .A2(new_n312), .A3(new_n291), .A4(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n290), .ZN(new_n315));
  INV_X1    g0115(.A(G45), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n311), .A2(new_n285), .B1(new_n317), .B2(new_n287), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n307), .B1(new_n318), .B2(new_n313), .ZN(new_n319));
  OAI21_X1  g0119(.A(G200), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n256), .A2(G77), .B1(new_n253), .B2(G50), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(new_n227), .B2(G68), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(KEYINPUT11), .A3(new_n261), .ZN(new_n323));
  INV_X1    g0123(.A(G68), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n269), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n264), .A2(G68), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT12), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT11), .B1(new_n322), .B2(new_n261), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n312), .A2(new_n291), .A3(new_n313), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT13), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n318), .A2(new_n307), .A3(new_n313), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(G190), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n320), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT71), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n320), .A2(new_n329), .A3(new_n333), .A4(KEYINPUT71), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(G169), .B1(new_n314), .B2(new_n319), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT14), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n331), .A2(G179), .A3(new_n332), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT14), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n342), .B(G169), .C1(new_n314), .C2(new_n319), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n329), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n338), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n299), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n270), .B1(new_n299), .B2(G179), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  XOR2_X1   g0152(.A(KEYINPUT15), .B(G87), .Z(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n253), .B(KEYINPUT69), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n354), .B1(new_n258), .B2(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(new_n261), .B1(new_n206), .B2(new_n265), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n206), .B2(new_n269), .ZN(new_n358));
  INV_X1    g0158(.A(G238), .ZN(new_n359));
  INV_X1    g0159(.A(G107), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n279), .A2(new_n359), .B1(new_n360), .B2(new_n276), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n274), .A2(new_n275), .ZN(new_n362));
  NOR3_X1   g0162(.A1(new_n362), .A2(new_n237), .A3(G1698), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n285), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n297), .A2(G244), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n291), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n358), .B1(new_n366), .B2(G179), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n366), .A2(new_n348), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n306), .A2(new_n347), .A3(new_n352), .A4(new_n370), .ZN(new_n371));
  OR2_X1    g0171(.A1(KEYINPUT72), .A2(G33), .ZN(new_n372));
  NAND2_X1  g0172(.A1(KEYINPUT72), .A2(G33), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n273), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT73), .B1(new_n255), .B2(KEYINPUT3), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(new_n273), .A3(G33), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n227), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT7), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(new_n227), .C1(new_n374), .C2(new_n378), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(G68), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G58), .A2(G68), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n227), .B1(new_n229), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n253), .A2(G159), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT74), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n384), .ZN(new_n389));
  OAI21_X1  g0189(.A(G20), .B1(new_n389), .B2(new_n201), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT74), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(new_n386), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  AND2_X1   g0196(.A1(KEYINPUT72), .A2(G33), .ZN(new_n397));
  NOR2_X1   g0197(.A1(KEYINPUT72), .A2(G33), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT3), .ZN(new_n399));
  INV_X1    g0199(.A(new_n275), .ZN(new_n400));
  OAI211_X1 g0200(.A(KEYINPUT7), .B(new_n227), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT7), .B1(new_n362), .B2(new_n227), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n324), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n396), .B1(new_n404), .B2(new_n393), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n395), .A2(new_n261), .A3(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n375), .A2(new_n377), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT3), .B1(new_n397), .B2(new_n398), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n217), .A2(G1698), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n280), .A2(new_n277), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n407), .A2(new_n408), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n284), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT76), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n295), .A2(G232), .A3(new_n296), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n291), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n414), .A3(new_n291), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n413), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OR2_X1    g0219(.A1(KEYINPUT77), .A2(G190), .ZN(new_n420));
  NAND2_X1  g0220(.A1(KEYINPUT77), .A2(G190), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n258), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n268), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT75), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n265), .A2(new_n261), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n427), .A2(new_n428), .B1(new_n265), .B2(new_n258), .ZN(new_n429));
  INV_X1    g0229(.A(new_n418), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(new_n416), .ZN(new_n431));
  OAI21_X1  g0231(.A(G200), .B1(new_n431), .B2(new_n413), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n406), .A2(new_n424), .A3(new_n429), .A4(new_n432), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n433), .A2(KEYINPUT17), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(KEYINPUT17), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n406), .A2(new_n429), .ZN(new_n436));
  INV_X1    g0236(.A(new_n413), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(G179), .C1(new_n416), .C2(new_n430), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n348), .B2(new_n419), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n436), .A2(KEYINPUT18), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT18), .B1(new_n436), .B2(new_n439), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n434), .A2(new_n435), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n366), .A2(new_n301), .ZN(new_n443));
  AOI211_X1 g0243(.A(new_n358), .B(new_n443), .C1(G200), .C2(new_n366), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n371), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n260), .A2(new_n226), .B1(G20), .B2(new_n208), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G283), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n447), .B(new_n227), .C1(G33), .C2(new_n213), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT86), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n446), .A2(new_n448), .B1(new_n449), .B2(KEYINPUT20), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n449), .B2(KEYINPUT20), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT20), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n446), .A2(KEYINPUT86), .A3(new_n448), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n265), .A2(new_n208), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n263), .A2(G33), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n428), .A2(G116), .A3(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n451), .A2(new_n453), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n457), .A2(G169), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT67), .ZN(new_n459));
  INV_X1    g0259(.A(G41), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT5), .ZN(new_n462));
  NAND2_X1  g0262(.A1(KEYINPUT67), .A2(G41), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n263), .A2(G45), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n460), .A2(KEYINPUT5), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n468), .A2(G270), .A3(new_n295), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n464), .A2(G274), .A3(new_n466), .A4(new_n467), .ZN(new_n470));
  INV_X1    g0270(.A(new_n295), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT85), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n362), .A2(G303), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n214), .A2(new_n277), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n407), .A2(new_n408), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n277), .A2(G264), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n285), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n465), .B1(new_n290), .B2(new_n462), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n480), .A2(G274), .A3(new_n295), .A4(new_n467), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n468), .A2(G270), .A3(new_n295), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT85), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n473), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n458), .A2(new_n485), .A3(KEYINPUT21), .ZN(new_n486));
  INV_X1    g0286(.A(G179), .ZN(new_n487));
  INV_X1    g0287(.A(new_n457), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT21), .B1(new_n458), .B2(new_n485), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n486), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n211), .A2(G20), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n407), .A2(KEYINPUT22), .A3(new_n408), .A4(new_n492), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n397), .A2(new_n398), .A3(new_n208), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n274), .A3(new_n275), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT22), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n227), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n227), .A2(G107), .ZN(new_n498));
  XNOR2_X1  g0298(.A(new_n498), .B(KEYINPUT23), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n493), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT87), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT87), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n493), .A2(new_n497), .A3(new_n502), .A4(new_n499), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(KEYINPUT24), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT24), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n500), .A2(KEYINPUT87), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n261), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n267), .A2(new_n264), .A3(new_n455), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G107), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n264), .A2(G107), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n511), .B(KEYINPUT25), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n507), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n214), .A2(G1698), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n212), .A2(new_n277), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n407), .A2(new_n408), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n372), .A2(G294), .A3(new_n373), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n284), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n468), .A2(G264), .A3(new_n295), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n519), .A2(new_n481), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT88), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n468), .A2(KEYINPUT88), .A3(G264), .A4(new_n295), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n519), .A2(new_n481), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n521), .A2(new_n348), .B1(new_n525), .B2(new_n487), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n513), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G200), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n519), .A2(new_n301), .A3(new_n481), .A4(new_n520), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n531), .A2(new_n510), .A3(new_n507), .A4(new_n512), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n485), .A2(G200), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n533), .B(new_n488), .C1(new_n485), .C2(new_n422), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n491), .A2(new_n527), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n468), .A2(G257), .A3(new_n295), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n481), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n207), .A2(G1698), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n408), .A2(new_n375), .A3(new_n377), .A4(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT4), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n540), .A2(KEYINPUT79), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT79), .B1(new_n540), .B2(new_n541), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n276), .A2(G250), .A3(G1698), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n276), .A2(KEYINPUT4), .A3(new_n539), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n545), .A3(new_n447), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(G190), .B(new_n538), .C1(new_n547), .C2(new_n284), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n265), .A2(new_n213), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n508), .B2(new_n213), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n253), .A2(G77), .ZN(new_n551));
  NAND2_X1  g0351(.A1(KEYINPUT6), .A2(G97), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT78), .B1(new_n552), .B2(G107), .ZN(new_n553));
  OR3_X1    g0353(.A1(new_n552), .A2(KEYINPUT78), .A3(G107), .ZN(new_n554));
  XOR2_X1   g0354(.A(G97), .B(G107), .Z(new_n555));
  OAI211_X1 g0355(.A(new_n553), .B(new_n554), .C1(new_n555), .C2(KEYINPUT6), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G20), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n372), .A2(new_n273), .A3(new_n373), .ZN(new_n558));
  AOI21_X1  g0358(.A(G20), .B1(new_n558), .B2(new_n275), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n402), .B1(new_n559), .B2(KEYINPUT7), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n551), .B(new_n557), .C1(new_n560), .C2(new_n360), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n550), .B1(new_n561), .B2(new_n261), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n548), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT80), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n481), .A2(new_n536), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n564), .B1(new_n481), .B2(new_n536), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n540), .A2(new_n541), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT79), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n544), .A2(new_n545), .A3(new_n447), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n540), .A2(KEYINPUT79), .A3(new_n541), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n285), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n528), .B1(new_n568), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT81), .B1(new_n563), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n257), .B2(new_n213), .ZN(new_n579));
  XNOR2_X1  g0379(.A(KEYINPUT83), .B(G87), .ZN(new_n580));
  NOR2_X1   g0380(.A1(G97), .A2(G107), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n227), .B1(new_n310), .B2(new_n578), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n407), .A2(new_n227), .A3(new_n408), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n579), .B(new_n584), .C1(new_n585), .C2(new_n324), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n261), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n353), .A2(new_n264), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n509), .A2(KEYINPUT84), .A3(new_n353), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT84), .ZN(new_n591));
  INV_X1    g0391(.A(new_n353), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n591), .B1(new_n508), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n587), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n207), .A2(G1698), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(G238), .B2(G1698), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n374), .A2(new_n378), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n285), .B1(new_n598), .B2(new_n494), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n295), .A2(G250), .A3(new_n465), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT82), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n295), .A2(KEYINPUT82), .A3(G250), .A4(new_n465), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n466), .A2(G274), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n599), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n348), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n595), .B(new_n607), .C1(G179), .C2(new_n606), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n508), .A2(new_n211), .ZN(new_n609));
  AOI211_X1 g0409(.A(new_n588), .B(new_n609), .C1(new_n586), .C2(new_n261), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n606), .A2(G200), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n599), .A2(new_n604), .A3(G190), .A4(new_n605), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n542), .A2(new_n543), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n284), .B1(new_n615), .B2(new_n572), .ZN(new_n616));
  INV_X1    g0416(.A(new_n567), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n565), .ZN(new_n618));
  OAI21_X1  g0418(.A(G200), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT81), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n619), .A2(new_n620), .A3(new_n562), .A4(new_n548), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n348), .B1(new_n616), .B2(new_n537), .ZN(new_n622));
  INV_X1    g0422(.A(new_n562), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n568), .A2(new_n575), .A3(new_n487), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n577), .A2(new_n614), .A3(new_n621), .A4(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n535), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n445), .A2(new_n627), .ZN(G372));
  AND3_X1   g0428(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT26), .B1(new_n629), .B2(new_n614), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n608), .A2(new_n613), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n625), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n608), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT90), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(KEYINPUT90), .B(new_n608), .C1(new_n630), .C2(new_n633), .ZN(new_n637));
  INV_X1    g0437(.A(new_n626), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n458), .A2(new_n485), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT21), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND4_X1   g0441(.A1(G179), .A2(new_n473), .A3(new_n479), .A4(new_n484), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n457), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n458), .A2(new_n485), .A3(KEYINPUT21), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT89), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT89), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n641), .A2(new_n643), .A3(new_n647), .A4(new_n644), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n527), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n638), .A2(new_n649), .A3(new_n532), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n636), .A2(new_n637), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n445), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n441), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n436), .A2(KEYINPUT18), .A3(new_n439), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n338), .A2(new_n369), .B1(new_n345), .B2(new_n344), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n433), .B(KEYINPUT17), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n655), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n351), .B1(new_n659), .B2(new_n306), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n652), .A2(new_n660), .ZN(G369));
  NAND4_X1  g0461(.A1(new_n534), .A2(new_n643), .A3(new_n641), .A4(new_n644), .ZN(new_n662));
  INV_X1    g0462(.A(G13), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G20), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n263), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G343), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n669), .B(KEYINPUT91), .Z(new_n670));
  AOI21_X1  g0470(.A(new_n662), .B1(new_n457), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n457), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n646), .B2(new_n648), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT92), .ZN(new_n675));
  XOR2_X1   g0475(.A(KEYINPUT93), .B(G330), .Z(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n532), .A2(new_n527), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n513), .A2(new_n670), .ZN(new_n680));
  INV_X1    g0480(.A(new_n670), .ZN(new_n681));
  OAI22_X1  g0481(.A1(new_n679), .A2(new_n680), .B1(new_n527), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n491), .A2(new_n527), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n684), .A2(new_n532), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n681), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT94), .ZN(G399));
  INV_X1    g0488(.A(new_n231), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n290), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G1), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n580), .A2(new_n208), .A3(new_n581), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n229), .A2(G50), .ZN(new_n694));
  OAI22_X1  g0494(.A1(new_n692), .A2(new_n693), .B1(new_n694), .B2(new_n691), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n634), .B1(new_n638), .B2(new_n685), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT29), .B1(new_n697), .B2(new_n670), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n651), .A2(new_n681), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(KEYINPUT29), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT97), .B1(new_n627), .B2(new_n681), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT97), .ZN(new_n702));
  NOR4_X1   g0502(.A1(new_n535), .A2(new_n626), .A3(new_n702), .A4(new_n670), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n481), .A2(new_n483), .A3(new_n482), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n483), .B1(new_n481), .B2(new_n482), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(G179), .B1(new_n706), .B2(new_n479), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n568), .A2(new_n575), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n707), .A2(new_n708), .A3(new_n606), .A4(new_n525), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT96), .ZN(new_n711));
  INV_X1    g0511(.A(new_n606), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n537), .B1(new_n574), .B2(new_n285), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n523), .A2(new_n524), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n518), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n642), .A2(new_n712), .A3(new_n713), .A4(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n711), .B1(new_n716), .B2(KEYINPUT95), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n710), .B1(new_n717), .B2(KEYINPUT30), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n706), .A2(new_n712), .A3(G179), .A4(new_n479), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n575), .A2(new_n715), .A3(new_n538), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT95), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT96), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n711), .B1(new_n719), .B2(new_n720), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT30), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  AOI211_X1 g0525(.A(KEYINPUT31), .B(new_n681), .C1(new_n718), .C2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n721), .A2(KEYINPUT96), .A3(KEYINPUT30), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n716), .B2(new_n711), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n728), .B(new_n709), .C1(new_n717), .C2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n727), .B1(new_n731), .B2(new_n670), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n701), .A2(new_n703), .B1(new_n726), .B2(new_n732), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n733), .A2(new_n676), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n700), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n696), .B1(new_n736), .B2(G1), .ZN(G364));
  AOI21_X1  g0537(.A(new_n263), .B1(new_n664), .B2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n690), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n678), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(new_n676), .B2(new_n675), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n528), .A2(G179), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n227), .A2(G190), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT100), .Z(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n360), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G179), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G159), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT32), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n743), .A2(G20), .A3(G190), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n748), .A2(G190), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n276), .B1(new_n753), .B2(new_n580), .C1(new_n756), .C2(new_n213), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n747), .A2(new_n752), .A3(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n227), .A2(new_n487), .A3(new_n528), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n423), .A2(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n227), .A2(new_n487), .A3(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n423), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G58), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n202), .A2(new_n760), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n761), .A2(new_n301), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT99), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT99), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n764), .B1(new_n768), .B2(G77), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n759), .A2(new_n301), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n758), .B(new_n769), .C1(new_n324), .C2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT101), .ZN(new_n772));
  INV_X1    g0572(.A(G303), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n753), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G294), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n756), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G317), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n777), .A2(KEYINPUT33), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(KEYINPUT33), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n770), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n760), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n776), .B(new_n780), .C1(G326), .C2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n746), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G283), .ZN(new_n784));
  INV_X1    g0584(.A(new_n762), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n785), .A2(G322), .B1(G311), .B2(new_n765), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n276), .B1(new_n750), .B2(G329), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n782), .A2(new_n784), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n772), .B1(new_n774), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n226), .B1(G20), .B2(new_n348), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n247), .A2(G45), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n407), .A2(new_n408), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n689), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n794), .B(new_n797), .C1(G45), .C2(new_n694), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n276), .A2(G355), .A3(new_n231), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(G116), .C2(new_n231), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n793), .B(new_n790), .C1(new_n800), .C2(KEYINPUT98), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(KEYINPUT98), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n789), .A2(new_n790), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n793), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n740), .B(new_n803), .C1(new_n675), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n742), .A2(new_n805), .ZN(G396));
  AND2_X1   g0606(.A1(new_n670), .A2(new_n358), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n370), .B1(new_n444), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n369), .A2(new_n681), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n699), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n651), .A2(new_n681), .A3(new_n810), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(new_n734), .ZN(new_n815));
  INV_X1    g0615(.A(new_n740), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G137), .A2(new_n781), .B1(new_n785), .B2(G143), .ZN(new_n818));
  INV_X1    g0618(.A(G150), .ZN(new_n819));
  INV_X1    g0619(.A(new_n768), .ZN(new_n820));
  INV_X1    g0620(.A(G159), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n818), .B1(new_n819), .B2(new_n770), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT34), .ZN(new_n823));
  INV_X1    g0623(.A(G132), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n796), .B1(new_n763), .B2(new_n756), .C1(new_n824), .C2(new_n749), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G68), .B2(new_n783), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n823), .B(new_n826), .C1(new_n202), .C2(new_n753), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n760), .A2(new_n773), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n770), .A2(KEYINPUT102), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n770), .A2(KEYINPUT102), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G116), .A2(new_n768), .B1(new_n832), .B2(G283), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n746), .A2(new_n211), .ZN(new_n834));
  INV_X1    g0634(.A(new_n753), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n834), .B1(G107), .B2(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n785), .A2(G294), .B1(G97), .B2(new_n755), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n276), .B1(new_n750), .B2(G311), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n833), .A2(new_n836), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n827), .B1(new_n828), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n790), .A2(new_n791), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n840), .A2(new_n790), .B1(new_n206), .B2(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n842), .B(new_n740), .C1(new_n792), .C2(new_n810), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n817), .A2(new_n843), .ZN(G384));
  INV_X1    g0644(.A(KEYINPUT104), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n436), .B1(new_n439), .B2(new_n668), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT37), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n846), .A2(new_n847), .A3(new_n433), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n395), .A2(new_n261), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT16), .B1(new_n383), .B2(new_n394), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n429), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n852), .A2(new_n853), .B1(new_n439), .B2(new_n668), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n847), .B1(new_n854), .B2(new_n433), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n845), .B1(new_n849), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n668), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n383), .A2(new_n394), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n396), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n859), .A2(new_n261), .A3(new_n395), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n857), .B1(new_n860), .B2(new_n429), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n442), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(G169), .B1(new_n431), .B2(new_n413), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n863), .A2(new_n438), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n864), .A2(new_n857), .B1(new_n860), .B2(new_n429), .ZN(new_n865));
  INV_X1    g0665(.A(new_n433), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT37), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(KEYINPUT104), .A3(new_n848), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n856), .A2(new_n862), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n856), .A2(new_n862), .A3(new_n868), .A4(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT105), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n338), .A2(new_n346), .A3(KEYINPUT103), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n681), .A2(new_n329), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n344), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n338), .A2(new_n880), .A3(KEYINPUT103), .A4(new_n877), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n879), .A2(new_n810), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n679), .A2(new_n662), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n638), .A2(new_n883), .A3(new_n681), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n702), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n627), .A2(KEYINPUT97), .A3(new_n681), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n732), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n731), .A2(new_n727), .A3(new_n670), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n882), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n871), .A2(KEYINPUT105), .A3(new_n872), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n875), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT40), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n436), .A2(new_n668), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n655), .B2(new_n657), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n847), .B1(new_n846), .B2(new_n433), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n849), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n870), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n894), .B1(new_n872), .B2(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n893), .A2(new_n894), .B1(new_n891), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n445), .A2(new_n733), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n901), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n676), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n879), .A2(new_n881), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n813), .B2(new_n809), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(new_n875), .A3(new_n892), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n653), .A2(new_n654), .A3(new_n857), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n346), .A2(new_n670), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n871), .B2(new_n872), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n872), .A2(new_n899), .A3(new_n910), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n907), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n700), .A2(new_n445), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n660), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n914), .B(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n904), .B(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n263), .B2(new_n664), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n208), .B1(new_n556), .B2(KEYINPUT35), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n920), .B(new_n228), .C1(KEYINPUT35), .C2(new_n556), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT36), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n384), .A2(G77), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n694), .A2(new_n923), .B1(G50), .B2(new_n324), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(G1), .A3(new_n663), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n919), .A2(new_n922), .A3(new_n925), .ZN(G367));
  AND3_X1   g0726(.A1(new_n577), .A2(new_n625), .A3(new_n621), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n562), .B2(new_n681), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n629), .A2(new_n670), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n679), .A2(new_n491), .A3(new_n670), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT42), .Z(new_n933));
  INV_X1    g0733(.A(KEYINPUT106), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n625), .B1(new_n928), .B2(new_n527), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n681), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n934), .B1(new_n933), .B2(new_n936), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n681), .A2(new_n610), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(new_n631), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n938), .A2(new_n939), .B1(KEYINPUT43), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n939), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n941), .B(KEYINPUT43), .Z(new_n945));
  NAND3_X1  g0745(.A1(new_n944), .A2(new_n937), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n678), .A2(new_n682), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n930), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT107), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n949), .A2(new_n950), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n931), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n491), .A2(new_n670), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n955), .B1(new_n682), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n677), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT108), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n677), .A2(new_n957), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(KEYINPUT108), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(new_n735), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n930), .A2(new_n686), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT45), .Z(new_n965));
  NOR2_X1   g0765(.A1(new_n686), .A2(new_n927), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT44), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n948), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n683), .A2(new_n965), .A3(new_n967), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n963), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n736), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n690), .B(KEYINPUT41), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n954), .B1(new_n975), .B2(new_n739), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G283), .A2(new_n768), .B1(new_n832), .B2(G294), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n750), .A2(G317), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n753), .A2(new_n208), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT46), .ZN(new_n980));
  INV_X1    g0780(.A(G311), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n980), .B1(new_n981), .B2(new_n760), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G303), .B2(new_n785), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n979), .A2(KEYINPUT46), .B1(new_n756), .B2(new_n360), .ZN(new_n984));
  INV_X1    g0784(.A(new_n745), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n796), .B(new_n984), .C1(G97), .C2(new_n985), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n977), .A2(new_n978), .A3(new_n983), .A4(new_n986), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G50), .A2(new_n768), .B1(new_n832), .B2(G159), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n276), .B1(new_n745), .B2(new_n206), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT110), .Z(new_n990));
  NOR2_X1   g0790(.A1(new_n756), .A2(new_n324), .ZN(new_n991));
  INV_X1    g0791(.A(G137), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n762), .A2(new_n819), .B1(new_n992), .B2(new_n749), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n991), .B(new_n993), .C1(G143), .C2(new_n781), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n988), .A2(new_n990), .A3(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n753), .A2(new_n763), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n987), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n998));
  XNOR2_X1  g0798(.A(new_n997), .B(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n816), .B1(new_n999), .B2(new_n790), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n793), .A2(new_n790), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n797), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1001), .B1(new_n231), .B2(new_n592), .C1(new_n243), .C2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT109), .Z(new_n1004));
  OAI211_X1 g0804(.A(new_n1000), .B(new_n1004), .C1(new_n942), .C2(new_n804), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n976), .A2(new_n1005), .ZN(G387));
  OR2_X1    g0806(.A1(new_n962), .A2(new_n735), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n962), .A2(new_n735), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n690), .A3(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n768), .A2(G303), .B1(G322), .B2(new_n781), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n981), .B2(new_n831), .C1(new_n777), .C2(new_n762), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT48), .ZN(new_n1012));
  INV_X1    g0812(.A(G283), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1012), .B1(new_n1013), .B2(new_n756), .C1(new_n775), .C2(new_n753), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT49), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n750), .A2(G326), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n796), .B1(G116), .B2(new_n985), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n756), .A2(new_n592), .B1(new_n770), .B2(new_n258), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n795), .B(new_n1021), .C1(G159), .C2(new_n781), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n835), .A2(G77), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n783), .A2(G97), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n765), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1025), .A2(new_n324), .B1(new_n762), .B2(new_n202), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(KEYINPUT114), .B(G150), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1026), .B1(new_n750), .B2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1020), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n693), .A2(new_n231), .A3(new_n276), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n258), .A2(G50), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT50), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n316), .C1(new_n324), .C2(new_n206), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n797), .B1(new_n1034), .B2(new_n693), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT113), .Z(new_n1036));
  NOR2_X1   g0836(.A1(new_n240), .A2(new_n316), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1031), .B1(G107), .B2(new_n231), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1030), .A2(new_n790), .B1(new_n1001), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1039), .B(new_n740), .C1(new_n682), .C2(new_n804), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT115), .Z(new_n1041));
  NAND4_X1  g0841(.A1(new_n959), .A2(new_n739), .A3(new_n960), .A4(new_n961), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT112), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1009), .A2(new_n1041), .A3(new_n1044), .ZN(G393));
  NAND2_X1  g0845(.A1(new_n971), .A2(new_n739), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1001), .B1(new_n213), .B2(new_n231), .C1(new_n250), .C2(new_n1002), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n750), .A2(G143), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n796), .B(new_n1048), .C1(new_n324), .C2(new_n753), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1049), .B(new_n834), .C1(G77), .C2(new_n755), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n832), .A2(G50), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n819), .A2(new_n760), .B1(new_n762), .B2(new_n821), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT51), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n768), .A2(new_n425), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n765), .A2(G294), .B1(G116), .B2(new_n755), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1056), .B(new_n362), .C1(new_n1013), .C2(new_n753), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n747), .B(new_n1057), .C1(G322), .C2(new_n750), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n773), .B2(new_n831), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n981), .A2(new_n762), .B1(new_n760), .B2(new_n777), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT52), .Z(new_n1061));
  OAI21_X1  g0861(.A(new_n1055), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n816), .B1(new_n1062), .B2(new_n790), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1047), .B(new_n1063), .C1(new_n930), .C2(new_n804), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1046), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT116), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1046), .A2(KEYINPUT116), .A3(new_n1064), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n971), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1007), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1071), .A2(new_n690), .A3(new_n972), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1069), .A2(new_n1072), .ZN(G390));
  NOR2_X1   g0873(.A1(new_n911), .A2(new_n912), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n906), .B2(new_n909), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n909), .B1(new_n872), .B2(new_n899), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n685), .A2(new_n638), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n634), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n670), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1079), .A2(new_n808), .B1(new_n369), .B2(new_n681), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1076), .B1(new_n1080), .B2(new_n905), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1075), .A2(new_n1081), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n879), .A2(new_n810), .A3(new_n881), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n733), .A2(G330), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(KEYINPUT117), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT117), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n733), .A2(new_n1083), .A3(new_n1086), .A4(G330), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1082), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n733), .A2(new_n676), .A3(new_n810), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1091), .A2(new_n905), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1075), .A2(new_n1081), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n445), .A2(G330), .A3(new_n733), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n915), .A2(new_n660), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1091), .A2(new_n905), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1085), .A2(new_n1097), .A3(new_n1087), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n813), .A2(new_n809), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n905), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n734), .A2(new_n810), .A3(new_n1101), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n733), .A2(G330), .A3(new_n810), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1102), .B(new_n1080), .C1(new_n1101), .C2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1096), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT118), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1094), .A2(new_n1106), .A3(new_n1105), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(new_n1094), .B2(new_n1105), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n690), .B1(new_n1094), .B2(new_n1105), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1074), .A2(new_n791), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n783), .A2(G68), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n785), .A2(G116), .B1(G77), .B2(new_n755), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n276), .B1(new_n835), .B2(G87), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n750), .A2(G294), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n820), .A2(new_n213), .B1(new_n360), .B2(new_n831), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1115), .B(new_n1116), .C1(G283), .C2(new_n781), .ZN(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT54), .B(G143), .Z(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n820), .A2(new_n1119), .B1(new_n992), .B2(new_n831), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n835), .A2(new_n1027), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT53), .Z(new_n1122));
  INV_X1    g0922(.A(G125), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1122), .B(new_n276), .C1(new_n1123), .C2(new_n749), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n745), .A2(new_n202), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G128), .A2(new_n781), .B1(new_n785), .B2(G132), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n821), .B2(new_n756), .ZN(new_n1127));
  NOR4_X1   g0927(.A1(new_n1120), .A2(new_n1124), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n790), .B1(new_n1117), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n841), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n740), .B1(new_n425), .B2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT119), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1110), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT120), .Z(new_n1134));
  NAND2_X1  g0934(.A1(new_n1094), .A2(new_n739), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1109), .A2(new_n1134), .A3(new_n1135), .ZN(G378));
  INV_X1    g0936(.A(KEYINPUT57), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1096), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1075), .A2(new_n1081), .A3(new_n1092), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1088), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(KEYINPUT118), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1094), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1096), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n306), .A2(new_n352), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n272), .A2(new_n857), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1147), .B(new_n1148), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1149), .A2(KEYINPUT55), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(KEYINPUT55), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1150), .A2(KEYINPUT56), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT56), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n893), .A2(new_n894), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n891), .A2(new_n900), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(G330), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n914), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n907), .A2(new_n908), .A3(new_n913), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n901), .A3(G330), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1154), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1154), .B1(new_n1160), .B2(new_n1158), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1137), .B1(new_n1146), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1139), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1154), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1161), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1166), .A2(KEYINPUT57), .A3(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1165), .A2(new_n690), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1154), .A2(new_n791), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n841), .A2(new_n202), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n756), .A2(new_n324), .B1(new_n1013), .B2(new_n749), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G107), .A2(new_n785), .B1(new_n781), .B2(G116), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n213), .B2(new_n770), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(G58), .C2(new_n985), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1023), .A2(new_n795), .A3(new_n315), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT121), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(new_n592), .C2(new_n1025), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT58), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1025), .A2(new_n992), .B1(new_n824), .B2(new_n770), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT122), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n756), .A2(new_n819), .B1(new_n1119), .B2(new_n753), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G128), .B2(new_n785), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(new_n1123), .C2(new_n760), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(G33), .A2(G41), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n985), .A2(G159), .B1(new_n750), .B2(G124), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n202), .B1(G33), .B2(G41), .C1(new_n796), .C2(new_n290), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1182), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n816), .B1(new_n1194), .B2(new_n790), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1173), .A2(new_n1174), .A3(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(KEYINPUT123), .B(new_n1196), .C1(new_n1164), .C2(new_n738), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT123), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n738), .B1(new_n1169), .B2(new_n1161), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1196), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1197), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1172), .A2(new_n1202), .ZN(G375));
  NAND3_X1  g1003(.A1(new_n1100), .A2(new_n1104), .A3(new_n1096), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1140), .A2(new_n974), .A3(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT124), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n832), .A2(new_n1118), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n824), .A2(new_n760), .B1(new_n762), .B2(new_n992), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G150), .B2(new_n765), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n750), .A2(G128), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n753), .A2(new_n821), .B1(new_n745), .B2(new_n763), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n795), .B(new_n1211), .C1(G50), .C2(new_n755), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1207), .A2(new_n1209), .A3(new_n1210), .A4(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G107), .A2(new_n768), .B1(new_n832), .B2(G116), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n756), .A2(new_n592), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n760), .A2(new_n775), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(G283), .C2(new_n785), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n362), .B1(new_n749), .B2(new_n773), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n783), .B2(G77), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1214), .A2(new_n1217), .A3(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n753), .A2(new_n213), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1213), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n790), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(G68), .B2(new_n1130), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n816), .B(new_n1224), .C1(new_n905), .C2(new_n791), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1138), .B2(new_n739), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1206), .A2(new_n1226), .ZN(G381));
  XNOR2_X1  g1027(.A(G375), .B(KEYINPUT125), .ZN(new_n1228));
  INV_X1    g1028(.A(G378), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(new_n1226), .A4(new_n1206), .ZN(new_n1230));
  INV_X1    g1030(.A(G396), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1009), .A2(new_n1041), .A3(new_n1044), .A4(new_n1231), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(G387), .A2(G384), .A3(G390), .A4(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1230), .A2(new_n1234), .ZN(G407));
  INV_X1    g1035(.A(G343), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1228), .A2(new_n1236), .A3(new_n1229), .ZN(new_n1237));
  OAI211_X1 g1037(.A(G213), .B(new_n1237), .C1(new_n1230), .C2(new_n1234), .ZN(G409));
  AND2_X1   g1038(.A1(new_n1236), .A2(G213), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1172), .A2(G378), .A3(new_n1202), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1166), .A2(new_n974), .A3(new_n1170), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1229), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1239), .B1(new_n1240), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT60), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1204), .A2(new_n1246), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1100), .A2(new_n1104), .A3(KEYINPUT60), .A4(new_n1096), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1247), .A2(new_n1140), .A3(new_n690), .A4(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(G384), .A3(new_n1226), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT126), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1226), .ZN(new_n1252));
  INV_X1    g1052(.A(G384), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT126), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1249), .A2(new_n1255), .A3(G384), .A4(new_n1226), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1251), .A2(new_n1254), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1239), .A2(G2897), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(KEYINPUT127), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(KEYINPUT127), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1259), .A2(KEYINPUT127), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1261), .B1(new_n1257), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(KEYINPUT63), .B1(new_n1245), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1245), .A2(new_n1258), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(G393), .A2(G396), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1232), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(G390), .A2(new_n1268), .A3(new_n1232), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(G387), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1271), .A2(new_n976), .A3(new_n1005), .A4(new_n1272), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1239), .B(new_n1257), .C1(new_n1240), .C2(new_n1244), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1276), .B1(new_n1277), .B2(KEYINPUT63), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1267), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT62), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1245), .A2(new_n1281), .A3(new_n1258), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1279), .B1(new_n1245), .B2(new_n1264), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1245), .B2(new_n1258), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1276), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1280), .B1(new_n1285), .B2(new_n1286), .ZN(G405));
  NAND2_X1  g1087(.A1(G375), .A2(new_n1229), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1240), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1258), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1288), .A2(new_n1240), .A3(new_n1257), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(new_n1276), .ZN(G402));
endmodule


