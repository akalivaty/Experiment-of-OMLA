//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT6), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT70), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G119), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT70), .A3(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(G119), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n194), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT69), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n200));
  INV_X1    g014(.A(G113), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT69), .B1(KEYINPUT2), .B2(G113), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n202), .A2(new_n203), .B1(KEYINPUT2), .B2(G113), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT5), .A4(new_n197), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n193), .A2(KEYINPUT5), .A3(G119), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(new_n201), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n198), .A2(new_n204), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT3), .B1(new_n209), .B2(G107), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G104), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n209), .A2(G107), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n210), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n209), .A2(G107), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n212), .A2(G104), .ZN(new_n218));
  OAI21_X1  g032(.A(G101), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n208), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n210), .A2(new_n213), .A3(new_n215), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(G101), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT81), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n223), .A2(KEYINPUT81), .A3(new_n224), .A4(G101), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n202), .A2(new_n203), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT2), .A2(G113), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n194), .A2(new_n196), .A3(new_n197), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n198), .A2(new_n204), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n224), .B1(new_n223), .B2(G101), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n216), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n222), .B1(new_n229), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  XOR2_X1   g055(.A(new_n241), .B(KEYINPUT84), .Z(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n191), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n222), .B(new_n242), .C1(new_n229), .C2(new_n239), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(KEYINPUT85), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT85), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n234), .A2(new_n235), .B1(new_n237), .B2(new_n216), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n227), .A2(new_n228), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n248), .A2(new_n249), .B1(new_n221), .B2(new_n208), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n247), .B1(new_n250), .B2(new_n242), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n244), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT86), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(G146), .ZN(new_n255));
  INV_X1    g069(.A(G146), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(G143), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  OAI22_X1  g073(.A1(new_n255), .A2(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(G143), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n254), .A2(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n260), .A2(G125), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n261), .A2(new_n262), .ZN(new_n266));
  INV_X1    g080(.A(G128), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n266), .A2(new_n267), .B1(KEYINPUT1), .B2(new_n257), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n269));
  XNOR2_X1  g083(.A(G143), .B(G146), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n267), .A2(KEYINPUT1), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AND4_X1   g086(.A1(new_n269), .A2(new_n271), .A3(new_n261), .A4(new_n262), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n268), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n265), .B1(new_n274), .B2(G125), .ZN(new_n275));
  INV_X1    g089(.A(G224), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G953), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n265), .B(new_n277), .C1(new_n274), .C2(G125), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n250), .A2(KEYINPUT6), .A3(new_n242), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n252), .A2(new_n253), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n242), .B(KEYINPUT8), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n221), .A2(new_n235), .ZN(new_n286));
  OR2_X1    g100(.A1(new_n205), .A2(KEYINPUT87), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n201), .B(new_n206), .C1(new_n205), .C2(KEYINPUT87), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n208), .A2(new_n221), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n285), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT7), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n275), .A2(new_n292), .A3(new_n278), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n278), .A2(new_n292), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n279), .A2(new_n280), .A3(new_n294), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n291), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n245), .A2(KEYINPUT85), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n250), .A2(new_n247), .A3(new_n242), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n284), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n282), .B1(new_n299), .B2(new_n244), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n253), .B1(new_n302), .B2(new_n281), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n190), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n252), .A2(new_n281), .A3(new_n283), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT86), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n306), .A2(new_n189), .A3(new_n284), .A4(new_n300), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n188), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT66), .B(G131), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(G237), .A2(G953), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(G143), .A3(G214), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(G143), .B1(new_n311), .B2(G214), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n310), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT88), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n310), .B(KEYINPUT88), .C1(new_n313), .C2(new_n314), .ZN(new_n318));
  INV_X1    g132(.A(G237), .ZN(new_n319));
  INV_X1    g133(.A(G953), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(G214), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n254), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(new_n309), .A3(new_n312), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n317), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G125), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G140), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n328), .A3(KEYINPUT16), .ZN(new_n329));
  OR3_X1    g143(.A1(new_n327), .A2(KEYINPUT16), .A3(G140), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n329), .A2(G146), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G125), .B(G140), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT19), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n331), .B1(new_n333), .B2(new_n256), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n324), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n322), .A2(new_n312), .ZN(new_n336));
  NAND2_X1  g150(.A1(KEYINPUT18), .A2(G131), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n336), .B(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n332), .A2(new_n256), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n332), .A2(KEYINPUT78), .A3(new_n256), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n332), .A2(new_n256), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n338), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n335), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G113), .B(G122), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT89), .B(G104), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n318), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT88), .B1(new_n336), .B2(new_n310), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT17), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT17), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n317), .A2(new_n354), .A3(new_n318), .A4(new_n323), .ZN(new_n355));
  AOI21_X1  g169(.A(G146), .B1(new_n329), .B2(new_n330), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n331), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n353), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n349), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n345), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n350), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(G475), .A2(G902), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(KEYINPUT90), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT20), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n361), .B(new_n362), .C1(KEYINPUT90), .C2(KEYINPUT20), .ZN(new_n367));
  INV_X1    g181(.A(G902), .ZN(new_n368));
  INV_X1    g182(.A(new_n360), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n359), .B1(new_n358), .B2(new_n345), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G475), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n367), .A3(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(KEYINPUT74), .B(G217), .Z(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT9), .B(G234), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n374), .A2(G953), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n193), .A2(G122), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n193), .A2(G122), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(new_n212), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n267), .A2(G143), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT92), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n383), .B1(new_n254), .B2(G128), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n267), .A2(KEYINPUT92), .A3(G143), .ZN(new_n385));
  AOI211_X1 g199(.A(G134), .B(new_n382), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G134), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n385), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n254), .A2(G128), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n381), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n380), .A2(KEYINPUT14), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT94), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT94), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT14), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n193), .B2(G122), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n394), .B1(new_n396), .B2(new_n380), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n393), .B1(new_n397), .B2(new_n392), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n391), .B1(G107), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n380), .ZN(new_n400));
  OAI21_X1  g214(.A(G107), .B1(new_n400), .B2(new_n378), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n381), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n388), .A2(new_n387), .A3(new_n389), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OR2_X1    g218(.A1(KEYINPUT91), .A2(KEYINPUT13), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT91), .A2(KEYINPUT13), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n389), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n388), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT93), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n388), .A2(new_n407), .A3(KEYINPUT93), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n405), .A2(new_n406), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n382), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n404), .B1(new_n414), .B2(G134), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n377), .B1(new_n399), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n398), .A2(G107), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n417), .B(new_n381), .C1(new_n386), .C2(new_n390), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n411), .A2(new_n413), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n387), .B1(new_n419), .B2(new_n410), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n418), .B(new_n376), .C1(new_n420), .C2(new_n404), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n368), .ZN(new_n423));
  INV_X1    g237(.A(G478), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(KEYINPUT15), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n422), .B(new_n368), .C1(KEYINPUT15), .C2(new_n424), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(G234), .A2(G237), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(G952), .A3(new_n320), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(G902), .A3(G953), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(G898), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n373), .A2(new_n428), .A3(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n308), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n311), .A2(G210), .ZN(new_n438));
  XOR2_X1   g252(.A(new_n438), .B(KEYINPUT27), .Z(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT71), .ZN(new_n440));
  XOR2_X1   g254(.A(KEYINPUT26), .B(G101), .Z(new_n441));
  XOR2_X1   g255(.A(new_n440), .B(new_n441), .Z(new_n442));
  INV_X1    g256(.A(KEYINPUT28), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT11), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n387), .B2(G137), .ZN(new_n445));
  INV_X1    g259(.A(G137), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT11), .A3(G134), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n387), .A2(G137), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n445), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(G134), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n448), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n449), .A2(new_n309), .B1(G131), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n274), .A2(KEYINPUT68), .A3(new_n452), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n309), .A2(new_n447), .A3(new_n448), .A4(new_n445), .ZN(new_n454));
  INV_X1    g268(.A(G131), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n449), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n259), .A2(new_n258), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n264), .B(KEYINPUT65), .C1(new_n457), .C2(new_n270), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT65), .B1(new_n260), .B2(new_n264), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT68), .B1(new_n274), .B2(new_n452), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n236), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n236), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n274), .A2(new_n452), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n260), .A2(new_n264), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n456), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n443), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n469), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(KEYINPUT28), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n442), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT68), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n254), .A2(KEYINPUT1), .A3(G146), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n475), .B1(new_n270), .B2(G128), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n271), .A2(new_n261), .A3(new_n262), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT67), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n270), .A2(new_n269), .A3(new_n271), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n451), .A2(G131), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n454), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n474), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n461), .A3(new_n453), .ZN(new_n484));
  XOR2_X1   g298(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n466), .A2(new_n468), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT30), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n236), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT31), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n440), .B(new_n441), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n469), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n473), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n489), .A2(new_n469), .A3(new_n491), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT31), .ZN(new_n495));
  AOI21_X1  g309(.A(G902), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT73), .ZN(new_n497));
  INV_X1    g311(.A(G472), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT32), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n495), .A2(new_n492), .A3(new_n473), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n500), .A2(KEYINPUT32), .A3(new_n498), .A4(new_n368), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT73), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n473), .A2(new_n492), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n484), .A2(new_n485), .B1(new_n487), .B2(KEYINPUT30), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n471), .B1(new_n504), .B2(new_n236), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n490), .B1(new_n505), .B2(new_n491), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n498), .B(new_n368), .C1(new_n503), .C2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT32), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n465), .B1(new_n466), .B2(new_n468), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n469), .B1(new_n510), .B2(KEYINPUT72), .ZN(new_n511));
  OR2_X1    g325(.A1(new_n469), .A2(KEYINPUT72), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n443), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(new_n472), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT29), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n442), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(G902), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n472), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n471), .B1(new_n236), .B2(new_n484), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n518), .B(new_n491), .C1(new_n519), .C2(new_n443), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n520), .B(new_n515), .C1(new_n505), .C2(new_n491), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G472), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n499), .A2(new_n502), .A3(new_n509), .A4(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT75), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(new_n195), .B2(G128), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n195), .A2(G128), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n267), .A2(KEYINPUT75), .A3(G119), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT24), .B(G110), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n331), .B2(new_n356), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT23), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n195), .B2(G128), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n267), .A2(KEYINPUT23), .A3(G119), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(new_n527), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G110), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT76), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(KEYINPUT76), .A3(G110), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n532), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n529), .A2(new_n530), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(G110), .B2(new_n536), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT77), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n331), .B1(new_n341), .B2(new_n342), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT77), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n543), .B(new_n547), .C1(G110), .C2(new_n536), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT22), .B(G137), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n320), .A2(G221), .A3(G234), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n551), .B(new_n552), .Z(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n542), .A2(new_n549), .A3(new_n553), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n374), .B1(G234), .B2(new_n368), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(G902), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT25), .ZN(new_n561));
  INV_X1    g375(.A(new_n556), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n553), .B1(new_n542), .B2(new_n549), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n561), .B(new_n368), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n558), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n561), .B1(new_n557), .B2(new_n368), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n560), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT79), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G469), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n274), .A2(new_n221), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n478), .A2(new_n479), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n220), .B1(new_n572), .B2(new_n268), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n456), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT12), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g390(.A(KEYINPUT12), .B(new_n456), .C1(new_n571), .C2(new_n573), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n237), .A2(new_n216), .B1(new_n260), .B2(new_n264), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n249), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n480), .B2(new_n220), .ZN(new_n582));
  INV_X1    g396(.A(new_n456), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n274), .A2(KEYINPUT10), .A3(new_n221), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n580), .A2(new_n582), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(G110), .B(G140), .ZN(new_n587));
  INV_X1    g401(.A(G227), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(G953), .ZN(new_n589));
  XOR2_X1   g403(.A(new_n587), .B(new_n589), .Z(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n480), .A2(new_n581), .A3(new_n220), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT10), .B1(new_n274), .B2(new_n221), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n583), .B1(new_n595), .B2(new_n580), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n585), .A2(new_n590), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n570), .B1(new_n599), .B2(new_n368), .ZN(new_n600));
  INV_X1    g414(.A(new_n585), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n591), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT82), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n585), .A2(new_n603), .A3(new_n590), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n578), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n603), .B1(new_n585), .B2(new_n590), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(new_n570), .A3(new_n368), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT83), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n597), .A2(KEYINPUT82), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n604), .A3(new_n578), .ZN(new_n611));
  AOI21_X1  g425(.A(G902), .B1(new_n611), .B2(new_n602), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT83), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n613), .A3(new_n570), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n600), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(G221), .B1(new_n375), .B2(G902), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT80), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n437), .A2(new_n524), .A3(new_n569), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  INV_X1    g434(.A(new_n308), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n435), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT95), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n496), .B1(new_n623), .B2(new_n498), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n368), .B1(new_n503), .B2(new_n506), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(KEYINPUT95), .A3(G472), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n569), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n423), .A2(G478), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n416), .A2(new_n421), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n629), .B1(new_n416), .B2(new_n421), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n368), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n628), .B1(new_n632), .B2(G478), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n366), .A2(new_n367), .A3(new_n372), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND4_X1   g450(.A1(new_n618), .A2(new_n622), .A3(new_n627), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT34), .B(G104), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  AOI21_X1  g453(.A(KEYINPUT20), .B1(new_n361), .B2(new_n362), .ZN(new_n640));
  INV_X1    g454(.A(new_n362), .ZN(new_n641));
  AOI211_X1 g455(.A(new_n365), .B(new_n641), .C1(new_n350), .C2(new_n360), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n643), .A2(new_n372), .A3(new_n428), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n621), .A2(new_n435), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n618), .A3(new_n627), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT96), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT35), .B(G107), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  AND2_X1   g463(.A1(new_n624), .A2(new_n626), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n553), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n550), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n559), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n653), .B1(new_n565), .B2(new_n566), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n437), .A2(new_n618), .A3(new_n650), .A4(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  INV_X1    g471(.A(new_n654), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n615), .A2(new_n617), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n433), .A2(new_n660), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n661), .A2(KEYINPUT97), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(KEYINPUT97), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n430), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n643), .A2(new_n428), .A3(new_n372), .A4(new_n664), .ZN(new_n665));
  AOI211_X1 g479(.A(new_n188), .B(new_n665), .C1(new_n304), .C2(new_n307), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n524), .A2(new_n659), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  XNOR2_X1  g482(.A(new_n664), .B(KEYINPUT39), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n618), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT40), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n511), .A2(new_n512), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n494), .B1(new_n491), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n498), .B1(new_n673), .B2(new_n368), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n507), .B2(new_n508), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n499), .A2(new_n502), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n304), .A2(new_n307), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT38), .Z(new_n679));
  INV_X1    g493(.A(new_n428), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n635), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n658), .A3(new_n187), .ZN(new_n682));
  OR4_X1    g496(.A1(new_n671), .A2(new_n677), .A3(new_n679), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  AND3_X1   g498(.A1(new_n373), .A2(new_n633), .A3(new_n664), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n308), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n524), .A3(new_n659), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT98), .B(G146), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G48));
  AND2_X1   g503(.A1(new_n524), .A2(new_n569), .ZN(new_n690));
  INV_X1    g504(.A(new_n617), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n612), .A2(new_n570), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n613), .B1(new_n612), .B2(new_n570), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n613), .A2(new_n607), .A3(new_n570), .A4(new_n368), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n691), .B(new_n692), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT99), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n612), .A2(new_n570), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n609), .B2(new_n614), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT99), .B1(new_n699), .B2(new_n691), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n690), .A2(new_n636), .A3(new_n701), .A4(new_n622), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT41), .B(G113), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  NAND3_X1  g518(.A1(new_n690), .A2(new_n645), .A3(new_n701), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  NOR3_X1   g520(.A1(new_n697), .A2(new_n700), .A3(new_n621), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n524), .A2(new_n436), .A3(new_n654), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT100), .B(G119), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G21));
  OAI21_X1  g525(.A(new_n442), .B1(new_n513), .B2(new_n472), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n495), .A2(new_n712), .A3(new_n492), .ZN(new_n713));
  NOR2_X1   g527(.A1(G472), .A2(G902), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n625), .A2(G472), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n435), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n567), .A2(KEYINPUT101), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT101), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n718), .B(new_n560), .C1(new_n565), .C2(new_n566), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n715), .A2(new_n716), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n695), .A2(new_n696), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n699), .A2(KEYINPUT99), .A3(new_n691), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n678), .A2(new_n187), .A3(new_n681), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT102), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT102), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n308), .A2(new_n727), .A3(new_n681), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  AND3_X1   g545(.A1(new_n715), .A2(new_n654), .A3(new_n685), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n701), .A2(KEYINPUT103), .A3(new_n308), .A4(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n722), .A3(new_n308), .A4(new_n723), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT103), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  INV_X1    g552(.A(new_n509), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n523), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n496), .A2(KEYINPUT106), .A3(KEYINPUT32), .A4(new_n498), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n501), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n507), .A2(new_n740), .A3(new_n508), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n742), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n720), .B1(new_n741), .B2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n304), .A2(new_n307), .A3(new_n691), .A4(new_n187), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n609), .A2(new_n614), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n592), .A2(G469), .A3(new_n598), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n570), .A2(new_n368), .ZN(new_n753));
  XOR2_X1   g567(.A(new_n753), .B(KEYINPUT104), .Z(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n750), .B1(new_n751), .B2(new_n756), .ZN(new_n757));
  AOI211_X1 g571(.A(KEYINPUT105), .B(new_n755), .C1(new_n609), .C2(new_n614), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n685), .B(new_n749), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT42), .B1(new_n747), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n756), .B1(new_n693), .B2(new_n694), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT105), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n751), .A2(new_n750), .A3(new_n756), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n748), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n685), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(KEYINPUT42), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n690), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n760), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G131), .ZN(G33));
  INV_X1    g583(.A(new_n665), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n764), .A2(new_n524), .A3(new_n569), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT108), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n690), .A2(new_n773), .A3(new_n770), .A4(new_n764), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  XNOR2_X1  g590(.A(new_n599), .B(KEYINPUT45), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(G469), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT109), .ZN(new_n779));
  INV_X1    g593(.A(new_n754), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(KEYINPUT46), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(KEYINPUT46), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n751), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n691), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n669), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n678), .A2(new_n188), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n634), .A2(new_n373), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT43), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n792), .A2(new_n650), .A3(new_n658), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n789), .B1(new_n793), .B2(KEYINPUT44), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(KEYINPUT44), .B2(new_n793), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n787), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(new_n446), .ZN(G39));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT47), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n798), .B1(new_n786), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n785), .A2(KEYINPUT111), .A3(KEYINPUT47), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n786), .B2(new_n799), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n785), .A2(KEYINPUT110), .A3(KEYINPUT47), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n800), .B(new_n801), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  OR4_X1    g619(.A1(new_n524), .A2(new_n789), .A3(new_n765), .A4(new_n569), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(KEYINPUT112), .B(G140), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(G42));
  XNOR2_X1  g623(.A(new_n699), .B(KEYINPUT49), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n691), .A2(new_n790), .A3(new_n720), .A4(new_n187), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n679), .A2(new_n677), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n715), .A2(new_n720), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n792), .A2(new_n430), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n788), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n699), .A2(new_n617), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n816), .B1(new_n805), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n815), .A2(new_n188), .A3(new_n679), .ZN(new_n820));
  INV_X1    g634(.A(new_n701), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n820), .A2(new_n819), .A3(new_n821), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n825), .A2(KEYINPUT117), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(KEYINPUT117), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n701), .A2(new_n431), .A3(new_n788), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n792), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n654), .A3(new_n715), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n677), .A2(new_n569), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n635), .A3(new_n634), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n826), .A2(new_n827), .A3(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(KEYINPUT118), .B(new_n813), .C1(new_n818), .C2(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n828), .A2(new_n747), .A3(new_n792), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT48), .Z(new_n838));
  NAND2_X1  g652(.A1(new_n815), .A2(new_n707), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(G952), .A3(new_n320), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n832), .B2(new_n636), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT119), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n834), .B(KEYINPUT51), .C1(new_n823), .C2(new_n824), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n836), .B(new_n843), .C1(new_n818), .C2(new_n844), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n818), .A2(new_n835), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT118), .B1(new_n846), .B2(new_n813), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n372), .A2(new_n664), .ZN(new_n848));
  NOR4_X1   g662(.A1(new_n848), .A2(new_n428), .A3(new_n640), .A4(new_n642), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n304), .A3(new_n187), .A4(new_n307), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n850), .A2(new_n615), .A3(new_n617), .A4(new_n658), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n851), .A2(new_n524), .B1(new_n764), .B2(new_n732), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n768), .A2(new_n775), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n727), .A2(new_n678), .A3(new_n187), .A4(new_n681), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n727), .B1(new_n308), .B2(new_n681), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n658), .A2(new_n691), .A3(new_n664), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n676), .B(new_n860), .C1(new_n757), .C2(new_n758), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n855), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n762), .B2(new_n763), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n729), .A2(KEYINPUT115), .A3(new_n676), .A4(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n687), .A2(new_n667), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n734), .A2(new_n735), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n734), .A2(new_n735), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n854), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n687), .A2(new_n667), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n733), .B2(new_n736), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n862), .A2(new_n864), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT52), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n853), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n702), .A2(new_n709), .A3(new_n705), .A4(new_n730), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT113), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n707), .A2(new_n708), .B1(new_n724), .B2(new_n729), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n879), .A2(KEYINPUT113), .A3(new_n702), .A4(new_n705), .ZN(new_n880));
  INV_X1    g694(.A(new_n636), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(new_n373), .B2(new_n680), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n622), .A2(new_n627), .A3(new_n618), .A4(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(new_n619), .A3(new_n655), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT114), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n883), .A2(new_n619), .A3(new_n655), .A4(KEYINPUT114), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n878), .A2(new_n880), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT53), .B1(new_n875), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n760), .A2(new_n852), .A3(new_n767), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n772), .B2(new_n774), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT52), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT52), .B1(new_n872), .B2(new_n873), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n878), .A2(new_n888), .A3(new_n880), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n890), .B1(new_n898), .B2(KEYINPUT116), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(KEYINPUT116), .B2(new_n898), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT54), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n876), .A2(new_n896), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n892), .A2(new_n888), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n893), .A2(new_n894), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n890), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n845), .A2(new_n847), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(G952), .A2(G953), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n812), .B1(new_n910), .B2(new_n911), .ZN(G75));
  NOR2_X1   g726(.A1(new_n320), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n906), .A2(new_n368), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT56), .B1(new_n915), .B2(G210), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n302), .B(new_n281), .ZN(new_n917));
  XOR2_X1   g731(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n914), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n916), .B2(new_n919), .ZN(G51));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n890), .A2(new_n905), .A3(KEYINPUT121), .A4(KEYINPUT54), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT54), .B1(new_n890), .B2(new_n905), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n923), .B1(new_n926), .B2(new_n908), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n754), .B(KEYINPUT57), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n922), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n906), .A2(new_n925), .A3(new_n907), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n870), .A2(new_n874), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n932), .A2(new_n888), .A3(new_n892), .A4(new_n902), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT121), .B1(new_n934), .B2(KEYINPUT54), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(KEYINPUT54), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n930), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n928), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n937), .A2(KEYINPUT122), .A3(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n929), .A2(KEYINPUT123), .A3(new_n607), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n915), .A2(new_n779), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n929), .A2(new_n607), .A3(new_n939), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT123), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n913), .B1(new_n942), .B2(new_n945), .ZN(G54));
  NAND3_X1  g760(.A1(new_n915), .A2(KEYINPUT58), .A3(G475), .ZN(new_n947));
  INV_X1    g761(.A(new_n361), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n913), .ZN(G60));
  NOR2_X1   g765(.A1(new_n630), .A2(new_n631), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT59), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n953), .B1(new_n909), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n953), .A2(new_n956), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n914), .B1(new_n927), .B2(new_n958), .ZN(new_n959));
  OR3_X1    g773(.A1(new_n957), .A2(KEYINPUT124), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT124), .B1(new_n957), .B2(new_n959), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(G63));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT60), .Z(new_n964));
  NAND2_X1  g778(.A1(new_n934), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n965), .A2(KEYINPUT125), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(KEYINPUT125), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT126), .B1(new_n969), .B2(new_n652), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n970), .A2(KEYINPUT61), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n913), .B1(new_n969), .B2(new_n652), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n967), .A2(new_n556), .A3(new_n555), .A4(new_n968), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n973), .B(new_n972), .C1(new_n970), .C2(KEYINPUT61), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(G66));
  NOR3_X1   g791(.A1(new_n434), .A2(new_n276), .A3(new_n320), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n889), .B2(new_n320), .ZN(new_n979));
  INV_X1    g793(.A(new_n302), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(G898), .B2(new_n320), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n979), .B(new_n981), .ZN(G69));
  XOR2_X1   g796(.A(new_n504), .B(new_n333), .Z(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(new_n588), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n984), .A2(new_n660), .A3(new_n320), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n787), .A2(new_n858), .A3(new_n747), .ZN(new_n986));
  INV_X1    g800(.A(new_n768), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n986), .A2(new_n796), .A3(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n807), .A2(new_n988), .A3(new_n775), .A4(new_n872), .ZN(new_n989));
  INV_X1    g803(.A(new_n983), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n683), .A2(new_n872), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT62), .Z(new_n993));
  AND4_X1   g807(.A1(new_n618), .A2(new_n788), .A3(new_n669), .A4(new_n882), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n796), .B1(new_n690), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n807), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n991), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n985), .B1(new_n997), .B2(new_n320), .ZN(G72));
  NAND2_X1  g812(.A1(new_n505), .A2(new_n442), .ZN(new_n999));
  OR2_X1    g813(.A1(new_n505), .A2(new_n442), .ZN(new_n1000));
  OAI22_X1  g814(.A1(new_n989), .A2(new_n999), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n889), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1000), .A2(new_n999), .ZN(new_n1003));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT63), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT127), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n913), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1002), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1008), .B1(new_n900), .B2(new_n1009), .ZN(G57));
endmodule


