//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n205));
  AND2_X1   g004(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(G190gat), .ZN(new_n207));
  INV_X1    g006(.A(G169gat), .ZN(new_n208));
  INV_X1    g007(.A(G176gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT23), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G169gat), .B2(G176gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n203), .B1(new_n207), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n205), .A2(new_n204), .ZN(new_n216));
  NAND3_X1  g015(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  AOI22_X1  g019(.A1(KEYINPUT65), .A2(new_n219), .B1(new_n220), .B2(KEYINPUT23), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n208), .A2(new_n209), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n203), .B1(new_n223), .B2(new_n211), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n218), .A2(new_n221), .A3(new_n222), .A4(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G183gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT27), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT27), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT28), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n227), .A2(new_n229), .A3(KEYINPUT28), .A4(new_n230), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n204), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n219), .B1(new_n223), .B2(KEYINPUT26), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT26), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n236), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n215), .A2(new_n225), .B1(new_n235), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n202), .B1(new_n241), .B2(KEYINPUT29), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n215), .A2(new_n225), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT27), .B(G183gat), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT28), .B1(new_n245), .B2(new_n230), .ZN(new_n246));
  INV_X1    g045(.A(new_n234), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n237), .A2(new_n239), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n204), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n244), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n235), .A2(KEYINPUT66), .A3(new_n240), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n243), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n242), .B(KEYINPUT74), .C1(new_n253), .C2(new_n202), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n215), .A2(new_n225), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n235), .A2(KEYINPUT66), .A3(new_n240), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT66), .B1(new_n235), .B2(new_n240), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT74), .ZN(new_n259));
  INV_X1    g058(.A(new_n202), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(G197gat), .A2(G204gat), .ZN(new_n263));
  AND2_X1   g062(.A1(G197gat), .A2(G204gat), .ZN(new_n264));
  AND2_X1   g063(.A1(G211gat), .A2(G218gat), .ZN(new_n265));
  OAI22_X1  g064(.A1(new_n263), .A2(new_n264), .B1(new_n265), .B2(KEYINPUT22), .ZN(new_n266));
  XNOR2_X1  g065(.A(G211gat), .B(G218gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n260), .A2(KEYINPUT29), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n258), .A2(new_n271), .B1(new_n260), .B2(new_n241), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n268), .ZN(new_n273));
  XNOR2_X1  g072(.A(G8gat), .B(G36gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n274), .B(new_n275), .Z(new_n276));
  NAND3_X1  g075(.A1(new_n270), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n276), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n268), .B1(new_n254), .B2(new_n261), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n272), .A2(new_n268), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n277), .A2(new_n281), .A3(KEYINPUT30), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n270), .A2(new_n283), .A3(new_n273), .A4(new_n276), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G1gat), .B(G29gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT0), .ZN(new_n287));
  XNOR2_X1  g086(.A(G57gat), .B(G85gat), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n287), .B(new_n288), .Z(new_n289));
  INV_X1    g088(.A(KEYINPUT1), .ZN(new_n290));
  INV_X1    g089(.A(G120gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(G113gat), .ZN(new_n292));
  INV_X1    g091(.A(G113gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(G120gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n290), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(G127gat), .B(G134gat), .Z(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n298));
  OR2_X1    g097(.A1(KEYINPUT67), .A2(G120gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n300));
  NAND2_X1  g099(.A1(KEYINPUT67), .A2(G120gat), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n299), .A2(new_n300), .A3(G113gat), .A4(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(KEYINPUT67), .A2(G120gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(KEYINPUT67), .A2(G120gat), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n303), .A2(new_n304), .A3(new_n293), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n292), .A2(KEYINPUT68), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n298), .B(new_n302), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n296), .A2(KEYINPUT1), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT67), .B(G120gat), .ZN(new_n310));
  OAI22_X1  g109(.A1(new_n310), .A2(new_n293), .B1(KEYINPUT68), .B2(new_n292), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n298), .B1(new_n311), .B2(new_n302), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n297), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G141gat), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G155gat), .ZN(new_n322));
  INV_X1    g121(.A(G162gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT76), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G162gat), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n322), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n318), .B(new_n321), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT75), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n319), .B2(new_n320), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n328), .A3(new_n317), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n313), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT79), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n316), .B(new_n317), .C1(new_n319), .C2(new_n320), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n325), .A2(G162gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n323), .A2(KEYINPUT76), .ZN(new_n340));
  OAI21_X1  g139(.A(G155gat), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n338), .B1(new_n341), .B2(KEYINPUT2), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n344), .B(new_n297), .C1(new_n309), .C2(new_n312), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n336), .A2(new_n337), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n313), .A2(KEYINPUT79), .A3(new_n335), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n297), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n307), .A2(new_n308), .ZN(new_n352));
  INV_X1    g151(.A(new_n312), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n329), .A2(new_n355), .A3(new_n334), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n355), .B1(new_n329), .B2(new_n334), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n354), .A2(new_n358), .A3(KEYINPUT4), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT3), .B1(new_n342), .B2(new_n343), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT77), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n335), .A2(new_n362), .A3(KEYINPUT3), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n361), .A2(new_n313), .A3(new_n363), .A4(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n345), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n359), .A2(new_n366), .A3(new_n347), .A4(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n369), .A3(KEYINPUT5), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n335), .A2(KEYINPUT78), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n329), .A2(new_n355), .A3(new_n334), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n367), .B1(new_n373), .B2(new_n313), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n354), .A2(KEYINPUT4), .A3(new_n344), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n348), .A2(KEYINPUT5), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n374), .A2(new_n375), .A3(new_n366), .A4(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n289), .B1(new_n370), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n285), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT39), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n374), .A2(new_n375), .A3(new_n366), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n382), .A3(new_n348), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n382), .B1(new_n381), .B2(new_n348), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n385), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n346), .A2(new_n349), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n380), .B1(new_n388), .B2(new_n347), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(new_n383), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n390), .A3(new_n289), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT40), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n386), .A2(new_n390), .A3(KEYINPUT40), .A4(new_n289), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(G22gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT31), .B(G50gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT29), .B1(new_n344), .B2(new_n364), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(new_n269), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n364), .B1(new_n268), .B2(KEYINPUT29), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n402), .A2(new_n335), .ZN(new_n403));
  OAI211_X1 g202(.A(G228gat), .B(G233gat), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n373), .A2(new_n402), .ZN(new_n405));
  NAND2_X1  g204(.A1(G228gat), .A2(G233gat), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n405), .B(new_n406), .C1(new_n269), .C2(new_n400), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n399), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n404), .A2(new_n407), .A3(new_n399), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n397), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n410), .ZN(new_n412));
  INV_X1    g211(.A(new_n397), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n412), .A2(new_n413), .A3(new_n408), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n277), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT37), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n270), .A2(new_n417), .A3(new_n273), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT83), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT83), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n270), .A2(new_n420), .A3(new_n417), .A4(new_n273), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n262), .A2(new_n268), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n417), .B1(new_n272), .B2(new_n269), .ZN(new_n424));
  AOI211_X1 g223(.A(KEYINPUT38), .B(new_n276), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n416), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n370), .A2(new_n377), .ZN(new_n427));
  INV_X1    g226(.A(new_n289), .ZN(new_n428));
  AND4_X1   g227(.A1(KEYINPUT81), .A2(new_n427), .A3(KEYINPUT6), .A4(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT81), .B1(new_n378), .B2(KEYINPUT6), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n378), .A2(KEYINPUT6), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n370), .A2(new_n289), .A3(new_n377), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT80), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n433), .A2(new_n434), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n432), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n426), .A2(new_n431), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT38), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT37), .B1(new_n279), .B2(new_n280), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT84), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n440), .A2(new_n441), .A3(new_n278), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n440), .B2(new_n278), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n439), .B1(new_n444), .B2(new_n422), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n395), .B(new_n415), .C1(new_n438), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n437), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n285), .ZN(new_n448));
  INV_X1    g247(.A(new_n415), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT70), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(new_n258), .B2(new_n313), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n251), .A2(new_n252), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n354), .A2(new_n453), .A3(KEYINPUT70), .A4(new_n255), .ZN(new_n454));
  NAND2_X1  g253(.A1(G227gat), .A2(G233gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT64), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n258), .A2(new_n313), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n452), .A2(new_n454), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT34), .B1(new_n459), .B2(KEYINPUT71), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT32), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n452), .A2(new_n454), .A3(new_n458), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n464), .B1(new_n465), .B2(new_n456), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT33), .B1(new_n465), .B2(new_n456), .ZN(new_n467));
  XOR2_X1   g266(.A(G15gat), .B(G43gat), .Z(new_n468));
  XNOR2_X1  g267(.A(G71gat), .B(G99gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n466), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  AOI221_X4 g271(.A(new_n464), .B1(KEYINPUT33), .B2(new_n470), .C1(new_n465), .C2(new_n456), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n463), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n465), .A2(new_n456), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT33), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n471), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n466), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n473), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n459), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(new_n460), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n474), .A2(KEYINPUT73), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT36), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT73), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n486), .B(new_n463), .C1(new_n472), .C2(new_n473), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT72), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(KEYINPUT72), .B(new_n463), .C1(new_n472), .C2(new_n473), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n490), .A2(KEYINPUT36), .A3(new_n483), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n446), .A2(new_n450), .A3(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n490), .A2(new_n483), .A3(new_n491), .A4(new_n415), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT86), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n491), .A2(new_n483), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n497), .A2(new_n498), .A3(new_n490), .A4(new_n415), .ZN(new_n499));
  INV_X1    g298(.A(new_n285), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n431), .B2(new_n437), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n496), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n484), .A2(new_n487), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT35), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n415), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  AND4_X1   g306(.A1(KEYINPUT85), .A2(new_n504), .A3(new_n501), .A4(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n506), .B1(new_n484), .B2(new_n487), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT85), .B1(new_n509), .B2(new_n501), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n494), .B1(new_n503), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G113gat), .B(G141gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G169gat), .B(G197gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n517), .B(KEYINPUT12), .Z(new_n518));
  XOR2_X1   g317(.A(G43gat), .B(G50gat), .Z(new_n519));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(KEYINPUT90), .B(G36gat), .Z(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT89), .B(G29gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(G29gat), .A2(G36gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT14), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(KEYINPUT88), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n526), .A2(KEYINPUT88), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n521), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n519), .A2(new_n520), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n519), .A2(new_n520), .ZN(new_n531));
  NOR4_X1   g330(.A1(new_n530), .A2(new_n531), .A3(new_n524), .A4(new_n526), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534));
  INV_X1    g333(.A(G1gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(KEYINPUT16), .A3(new_n535), .ZN(new_n536));
  OR2_X1    g335(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n536), .B(new_n537), .C1(new_n535), .C2(new_n534), .ZN(new_n538));
  NAND2_X1  g337(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n538), .B(new_n539), .Z(new_n540));
  NOR2_X1   g339(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n533), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT17), .B1(new_n529), .B2(new_n532), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n538), .B(new_n539), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n541), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT93), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT18), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n541), .A2(KEYINPUT94), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n541), .A2(KEYINPUT94), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n533), .A2(new_n540), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n550), .B(KEYINPUT13), .Z(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(new_n551), .B2(new_n552), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n518), .B1(new_n554), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n549), .A2(new_n550), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT18), .B1(new_n563), .B2(KEYINPUT93), .ZN(new_n564));
  INV_X1    g363(.A(new_n518), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n564), .A2(new_n553), .A3(new_n560), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G85gat), .A2(G92gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT7), .ZN(new_n570));
  INV_X1    g369(.A(G99gat), .ZN(new_n571));
  INV_X1    g370(.A(G106gat), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT8), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT98), .B(G85gat), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n570), .B(new_n573), .C1(G92gat), .C2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G99gat), .B(G106gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  INV_X1    g376(.A(KEYINPUT99), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n575), .B(new_n576), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT99), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n579), .B(new_n581), .C1(new_n529), .C2(new_n532), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT100), .ZN(new_n583));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT41), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n582), .A2(new_n583), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n583), .B1(new_n582), .B2(new_n587), .ZN(new_n589));
  INV_X1    g388(.A(new_n545), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n579), .A2(new_n581), .ZN(new_n591));
  OAI22_X1  g390(.A1(new_n588), .A2(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT101), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n584), .A2(new_n585), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n595), .B(G134gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(new_n323), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n590), .A2(new_n591), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n587), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT100), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n582), .A2(new_n583), .A3(new_n587), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n593), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n592), .A2(new_n593), .ZN(new_n606));
  OAI22_X1  g405(.A1(new_n594), .A2(new_n598), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n604), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n608), .A2(new_n609), .A3(KEYINPUT101), .A4(new_n597), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G71gat), .B(G78gat), .Z(new_n612));
  XNOR2_X1  g411(.A(G57gat), .B(G64gat), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT95), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT9), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n612), .B1(new_n618), .B2(new_n613), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G127gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n620), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n546), .B1(KEYINPUT21), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT97), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n625), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G155gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G183gat), .B(G211gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n629), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n611), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n579), .A2(KEYINPUT10), .A3(new_n581), .A4(new_n626), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n577), .A2(new_n620), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n580), .A2(new_n626), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(G230gat), .ZN(new_n643));
  INV_X1    g442(.A(G233gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n638), .A2(new_n640), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n647), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n647), .B(new_n652), .C1(new_n646), .C2(new_n648), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n649), .A2(KEYINPUT102), .A3(new_n653), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n636), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n512), .A2(new_n568), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n447), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g463(.A(KEYINPUT16), .B(G8gat), .Z(new_n665));
  NAND3_X1  g464(.A1(new_n661), .A2(new_n500), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n661), .ZN(new_n669));
  OAI21_X1  g468(.A(G8gat), .B1(new_n669), .B2(new_n285), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n666), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n668), .B1(new_n671), .B2(KEYINPUT42), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT103), .ZN(G1325gat));
  INV_X1    g472(.A(new_n504), .ZN(new_n674));
  OR3_X1    g473(.A1(new_n669), .A2(G15gat), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n493), .B(KEYINPUT104), .Z(new_n676));
  OAI21_X1  g475(.A(G15gat), .B1(new_n669), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT105), .Z(G1326gat));
  NAND2_X1  g478(.A1(new_n661), .A2(new_n449), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  INV_X1    g481(.A(new_n659), .ZN(new_n683));
  INV_X1    g482(.A(new_n611), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n634), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR4_X1   g485(.A1(new_n512), .A2(new_n568), .A3(new_n683), .A4(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(new_n662), .A3(new_n523), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT45), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n659), .B(KEYINPUT106), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n690), .A2(new_n568), .A3(new_n634), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n494), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n509), .A2(new_n501), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT85), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n509), .A2(KEYINPUT85), .A3(new_n501), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n693), .B1(new_n694), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(new_n701), .A3(new_n611), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT44), .B1(new_n512), .B2(new_n684), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n692), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n447), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n689), .B1(new_n523), .B2(new_n706), .ZN(G1328gat));
  NAND3_X1  g506(.A1(new_n687), .A2(new_n522), .A3(new_n500), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT46), .Z(new_n709));
  NOR2_X1   g508(.A1(new_n705), .A2(new_n285), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n522), .B2(new_n710), .ZN(G1329gat));
  OR2_X1    g510(.A1(new_n705), .A2(new_n676), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n674), .A2(G43gat), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n712), .A2(G43gat), .B1(new_n687), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(G43gat), .ZN(new_n715));
  INV_X1    g514(.A(new_n493), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n704), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n687), .A2(new_n713), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT47), .ZN(new_n719));
  OAI22_X1  g518(.A1(new_n714), .A2(KEYINPUT47), .B1(new_n717), .B2(new_n719), .ZN(G1330gat));
  INV_X1    g519(.A(KEYINPUT48), .ZN(new_n721));
  INV_X1    g520(.A(G50gat), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n704), .B2(new_n449), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n687), .A2(new_n722), .A3(new_n449), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n721), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n705), .B2(new_n415), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n704), .A2(KEYINPUT107), .A3(new_n449), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n727), .A2(G50gat), .A3(new_n728), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n724), .A2(new_n721), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n725), .B1(new_n729), .B2(new_n730), .ZN(G1331gat));
  NAND2_X1  g530(.A1(new_n511), .A2(new_n503), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n567), .B1(new_n732), .B2(new_n693), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(new_n636), .A3(new_n690), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n447), .B(KEYINPUT108), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g537(.A1(new_n734), .A2(new_n285), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n734), .B2(new_n676), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n674), .A2(G71gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n734), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g546(.A1(new_n735), .A2(new_n449), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G78gat), .ZN(G1335gat));
  NAND4_X1  g548(.A1(new_n700), .A2(KEYINPUT51), .A3(new_n568), .A4(new_n685), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n733), .A2(KEYINPUT110), .A3(KEYINPUT51), .A4(new_n685), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n700), .A2(new_n568), .A3(new_n685), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n752), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n447), .A2(new_n574), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n757), .A2(new_n683), .A3(new_n758), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n567), .A2(new_n634), .A3(new_n659), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n701), .B1(new_n700), .B2(new_n611), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n512), .A2(KEYINPUT44), .A3(new_n684), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT109), .B1(new_n763), .B2(new_n447), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n574), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n763), .A2(KEYINPUT109), .A3(new_n447), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n759), .B1(new_n765), .B2(new_n766), .ZN(G1336gat));
  INV_X1    g566(.A(new_n690), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n768), .A2(G92gat), .A3(new_n285), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n757), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G92gat), .B1(new_n763), .B2(new_n285), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT113), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n772), .A2(KEYINPUT113), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n770), .A2(new_n771), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n512), .A2(new_n567), .A3(new_n686), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n755), .B1(new_n777), .B2(KEYINPUT111), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n754), .A2(new_n779), .A3(KEYINPUT51), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n778), .A2(new_n780), .A3(new_n769), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n771), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n776), .B1(new_n782), .B2(KEYINPUT52), .ZN(new_n783));
  AOI211_X1 g582(.A(KEYINPUT112), .B(new_n772), .C1(new_n771), .C2(new_n781), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n775), .B1(new_n783), .B2(new_n784), .ZN(G1337gat));
  NAND4_X1  g584(.A1(new_n757), .A2(new_n571), .A3(new_n504), .A4(new_n683), .ZN(new_n786));
  OAI21_X1  g585(.A(G99gat), .B1(new_n763), .B2(new_n676), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(G1338gat));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n449), .B(new_n760), .C1(new_n761), .C2(new_n762), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT53), .B1(new_n790), .B2(G106gat), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n768), .A2(G106gat), .A3(new_n415), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n757), .A2(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n790), .A2(G106gat), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n778), .A2(new_n780), .A3(new_n792), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n789), .B1(new_n794), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n791), .A2(new_n793), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n796), .A2(new_n797), .ZN(new_n801));
  OAI211_X1 g600(.A(KEYINPUT114), .B(new_n800), .C1(new_n801), .C2(new_n795), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n802), .ZN(G1339gat));
  NAND3_X1  g602(.A1(new_n637), .A2(new_n645), .A3(new_n641), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n647), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n645), .B1(new_n637), .B2(new_n641), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n652), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n805), .A2(KEYINPUT55), .A3(new_n808), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n656), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT115), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n811), .A2(new_n815), .A3(new_n656), .A4(new_n812), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n567), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n558), .A2(new_n559), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n549), .A2(new_n550), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n517), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n566), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n683), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n611), .B1(new_n817), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n610), .A3(new_n607), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n814), .A2(new_n816), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n635), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n636), .A2(new_n568), .A3(new_n659), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n736), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n496), .A2(new_n499), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n285), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n293), .A3(new_n567), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n449), .B1(new_n827), .B2(new_n828), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n662), .A2(new_n285), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n674), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n568), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n836), .A2(new_n842), .ZN(G1340gat));
  NOR2_X1   g642(.A1(new_n659), .A2(new_n310), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n835), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n291), .B1(new_n840), .B2(new_n690), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n846), .B(KEYINPUT117), .Z(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(G1341gat));
  AND3_X1   g647(.A1(new_n840), .A2(G127gat), .A3(new_n634), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n635), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT118), .ZN(new_n851));
  AOI21_X1  g650(.A(G127gat), .B1(new_n850), .B2(KEYINPUT118), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(G1342gat));
  NAND2_X1  g652(.A1(new_n611), .A2(new_n285), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT119), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(G134gat), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n832), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT56), .Z(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n841), .B2(new_n684), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1343gat));
  INV_X1    g659(.A(new_n828), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n822), .B1(new_n568), .B2(new_n813), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n684), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n825), .B2(new_n824), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n861), .B1(new_n864), .B2(new_n635), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT57), .B1(new_n865), .B2(new_n415), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n716), .A2(new_n838), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n829), .A2(new_n449), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n866), .B(new_n867), .C1(KEYINPUT57), .C2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G141gat), .B1(new_n869), .B2(new_n568), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n676), .A2(new_n449), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n830), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n500), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n567), .A2(new_n314), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT120), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT58), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n870), .A2(new_n879), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1344gat));
  NAND2_X1  g680(.A1(new_n868), .A2(KEYINPUT57), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n415), .A2(KEYINPUT57), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n824), .A2(new_n813), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n634), .B1(new_n863), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n883), .B1(new_n885), .B2(new_n861), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n882), .A2(new_n683), .A3(new_n867), .A4(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(G148gat), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT59), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n315), .A2(KEYINPUT59), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n869), .B2(new_n659), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n873), .A2(new_n315), .A3(new_n683), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1345gat));
  OAI21_X1  g695(.A(G155gat), .B1(new_n869), .B2(new_n635), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n873), .A2(new_n322), .A3(new_n634), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1346gat));
  NAND2_X1  g698(.A1(new_n324), .A2(new_n326), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n900), .B1(new_n869), .B2(new_n684), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n855), .A2(new_n900), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n872), .B2(new_n902), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n662), .A2(new_n285), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n829), .A2(new_n831), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n208), .A3(new_n567), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT122), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n736), .A2(new_n674), .A3(new_n285), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n837), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n568), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n910), .ZN(G1348gat));
  NAND3_X1  g710(.A1(new_n905), .A2(new_n209), .A3(new_n683), .ZN(new_n912));
  OAI21_X1  g711(.A(G176gat), .B1(new_n909), .B2(new_n768), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1349gat));
  NAND3_X1  g713(.A1(new_n905), .A2(new_n245), .A3(new_n634), .ZN(new_n915));
  OAI21_X1  g714(.A(G183gat), .B1(new_n909), .B2(new_n635), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n909), .B2(new_n684), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n919), .A2(KEYINPUT123), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(KEYINPUT123), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(KEYINPUT61), .A3(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n919), .A2(KEYINPUT123), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n905), .A2(new_n230), .A3(new_n611), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(G1351gat));
  NOR2_X1   g725(.A1(new_n736), .A2(new_n285), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n676), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT57), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n415), .B1(new_n827), .B2(new_n828), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n886), .B(new_n928), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(G197gat), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n931), .A2(new_n932), .A3(new_n568), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n829), .A2(new_n904), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n676), .A2(new_n449), .ZN(new_n935));
  OAI21_X1  g734(.A(KEYINPUT124), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n871), .A2(new_n829), .A3(new_n937), .A4(new_n904), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n567), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n933), .B1(new_n940), .B2(new_n932), .ZN(G1352gat));
  NOR4_X1   g740(.A1(new_n934), .A2(new_n935), .A3(G204gat), .A4(new_n659), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT62), .ZN(new_n943));
  OAI21_X1  g742(.A(G204gat), .B1(new_n931), .B2(new_n768), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1353gat));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n946));
  OAI211_X1 g745(.A(KEYINPUT63), .B(G211gat), .C1(new_n931), .C2(new_n635), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n882), .A2(new_n634), .A3(new_n886), .A4(new_n928), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT63), .B1(new_n949), .B2(G211gat), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n635), .A2(G211gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n938), .A3(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n936), .A2(new_n938), .A3(KEYINPUT125), .A4(new_n952), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n946), .B1(new_n951), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n955), .A2(new_n956), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n959), .B(KEYINPUT126), .C1(new_n950), .C2(new_n948), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1354gat));
  AOI21_X1  g760(.A(G218gat), .B1(new_n939), .B2(new_n611), .ZN(new_n962));
  INV_X1    g761(.A(new_n931), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n611), .A2(G218gat), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT127), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n962), .B1(new_n963), .B2(new_n965), .ZN(G1355gat));
endmodule


