//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G137), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT11), .A3(G134), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G131), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT64), .A2(G131), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT64), .A2(G131), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n200), .A2(new_n192), .A3(new_n194), .A4(new_n195), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n203), .A2(KEYINPUT3), .A3(G107), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G104), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(G104), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT83), .B1(new_n209), .B2(KEYINPUT3), .ZN(new_n210));
  OAI211_X1 g024(.A(KEYINPUT83), .B(KEYINPUT3), .C1(new_n203), .C2(G107), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n207), .B(new_n208), .C1(new_n210), .C2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n203), .A2(G107), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n208), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  INV_X1    g032(.A(G143), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G146), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n218), .B(new_n220), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n220), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(G128), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n213), .A2(new_n216), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT84), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n213), .A2(new_n222), .A3(new_n225), .A4(new_n216), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n213), .A2(new_n216), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(new_n222), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n202), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT12), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n228), .A2(new_n227), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n230), .A2(new_n231), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n232), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT12), .A3(new_n202), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT83), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n211), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n208), .B1(new_n246), .B2(new_n207), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n218), .A2(new_n220), .A3(KEYINPUT0), .A4(G128), .ZN(new_n250));
  XNOR2_X1  g064(.A(G143), .B(G146), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT0), .B(G128), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n213), .A2(KEYINPUT4), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n249), .B(new_n254), .C1(new_n247), .C2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n202), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT10), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n228), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n214), .B1(new_n209), .B2(KEYINPUT3), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n245), .B2(new_n211), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n215), .B1(new_n261), .B2(new_n208), .ZN(new_n262));
  INV_X1    g076(.A(new_n231), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(KEYINPUT10), .A3(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n256), .A2(new_n257), .A3(new_n259), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n242), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G227), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT82), .ZN(new_n269));
  XNOR2_X1  g083(.A(G110), .B(G140), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n256), .A2(new_n259), .A3(new_n264), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n202), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n265), .A2(new_n271), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n266), .A2(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(G469), .B1(new_n276), .B2(G902), .ZN(new_n277));
  INV_X1    g091(.A(G469), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT71), .B(G902), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n265), .A2(new_n271), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n236), .B2(new_n241), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n271), .B1(new_n274), .B2(new_n265), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n278), .B(new_n279), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n189), .B1(new_n277), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G125), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n231), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n253), .A2(G125), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G224), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n289), .A2(G953), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n288), .A2(new_n290), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n290), .A2(KEYINPUT7), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(G110), .B(G122), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n296), .B(KEYINPUT8), .ZN(new_n297));
  INV_X1    g111(.A(G119), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G116), .ZN(new_n299));
  INV_X1    g113(.A(G116), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G119), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT2), .B(G113), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT66), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(G116), .B(G119), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT66), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(G113), .ZN(new_n308));
  INV_X1    g122(.A(G113), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(KEYINPUT2), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n305), .B(new_n306), .C1(new_n308), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n305), .A2(KEYINPUT5), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT5), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(new_n298), .A3(G116), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n313), .A2(KEYINPUT85), .A3(G113), .A4(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT85), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n299), .A2(new_n301), .A3(KEYINPUT5), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n315), .A2(G113), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n312), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n297), .B1(new_n321), .B2(new_n262), .ZN(new_n322));
  OAI211_X1 g136(.A(G113), .B(new_n315), .C1(new_n302), .C2(new_n314), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n312), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n322), .B1(new_n262), .B2(new_n324), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n288), .A2(new_n294), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n295), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT86), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n321), .B2(new_n230), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n311), .A2(new_n304), .B1(new_n323), .B2(new_n317), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n330), .A2(new_n262), .A3(KEYINPUT86), .A4(new_n316), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n248), .B1(new_n261), .B2(new_n208), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n333), .B1(new_n208), .B2(new_n261), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n302), .A2(new_n303), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n248), .A2(new_n247), .B1(new_n312), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n332), .A2(new_n296), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT87), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n329), .A2(new_n331), .B1(new_n334), .B2(new_n336), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT87), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(new_n296), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(G902), .B1(new_n327), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n332), .A2(new_n337), .ZN(new_n345));
  INV_X1    g159(.A(new_n296), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT6), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AND4_X1   g163(.A1(new_n341), .A2(new_n332), .A3(new_n296), .A4(new_n337), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n341), .B1(new_n340), .B2(new_n296), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT6), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n349), .B1(new_n352), .B2(new_n347), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n344), .B1(new_n353), .B2(new_n293), .ZN(new_n354));
  OAI21_X1  g168(.A(G210), .B1(G237), .B2(G902), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n349), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n348), .B1(new_n339), .B2(new_n342), .ZN(new_n359));
  INV_X1    g173(.A(new_n347), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n293), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n355), .A3(new_n344), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n357), .A2(KEYINPUT88), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G214), .B1(G237), .B2(G902), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n355), .B1(new_n363), .B2(new_n344), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT88), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AND4_X1   g183(.A1(new_n284), .A2(new_n365), .A3(new_n366), .A4(new_n369), .ZN(new_n370));
  XOR2_X1   g184(.A(KEYINPUT73), .B(G217), .Z(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(G234), .B2(new_n279), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(KEYINPUT25), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT78), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT22), .B(G137), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(KEYINPUT79), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT75), .B1(new_n285), .B2(G140), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT74), .B(G140), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n381), .B1(new_n382), .B2(new_n285), .ZN(new_n383));
  INV_X1    g197(.A(G140), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n384), .A2(KEYINPUT74), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(KEYINPUT74), .ZN(new_n386));
  OAI211_X1 g200(.A(KEYINPUT75), .B(G125), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(G125), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT16), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(new_n217), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT76), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n388), .A2(new_n391), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G146), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n388), .A2(KEYINPUT76), .A3(new_n217), .A4(new_n391), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT23), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n298), .B2(G128), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n221), .A2(KEYINPUT23), .A3(G119), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n400), .B(new_n401), .C1(G119), .C2(new_n221), .ZN(new_n402));
  XNOR2_X1  g216(.A(G119), .B(G128), .ZN(new_n403));
  XOR2_X1   g217(.A(KEYINPUT24), .B(G110), .Z(new_n404));
  AOI22_X1  g218(.A1(new_n402), .A2(G110), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n217), .B1(new_n388), .B2(new_n391), .ZN(new_n407));
  OAI22_X1  g221(.A1(new_n402), .A2(G110), .B1(new_n403), .B2(new_n404), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n285), .A2(G140), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT77), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n389), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n410), .B1(new_n389), .B2(new_n409), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n408), .B1(G146), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n407), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n380), .B1(new_n406), .B2(new_n416), .ZN(new_n417));
  AOI211_X1 g231(.A(new_n415), .B(new_n379), .C1(new_n398), .C2(new_n405), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n375), .B1(new_n419), .B2(new_n279), .ZN(new_n420));
  INV_X1    g234(.A(new_n279), .ZN(new_n421));
  NOR4_X1   g235(.A1(new_n417), .A2(new_n418), .A3(new_n421), .A4(new_n374), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n372), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(KEYINPUT81), .B(new_n372), .C1(new_n420), .C2(new_n422), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n372), .A2(G902), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n419), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(G134), .B(G137), .ZN(new_n430));
  INV_X1    g244(.A(G131), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT65), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n193), .A2(G134), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n195), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT65), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(G131), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n201), .A2(new_n432), .A3(new_n436), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n437), .A2(new_n231), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n254), .A2(new_n202), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n254), .B2(new_n202), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n438), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n312), .A2(new_n335), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n443), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n445), .B(new_n438), .C1(new_n440), .C2(new_n441), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(KEYINPUT69), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT69), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n442), .A2(new_n448), .A3(new_n443), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(KEYINPUT28), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n254), .A2(new_n202), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n438), .A2(new_n445), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT28), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT70), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT26), .B(G101), .ZN(new_n456));
  NOR2_X1   g270(.A1(G237), .A2(G953), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G210), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n456), .B(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT29), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n450), .A2(new_n455), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT30), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n438), .A2(new_n466), .A3(new_n451), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n437), .A2(new_n231), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n451), .A2(KEYINPUT67), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n253), .B1(new_n201), .B2(new_n197), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n439), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n468), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n467), .B1(new_n472), .B2(new_n466), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n443), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n461), .B1(new_n474), .B2(new_n446), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n443), .B1(new_n468), .B2(new_n470), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n454), .B(new_n476), .C1(new_n453), .C2(new_n446), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n463), .B1(new_n477), .B2(new_n462), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n465), .B(new_n279), .C1(new_n475), .C2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT72), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n479), .A2(new_n480), .A3(G472), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n480), .B1(new_n479), .B2(G472), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT30), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n442), .B2(KEYINPUT30), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n461), .B(new_n446), .C1(new_n485), .C2(new_n445), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT31), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT31), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n474), .A2(new_n488), .A3(new_n461), .A4(new_n446), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n477), .A2(new_n462), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(G472), .A2(G902), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT32), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT32), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n491), .A2(new_n495), .A3(new_n492), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n429), .B1(new_n483), .B2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT64), .B(G131), .ZN(new_n499));
  INV_X1    g313(.A(G237), .ZN(new_n500));
  AND4_X1   g314(.A1(G143), .A2(new_n500), .A3(new_n267), .A4(G214), .ZN(new_n501));
  AOI21_X1  g315(.A(G143), .B1(new_n457), .B2(G214), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n267), .A3(G214), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n219), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n457), .A2(G143), .A3(G214), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n200), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n503), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n507), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT17), .A3(new_n499), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n394), .A2(new_n396), .A3(new_n512), .A4(new_n397), .ZN(new_n513));
  XNOR2_X1  g327(.A(G113), .B(G122), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(new_n203), .ZN(new_n515));
  OAI211_X1 g329(.A(KEYINPUT18), .B(G131), .C1(new_n510), .C2(KEYINPUT89), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n510), .A2(KEYINPUT89), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n383), .A2(G146), .A3(new_n387), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n519), .B1(G146), .B2(new_n413), .ZN(new_n520));
  NAND2_X1  g334(.A1(KEYINPUT18), .A2(G131), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n518), .B(new_n520), .C1(new_n517), .C2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n513), .A2(new_n515), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT91), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n513), .A2(new_n525), .A3(new_n515), .A4(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT19), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n383), .B2(new_n387), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT19), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n217), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n396), .A2(KEYINPUT90), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n503), .A2(new_n508), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT90), .B1(new_n396), .B2(new_n531), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n522), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n515), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n527), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT92), .ZN(new_n540));
  NOR2_X1   g354(.A1(G475), .A2(G902), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT92), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n527), .A2(new_n542), .A3(new_n538), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n541), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(KEYINPUT20), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n544), .A2(KEYINPUT20), .B1(new_n539), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G475), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n515), .B1(new_n513), .B2(new_n522), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n549), .A2(KEYINPUT93), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(KEYINPUT93), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n527), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(G902), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n548), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n300), .A2(G122), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT14), .ZN(new_n556));
  AND2_X1   g370(.A1(KEYINPUT94), .A2(G122), .ZN(new_n557));
  NOR2_X1   g371(.A1(KEYINPUT94), .A2(G122), .ZN(new_n558));
  OAI21_X1  g372(.A(G116), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G107), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n205), .A3(new_n555), .ZN(new_n562));
  XNOR2_X1  g376(.A(G128), .B(G143), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(new_n191), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n559), .A2(new_n555), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G107), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n562), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT13), .B1(new_n221), .B2(G143), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(new_n191), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(new_n563), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n568), .A2(new_n571), .A3(KEYINPUT95), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT95), .B1(new_n568), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n565), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n371), .A2(G953), .A3(new_n187), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n565), .B(new_n575), .C1(new_n572), .C2(new_n573), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(KEYINPUT96), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n574), .A2(new_n580), .A3(new_n576), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n279), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G478), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(KEYINPUT15), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n584), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n547), .A2(new_n554), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(G952), .ZN(new_n589));
  AOI211_X1 g403(.A(G953), .B(new_n589), .C1(G234), .C2(G237), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT21), .B(G898), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT97), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  AOI211_X1 g407(.A(new_n267), .B(new_n279), .C1(G234), .C2(G237), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n590), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT98), .B1(new_n588), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n539), .A2(new_n546), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n527), .A2(new_n542), .A3(new_n538), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n542), .B1(new_n527), .B2(new_n538), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n599), .A2(new_n600), .A3(new_n545), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT20), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n554), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n585), .A2(new_n586), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n603), .A2(new_n596), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n370), .B(new_n498), .C1(new_n597), .C2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  NOR2_X1   g424(.A1(new_n354), .A2(new_n356), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n596), .B(new_n366), .C1(new_n611), .C2(new_n367), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n579), .A2(new_n613), .A3(new_n581), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n577), .A2(KEYINPUT33), .A3(new_n578), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n617), .A2(G478), .A3(new_n279), .ZN(new_n618));
  INV_X1    g432(.A(new_n582), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n618), .B1(G478), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n547), .B2(new_n554), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n612), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n276), .A2(G469), .ZN(new_n623));
  NAND2_X1  g437(.A1(G469), .A2(G902), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n283), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n188), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n491), .A2(new_n279), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(G472), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n493), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n429), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n622), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n634));
  INV_X1    g448(.A(new_n366), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n595), .B(new_n635), .C1(new_n357), .C2(new_n364), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n601), .A2(new_n602), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n544), .A2(KEYINPUT20), .ZN(new_n638));
  AOI211_X1 g452(.A(new_n554), .B(new_n605), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n634), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n599), .A2(new_n600), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n602), .B1(new_n641), .B2(new_n541), .ZN(new_n642));
  NOR4_X1   g456(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT20), .A4(new_n545), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n604), .B(new_n587), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n612), .A2(new_n644), .A3(KEYINPUT99), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n630), .B1(new_n640), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  INV_X1    g462(.A(new_n380), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(KEYINPUT36), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n406), .A2(new_n416), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n427), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n425), .A2(new_n426), .A3(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n629), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n370), .B(new_n656), .C1(new_n597), .C2(new_n608), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  OAI21_X1  g473(.A(new_n366), .B1(new_n611), .B2(new_n367), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n655), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n626), .B1(new_n483), .B2(new_n497), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n590), .B1(new_n594), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n644), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  XOR2_X1   g482(.A(new_n665), .B(KEYINPUT39), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n284), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n670), .A2(KEYINPUT40), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n547), .A2(new_n554), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n670), .B2(KEYINPUT40), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n474), .A2(new_n446), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n461), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n447), .A2(new_n449), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n676), .B(new_n553), .C1(new_n461), .C2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(G472), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n497), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n655), .A2(new_n680), .A3(new_n587), .A4(new_n366), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n674), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n365), .A2(new_n369), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n682), .A2(KEYINPUT101), .A3(new_n685), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n219), .ZN(G45));
  INV_X1    g505(.A(new_n665), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n620), .B(new_n692), .C1(new_n547), .C2(new_n554), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n663), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  NAND3_X1  g510(.A1(new_n479), .A2(new_n480), .A3(G472), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n279), .B1(new_n475), .B2(new_n478), .ZN(new_n698));
  INV_X1    g512(.A(new_n465), .ZN(new_n699));
  OAI21_X1  g513(.A(G472), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT72), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n497), .A2(new_n697), .A3(new_n701), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT12), .B1(new_n240), .B2(new_n202), .ZN(new_n704));
  AOI211_X1 g518(.A(new_n235), .B(new_n257), .C1(new_n239), .C2(new_n232), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n275), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n274), .A2(new_n265), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n272), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AOI211_X1 g523(.A(KEYINPUT102), .B(new_n278), .C1(new_n709), .C2(new_n279), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n279), .B1(new_n281), .B2(new_n282), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(G469), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(KEYINPUT102), .A3(new_n283), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n189), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n702), .A2(new_n703), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n622), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  OAI21_X1  g533(.A(new_n716), .B1(new_n640), .B2(new_n645), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  INV_X1    g535(.A(new_n715), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n660), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n702), .A2(new_n654), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n723), .B(new_n724), .C1(new_n597), .C2(new_n608), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  OAI211_X1 g540(.A(new_n587), .B(new_n366), .C1(new_n611), .C2(new_n367), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n672), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n283), .A2(KEYINPUT102), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n278), .B1(new_n709), .B2(new_n279), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n596), .B(new_n188), .C1(new_n731), .C2(new_n710), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n492), .B(KEYINPUT103), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n487), .A2(new_n489), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n461), .B1(new_n450), .B2(new_n455), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT104), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n738), .B(new_n733), .C1(new_n734), .C2(new_n735), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n737), .A2(new_n628), .A3(new_n739), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n732), .A2(new_n429), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n728), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NAND2_X1  g557(.A1(new_n693), .A2(KEYINPUT105), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n603), .A2(new_n604), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n746), .A3(new_n620), .A4(new_n692), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n655), .A2(new_n740), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n723), .A2(new_n744), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  AOI21_X1  g564(.A(new_n635), .B1(new_n365), .B2(new_n369), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n625), .A2(KEYINPUT106), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT106), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n277), .A2(new_n753), .A3(new_n283), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n752), .A2(new_n188), .A3(new_n754), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n751), .A2(new_n498), .A3(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n744), .A2(new_n747), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n757), .A3(KEYINPUT42), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT42), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n751), .A2(new_n498), .A3(new_n755), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n744), .A2(new_n747), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  AND4_X1   g578(.A1(new_n498), .A2(new_n666), .A3(new_n751), .A4(new_n755), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n191), .ZN(G36));
  NAND2_X1  g580(.A1(new_n275), .A2(new_n274), .ZN(new_n767));
  INV_X1    g581(.A(new_n266), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n767), .B1(new_n768), .B2(new_n271), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n278), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n276), .A2(KEYINPUT45), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n624), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT107), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n624), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n775), .A2(new_n283), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n781), .A2(new_n188), .A3(new_n669), .A4(new_n751), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n672), .A2(new_n620), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT43), .B1(new_n672), .B2(KEYINPUT108), .ZN(new_n784));
  XOR2_X1   g598(.A(new_n783), .B(new_n784), .Z(new_n785));
  NAND2_X1  g599(.A1(new_n654), .A2(new_n629), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT44), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n782), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n785), .A2(KEYINPUT44), .A3(new_n787), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  XOR2_X1   g607(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n794));
  AND3_X1   g608(.A1(new_n781), .A2(new_n188), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n781), .A2(new_n188), .B1(KEYINPUT109), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n751), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n799), .A2(new_n703), .A3(new_n702), .A4(new_n693), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G140), .ZN(G42));
  INV_X1    g616(.A(new_n685), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n731), .A2(new_n710), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n804), .B(KEYINPUT49), .Z(new_n805));
  NOR4_X1   g619(.A1(new_n680), .A2(new_n429), .A3(new_n189), .A4(new_n635), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n803), .A2(new_n783), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT110), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n783), .B(new_n784), .ZN(new_n810));
  INV_X1    g624(.A(new_n590), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n799), .A2(new_n722), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n814), .B(new_n815), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n809), .B(KEYINPUT48), .C1(new_n816), .C2(new_n498), .ZN(new_n817));
  XNOR2_X1  g631(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n816), .A2(new_n498), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n429), .A2(new_n740), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n812), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n821), .A2(new_n660), .A3(new_n722), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n680), .A2(new_n429), .A3(new_n811), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n813), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(G952), .B(new_n267), .C1(new_n824), .C2(new_n621), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n817), .A2(new_n819), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n821), .A2(new_n366), .A3(new_n685), .A4(new_n722), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT50), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n816), .A2(new_n748), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n824), .A2(new_n745), .A3(new_n620), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n821), .A2(new_n799), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n795), .A2(new_n797), .B1(new_n188), .B2(new_n804), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n828), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n826), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n683), .A2(new_n635), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n620), .B1(new_n603), .B2(new_n604), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n588), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n838), .A2(new_n840), .A3(new_n596), .A4(new_n630), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n609), .A2(new_n657), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n744), .A2(new_n748), .A3(new_n747), .A4(new_n755), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n655), .A2(new_n587), .A3(new_n665), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n554), .B1(new_n637), .B2(new_n638), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n845), .A3(new_n662), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n799), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n622), .A2(new_n716), .B1(new_n728), .B2(new_n741), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n720), .A2(new_n849), .A3(new_n725), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n765), .B1(new_n758), .B2(new_n762), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n720), .A2(new_n849), .A3(new_n725), .A4(KEYINPUT111), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n848), .A2(new_n852), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n425), .A2(new_n426), .A3(new_n653), .A4(new_n692), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT113), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(new_n680), .A3(new_n728), .A4(new_n755), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n661), .B(new_n662), .C1(new_n666), .C2(new_n694), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n859), .A3(new_n749), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT52), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n860), .B(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n864), .B2(KEYINPUT112), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n862), .B(new_n865), .Z(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT54), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(new_n855), .B2(new_n861), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n850), .A2(new_n868), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n864), .A2(new_n853), .A3(new_n848), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n834), .A2(new_n835), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n837), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(G952), .A2(G953), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n808), .B1(new_n876), .B2(new_n877), .ZN(G75));
  NAND2_X1  g692(.A1(new_n353), .A2(new_n293), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n363), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT55), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n279), .B(new_n355), .C1(new_n869), .C2(new_n872), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n881), .B1(new_n882), .B2(KEYINPUT56), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n267), .A2(G952), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n882), .A2(KEYINPUT116), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n881), .A2(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n882), .A2(KEYINPUT116), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n883), .B(new_n885), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT117), .ZN(G51));
  NAND2_X1  g705(.A1(new_n869), .A2(new_n872), .ZN(new_n892));
  INV_X1    g706(.A(new_n773), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n421), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT119), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n892), .A2(new_n896), .A3(new_n421), .A4(new_n893), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n709), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n624), .B(KEYINPUT57), .Z(new_n900));
  AND3_X1   g714(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n870), .B1(new_n869), .B2(new_n872), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n899), .B1(new_n903), .B2(KEYINPUT118), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT118), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n905), .B(new_n900), .C1(new_n901), .C2(new_n902), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n898), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT120), .B1(new_n907), .B2(new_n884), .ZN(new_n908));
  INV_X1    g722(.A(new_n898), .ZN(new_n909));
  INV_X1    g723(.A(new_n900), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n892), .A2(KEYINPUT54), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n910), .B1(new_n911), .B2(new_n873), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n709), .B1(new_n912), .B2(new_n905), .ZN(new_n913));
  INV_X1    g727(.A(new_n906), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n909), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT120), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n916), .A3(new_n885), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n908), .A2(new_n917), .ZN(G54));
  NAND4_X1  g732(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .A4(new_n421), .ZN(new_n919));
  INV_X1    g733(.A(new_n641), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n921), .A2(KEYINPUT121), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n921), .A2(KEYINPUT121), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n885), .B1(new_n919), .B2(new_n920), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(G60));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT59), .Z(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n617), .B1(new_n874), .B2(new_n928), .ZN(new_n929));
  AOI211_X1 g743(.A(new_n616), .B(new_n927), .C1(new_n911), .C2(new_n873), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n884), .A3(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT60), .Z(new_n933));
  AND2_X1   g747(.A1(new_n892), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n885), .B1(new_n934), .B2(new_n419), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n652), .B2(new_n934), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT61), .ZN(G66));
  AOI21_X1  g751(.A(new_n267), .B1(new_n592), .B2(G224), .ZN(new_n938));
  INV_X1    g752(.A(new_n842), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n852), .A2(new_n939), .A3(new_n854), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT122), .Z(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n938), .B1(new_n942), .B2(new_n267), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n353), .B1(G898), .B2(new_n267), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n943), .B(new_n944), .Z(G69));
  NAND2_X1  g759(.A1(new_n749), .A2(new_n859), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n688), .A2(new_n689), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT62), .ZN(new_n949));
  INV_X1    g763(.A(new_n670), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n840), .A2(new_n498), .A3(new_n950), .A4(new_n751), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n792), .A2(new_n801), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n267), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n529), .A2(new_n530), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n473), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT123), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n953), .A2(KEYINPUT123), .A3(new_n955), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n267), .B1(G227), .B2(G900), .ZN(new_n960));
  AOI22_X1  g774(.A1(new_n790), .A2(new_n791), .B1(new_n798), .B2(new_n800), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n781), .A2(new_n188), .A3(new_n669), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n728), .A2(new_n498), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n946), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n961), .A2(new_n267), .A3(new_n853), .A4(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n955), .B1(G900), .B2(G953), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n960), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n958), .A2(new_n959), .A3(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n965), .A2(new_n969), .A3(new_n966), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(new_n965), .B2(new_n966), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n972), .A2(new_n958), .A3(new_n959), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n973), .A2(new_n974), .A3(new_n960), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n973), .B2(new_n960), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n968), .B1(new_n975), .B2(new_n976), .ZN(G72));
  NAND2_X1  g791(.A1(G472), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT63), .Z(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT126), .Z(new_n980));
  OR2_X1    g794(.A1(new_n949), .A2(new_n952), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n980), .B1(new_n981), .B2(new_n942), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n982), .A2(new_n461), .A3(new_n675), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n961), .A2(new_n853), .A3(new_n964), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n980), .B1(new_n942), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n675), .A2(new_n461), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n884), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n986), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n866), .A2(new_n676), .A3(new_n979), .A4(new_n988), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n983), .A2(new_n987), .A3(new_n989), .ZN(G57));
endmodule


