//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n450, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(new_n461));
  INV_X1    g036(.A(new_n455), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n461), .B1(G2106), .B2(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n471), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT68), .Z(new_n486));
  AOI21_X1  g061(.A(G2105), .B1(new_n480), .B2(new_n481), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n478), .B(new_n486), .C1(G136), .C2(new_n487), .ZN(G162));
  NOR2_X1   g063(.A1(new_n464), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n492), .A2(new_n464), .A3(KEYINPUT4), .A4(G138), .ZN(new_n493));
  NAND2_X1  g068(.A1(G126), .A2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n495), .B2(new_n482), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(KEYINPUT69), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  OR2_X1    g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND3_X1   g082(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT6), .B1(KEYINPUT70), .B2(G651), .ZN(new_n509));
  INV_X1    g084(.A(new_n503), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI21_X1  g088(.A(G543), .B1(new_n508), .B2(new_n509), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n507), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND3_X1  g093(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(G51), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n519), .B(new_n521), .C1(new_n522), .C2(new_n514), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT70), .A2(G651), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n526), .A2(new_n527), .B1(new_n502), .B2(new_n503), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n528), .A2(G89), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n523), .A2(new_n529), .ZN(G168));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n510), .A2(new_n511), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(G651), .B1(new_n528), .B2(G90), .ZN(new_n535));
  INV_X1    g110(.A(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(new_n526), .B2(new_n527), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n535), .A2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n532), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n537), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n528), .A2(G81), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(KEYINPUT71), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n544), .A2(new_n549), .A3(new_n545), .A4(new_n546), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OAI211_X1 g134(.A(KEYINPUT72), .B(new_n558), .C1(new_n514), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n528), .A2(G91), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n502), .B2(new_n503), .ZN(new_n563));
  INV_X1    g138(.A(G78), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n536), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n558), .A2(KEYINPUT72), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n559), .B1(new_n568), .B2(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n537), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n560), .A2(new_n561), .A3(new_n566), .A4(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(KEYINPUT73), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(KEYINPUT73), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  NAND2_X1  g152(.A1(new_n528), .A2(G87), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n537), .A2(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(new_n504), .A2(G61), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(KEYINPUT74), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n582), .A2(KEYINPUT74), .B1(G73), .B2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n506), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  INV_X1    g161(.A(G48), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n512), .A2(new_n586), .B1(new_n514), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n506), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(KEYINPUT75), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(KEYINPUT75), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n528), .A2(G85), .B1(new_n537), .B2(G47), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n528), .A2(G92), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT10), .Z(new_n599));
  INV_X1    g174(.A(G79), .ZN(new_n600));
  OR3_X1    g175(.A1(new_n600), .A2(new_n536), .A3(KEYINPUT76), .ZN(new_n601));
  OAI21_X1  g176(.A(KEYINPUT76), .B1(new_n600), .B2(new_n536), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n601), .B(new_n602), .C1(new_n532), .C2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(G54), .B2(new_n537), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n597), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n597), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n575), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(new_n575), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n607), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n607), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n482), .A2(new_n472), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT77), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n623), .A2(G2100), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT78), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n487), .A2(G135), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n464), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(G123), .ZN(new_n629));
  OAI221_X1 g204(.A(new_n626), .B1(new_n627), .B2(new_n628), .C1(new_n629), .C2(new_n483), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2096), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n623), .B2(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n625), .A2(new_n632), .ZN(G156));
  XOR2_X1   g208(.A(G1341), .B(G1348), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT79), .ZN(new_n635));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n635), .B(new_n637), .Z(new_n638));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n638), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2067), .B(G2678), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT80), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT81), .B(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n652), .A2(new_n653), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n653), .B(KEYINPUT17), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n659), .B(new_n655), .C1(new_n652), .C2(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(new_n652), .A3(new_n654), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT82), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT20), .Z(new_n675));
  OR2_X1    g250(.A1(new_n668), .A2(new_n670), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n676), .A2(new_n673), .A3(new_n671), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n675), .B(new_n677), .C1(new_n673), .C2(new_n676), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G229));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G22), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT85), .Z(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G166), .B2(new_n685), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(G1971), .Z(new_n689));
  MUX2_X1   g264(.A(G23), .B(G288), .S(G16), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT33), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(G6), .A2(G16), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n589), .B2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT32), .B(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  OR3_X1    g272(.A1(new_n693), .A2(KEYINPUT34), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(KEYINPUT34), .B1(new_n693), .B2(new_n697), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n685), .A2(G24), .ZN(new_n700));
  INV_X1    g275(.A(G290), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n685), .ZN(new_n702));
  INV_X1    g277(.A(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n487), .A2(G131), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT84), .Z(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n707));
  INV_X1    g282(.A(G107), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G2105), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n484), .B2(G119), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G29), .ZN(new_n712));
  INV_X1    g287(.A(G25), .ZN(new_n713));
  OR3_X1    g288(.A1(new_n713), .A2(KEYINPUT83), .A3(G29), .ZN(new_n714));
  OAI21_X1  g289(.A(KEYINPUT83), .B1(new_n713), .B2(G29), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT35), .B(G1991), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n698), .A2(new_n699), .A3(new_n704), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT36), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n685), .A2(G19), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n552), .B2(new_n685), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1341), .ZN(new_n723));
  NOR2_X1   g298(.A1(G168), .A2(new_n685), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n685), .B2(G21), .ZN(new_n725));
  INV_X1    g300(.A(G1966), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT90), .ZN(new_n728));
  INV_X1    g303(.A(G29), .ZN(new_n729));
  OR3_X1    g304(.A1(new_n630), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n728), .B1(new_n630), .B2(new_n729), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G11), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n729), .B1(new_n734), .B2(G28), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(KEYINPUT91), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(KEYINPUT91), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n734), .B2(G28), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n733), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n730), .A2(new_n731), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n727), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n726), .B2(new_n725), .ZN(new_n742));
  INV_X1    g317(.A(G1961), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n685), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n685), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT92), .Z(new_n746));
  AOI211_X1 g321(.A(new_n723), .B(new_n742), .C1(new_n743), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n729), .A2(G35), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G162), .B2(new_n729), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT29), .B(G2090), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n607), .A2(new_n685), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G4), .B2(new_n685), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n751), .B1(G1348), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n729), .A2(G26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT28), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n487), .A2(G140), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n464), .A2(G116), .ZN(new_n759));
  OAI21_X1  g334(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n760));
  INV_X1    g335(.A(G128), .ZN(new_n761));
  OAI221_X1 g336(.A(new_n758), .B1(new_n759), .B2(new_n760), .C1(new_n761), .C2(new_n483), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT86), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n757), .B1(new_n765), .B2(new_n729), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT87), .B(G2067), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n754), .A2(G1348), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n767), .B2(new_n768), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT25), .Z(new_n772));
  INV_X1    g347(.A(new_n487), .ZN(new_n773));
  INV_X1    g348(.A(G139), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n482), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n772), .B1(new_n773), .B2(new_n774), .C1(new_n775), .C2(new_n464), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(G29), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n729), .A2(G33), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(new_n442), .ZN(new_n780));
  INV_X1    g355(.A(G2084), .ZN(new_n781));
  NAND2_X1  g356(.A1(G160), .A2(G29), .ZN(new_n782));
  INV_X1    g357(.A(G34), .ZN(new_n783));
  AOI21_X1  g358(.A(G29), .B1(new_n783), .B2(KEYINPUT24), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(KEYINPUT24), .B2(new_n783), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n780), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n484), .A2(G129), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n487), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n789));
  NAND3_X1  g364(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT26), .Z(new_n791));
  AND3_X1   g366(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n792), .A2(new_n729), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n729), .B2(G32), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT27), .B(G1996), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT88), .ZN(new_n796));
  OAI22_X1  g371(.A1(new_n794), .A2(new_n796), .B1(new_n779), .B2(new_n442), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n787), .A2(new_n797), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n794), .A2(new_n796), .B1(new_n781), .B2(new_n786), .ZN(new_n799));
  NOR2_X1   g374(.A1(G27), .A2(G29), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G164), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(new_n443), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n798), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n755), .A2(new_n770), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n746), .A2(new_n743), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT93), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n685), .A2(G20), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT23), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n575), .B2(new_n685), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1956), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n720), .A2(new_n747), .A3(new_n804), .A4(new_n811), .ZN(G150));
  INV_X1    g387(.A(G150), .ZN(G311));
  NOR2_X1   g388(.A1(new_n606), .A2(new_n613), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n528), .A2(G93), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n537), .A2(G55), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n817), .B(new_n818), .C1(new_n506), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n551), .A2(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n547), .A2(new_n820), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n816), .B(new_n824), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n826), .A2(new_n827), .A3(G860), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n820), .A2(G860), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT37), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n828), .A2(new_n830), .ZN(G145));
  XNOR2_X1  g406(.A(new_n764), .B(new_n500), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n792), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(new_n776), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n711), .B(new_n620), .ZN(new_n835));
  INV_X1    g410(.A(G130), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n464), .A2(G118), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n483), .A2(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G142), .B2(new_n487), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n835), .B(new_n840), .Z(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(KEYINPUT96), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n833), .A2(new_n776), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n834), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(G160), .B(KEYINPUT95), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n630), .ZN(new_n846));
  XNOR2_X1  g421(.A(G162), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n843), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n833), .A2(new_n776), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n841), .A2(KEYINPUT96), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n841), .A2(KEYINPUT96), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n844), .B(new_n847), .C1(new_n850), .C2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(G37), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n851), .B(new_n852), .C1(new_n848), .C2(new_n849), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n844), .ZN(new_n858));
  INV_X1    g433(.A(new_n847), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT97), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n861));
  AOI211_X1 g436(.A(new_n861), .B(new_n847), .C1(new_n857), .C2(new_n844), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n856), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g439(.A(new_n575), .B(new_n607), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n865), .A2(KEYINPUT41), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(KEYINPUT41), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n615), .B(new_n823), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OR3_X1    g445(.A1(new_n869), .A2(KEYINPUT98), .A3(new_n865), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT98), .B1(new_n869), .B2(new_n865), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT101), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(KEYINPUT101), .ZN(new_n875));
  XNOR2_X1  g450(.A(G303), .B(KEYINPUT99), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G305), .ZN(new_n877));
  XOR2_X1   g452(.A(G290), .B(G288), .Z(new_n878));
  OR2_X1    g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT42), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT100), .B1(new_n879), .B2(new_n880), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n879), .A2(KEYINPUT100), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n881), .B1(new_n885), .B2(KEYINPUT42), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n874), .A2(new_n875), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n886), .B1(new_n874), .B2(new_n875), .ZN(new_n888));
  OAI21_X1  g463(.A(G868), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G868), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n820), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(G295));
  NAND2_X1  g467(.A1(new_n889), .A2(new_n891), .ZN(G331));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n894));
  AOI21_X1  g469(.A(G168), .B1(G301), .B2(KEYINPUT102), .ZN(new_n895));
  NOR2_X1   g470(.A1(G301), .A2(KEYINPUT102), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n895), .B(new_n896), .Z(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n823), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n898), .A2(new_n865), .ZN(new_n899));
  INV_X1    g474(.A(new_n868), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n897), .B(new_n824), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n855), .B1(new_n902), .B2(new_n885), .ZN(new_n903));
  INV_X1    g478(.A(new_n884), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n901), .B1(new_n867), .B2(new_n866), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n898), .A2(new_n865), .ZN(new_n906));
  OAI22_X1  g481(.A1(new_n904), .A2(new_n882), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n894), .B1(new_n903), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n904), .A2(new_n882), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n905), .A2(new_n906), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n907), .A2(KEYINPUT103), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n914), .B1(new_n902), .B2(new_n885), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n912), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n909), .B1(new_n916), .B2(new_n894), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT44), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n912), .B(new_n894), .C1(new_n913), .C2(new_n915), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n903), .B2(new_n908), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(new_n923), .ZN(G397));
  INV_X1    g499(.A(G2067), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n764), .B(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G1996), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n926), .B1(new_n927), .B2(new_n792), .ZN(new_n928));
  INV_X1    g503(.A(G1384), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n489), .A2(new_n490), .ZN(new_n930));
  INV_X1    g505(.A(new_n494), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n498), .A2(KEYINPUT69), .ZN(new_n932));
  INV_X1    g507(.A(G138), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n933), .A2(G2105), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n931), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n465), .A2(new_n466), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n930), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n932), .B1(new_n487), .B2(G138), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n929), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G125), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n480), .B2(new_n481), .ZN(new_n943));
  INV_X1    g518(.A(new_n468), .ZN(new_n944));
  OAI21_X1  g519(.A(G2105), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n945), .A2(G40), .A3(new_n473), .A4(new_n470), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT104), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n927), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n928), .A2(new_n948), .B1(new_n792), .B2(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n706), .A2(new_n717), .A3(new_n710), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(G2067), .B2(new_n764), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n954), .A2(KEYINPUT124), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(KEYINPUT124), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n948), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n950), .A2(KEYINPUT46), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT125), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n926), .A2(new_n792), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n948), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n959), .B(new_n961), .C1(KEYINPUT46), .C2(new_n950), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n962), .A2(KEYINPUT47), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(KEYINPUT47), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n717), .B1(new_n706), .B2(new_n710), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n948), .B1(new_n965), .B2(new_n952), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n951), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(G290), .A2(G1986), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n947), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(KEYINPUT126), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT48), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n963), .A2(new_n964), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n957), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT127), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT127), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n957), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1956), .ZN(new_n978));
  INV_X1    g553(.A(G40), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n469), .A2(new_n474), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n496), .B2(new_n499), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n939), .A2(KEYINPUT50), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n978), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI22_X1  g560(.A1(new_n532), .A2(new_n562), .B1(new_n564), .B2(new_n536), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n986), .A2(G651), .B1(new_n528), .B2(G91), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT57), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n987), .A2(new_n988), .A3(new_n570), .A4(new_n560), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n571), .A2(KEYINPUT57), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(KEYINPUT45), .B(new_n929), .C1(new_n937), .C2(new_n938), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT56), .B(G2072), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n941), .A2(new_n980), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n985), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n991), .B1(new_n985), .B2(new_n994), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT61), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n985), .A2(new_n994), .ZN(new_n998));
  INV_X1    g573(.A(new_n991), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT61), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n985), .A2(new_n991), .A3(new_n994), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n997), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n941), .A2(new_n927), .A3(new_n980), .A4(new_n992), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n980), .A2(new_n981), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT58), .B(G1341), .Z(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1005), .B1(new_n1010), .B2(new_n552), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1005), .A3(new_n552), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(KEYINPUT59), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT59), .ZN(new_n1015));
  AOI211_X1 g590(.A(KEYINPUT116), .B(new_n551), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n1011), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1004), .A2(new_n1014), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1004), .A2(KEYINPUT117), .A3(new_n1014), .A4(new_n1017), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT106), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1022), .B1(new_n981), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n939), .A2(KEYINPUT106), .A3(KEYINPUT50), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n981), .A2(new_n982), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n980), .ZN(new_n1027));
  INV_X1    g602(.A(G1348), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1007), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1027), .A2(new_n1028), .B1(new_n925), .B2(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1030), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n606), .B1(new_n1030), .B2(KEYINPUT60), .ZN(new_n1032));
  OAI22_X1  g607(.A1(new_n1031), .A2(new_n1032), .B1(KEYINPUT60), .B2(new_n1030), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1020), .A2(new_n1021), .A3(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1030), .A2(new_n606), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1002), .B1(new_n1035), .B2(new_n996), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT113), .B(G2084), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n946), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1023), .B1(new_n500), .B2(new_n929), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1043), .A2(KEYINPUT106), .B1(new_n981), .B2(new_n982), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1044), .A2(KEYINPUT114), .A3(new_n1024), .A4(new_n1039), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n992), .A2(KEYINPUT112), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n981), .A2(new_n1047), .A3(KEYINPUT45), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n980), .B1(new_n981), .B2(KEYINPUT45), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT111), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1052), .B(new_n980), .C1(new_n981), .C2(KEYINPUT45), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1049), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1042), .B(new_n1045), .C1(new_n1054), .C2(G1966), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G8), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n1057));
  NAND2_X1  g632(.A1(G286), .A2(G8), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT118), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1056), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT51), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1059), .B1(new_n1055), .B2(G8), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1061), .B(new_n1062), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1057), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1068));
  INV_X1    g643(.A(G8), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n992), .A2(KEYINPUT112), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1047), .B1(new_n981), .B2(KEYINPUT45), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1052), .B1(new_n941), .B2(new_n980), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1053), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AND4_X1   g650(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1039), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1075), .A2(new_n726), .B1(KEYINPUT114), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1069), .B1(new_n1077), .B2(new_n1042), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1068), .B1(new_n1078), .B2(new_n1059), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1062), .B1(new_n1079), .B2(new_n1061), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1067), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(G2078), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1054), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1027), .A2(new_n743), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n941), .A2(new_n980), .A3(new_n992), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1083), .B1(new_n1089), .B2(G2078), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1086), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1091), .A2(G171), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1089), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(KEYINPUT53), .A3(new_n443), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1090), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1027), .A2(KEYINPUT121), .A3(new_n743), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1087), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1096), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT54), .B1(new_n1100), .B2(G301), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1082), .B1(new_n1093), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1099), .A2(new_n1097), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1104), .A2(new_n1090), .A3(new_n1095), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1103), .B1(new_n1105), .B2(G171), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT120), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(new_n1090), .A3(new_n1088), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1106), .B(KEYINPUT122), .C1(G171), .C2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1102), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1029), .A2(new_n1069), .ZN(new_n1112));
  INV_X1    g687(.A(G1976), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT52), .B1(G288), .B2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1112), .B(new_n1114), .C1(new_n1113), .C2(G288), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1112), .B1(new_n1113), .B2(G288), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1115), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(G1981), .B1(new_n585), .B2(KEYINPUT109), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(new_n589), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT49), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1112), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1119), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(KEYINPUT108), .A2(KEYINPUT55), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(G166), .B2(new_n1069), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT108), .B(KEYINPUT55), .ZN(new_n1129));
  NAND3_X1  g704(.A1(G303), .A2(G8), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1027), .A2(G2090), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1132), .A2(KEYINPUT107), .B1(G1971), .B2(new_n1094), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1132), .A2(KEYINPUT107), .ZN(new_n1134));
  OAI211_X1 g709(.A(G8), .B(new_n1131), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1094), .A2(G1971), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n983), .A2(new_n984), .A3(G2090), .ZN(new_n1137));
  OAI21_X1  g712(.A(G8), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1131), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1126), .A2(new_n1135), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(G171), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1100), .A2(G301), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1141), .B1(new_n1144), .B2(new_n1103), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1037), .A2(new_n1081), .A3(new_n1111), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1067), .B2(new_n1080), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1061), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT119), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1150), .A2(KEYINPUT62), .A3(new_n1066), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1148), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1126), .ZN(new_n1154));
  NOR2_X1   g729(.A1(G305), .A2(G1981), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1156));
  NOR2_X1   g731(.A1(G288), .A2(G1976), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n1112), .B(KEYINPUT110), .Z(new_n1159));
  OAI22_X1  g734(.A1(new_n1154), .A2(new_n1135), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  XOR2_X1   g735(.A(KEYINPUT115), .B(KEYINPUT63), .Z(new_n1161));
  NAND2_X1  g736(.A1(new_n1078), .A2(G168), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1161), .B1(new_n1141), .B2(new_n1162), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1078), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1164));
  OAI21_X1  g739(.A(G8), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1139), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1164), .A2(new_n1166), .A3(new_n1135), .A4(new_n1126), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1160), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1146), .A2(new_n1153), .A3(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n701), .A2(new_n703), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n947), .B1(new_n1170), .B2(new_n968), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n967), .A2(new_n1171), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1169), .A2(KEYINPUT123), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(KEYINPUT123), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n977), .B1(new_n1173), .B2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g750(.A1(new_n649), .A2(new_n665), .A3(G319), .ZN(new_n1177));
  NOR2_X1   g751(.A1(G229), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g752(.A1(new_n921), .A2(new_n863), .A3(new_n1178), .ZN(G225));
  INV_X1    g753(.A(G225), .ZN(G308));
endmodule


