//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948;
  INV_X1    g000(.A(G141gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G148gat), .ZN(new_n203));
  INV_X1    g002(.A(G148gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G141gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT2), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n206), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(KEYINPUT80), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT80), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(G155gat), .A3(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT79), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G155gat), .B2(G162gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n213), .A2(new_n218), .A3(new_n215), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n211), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n212), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n225));
  AND2_X1   g024(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n225), .B1(new_n228), .B2(G204gat), .ZN(new_n229));
  INV_X1    g028(.A(G211gat), .ZN(new_n230));
  INV_X1    g029(.A(G218gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G211gat), .A2(G218gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G204gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(new_n226), .B2(new_n227), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n229), .A2(KEYINPUT77), .A3(new_n234), .A4(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT74), .ZN(new_n238));
  INV_X1    g037(.A(G197gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(G204gat), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n225), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n236), .A2(new_n242), .A3(new_n234), .A4(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT77), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n237), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n233), .ZN(new_n248));
  NOR2_X1   g047(.A1(G211gat), .A2(G218gat), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT75), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT75), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n232), .A2(new_n251), .A3(new_n233), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n242), .A3(new_n243), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n253), .A2(KEYINPUT76), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT76), .B1(new_n253), .B2(new_n254), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n247), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT87), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n258), .B1(new_n257), .B2(new_n259), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n224), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G228gat), .A2(G233gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT82), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n213), .A2(new_n218), .A3(new_n215), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n218), .B1(new_n213), .B2(new_n215), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n223), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n203), .A2(new_n205), .B1(KEYINPUT2), .B2(new_n210), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n209), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(KEYINPUT81), .B(KEYINPUT3), .Z(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n266), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  AOI211_X1 g074(.A(KEYINPUT82), .B(new_n273), .C1(new_n269), .C2(new_n271), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n259), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n257), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n265), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n270), .B1(new_n220), .B2(new_n221), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n281), .A2(KEYINPUT83), .A3(new_n212), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT83), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n283), .B1(new_n269), .B2(new_n271), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n234), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n237), .A2(new_n246), .B1(new_n286), .B2(new_n254), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n274), .B1(new_n287), .B2(KEYINPUT29), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n277), .A2(new_n278), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n265), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n289), .A2(KEYINPUT86), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT86), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n254), .A2(new_n286), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT29), .B1(new_n247), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n285), .B1(new_n294), .B2(new_n273), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT82), .B1(new_n224), .B2(new_n273), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n272), .A2(new_n266), .A3(new_n274), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT29), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n295), .B1(new_n298), .B2(new_n257), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n292), .B1(new_n299), .B2(new_n265), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n280), .B1(new_n291), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G22gat), .ZN(new_n302));
  INV_X1    g101(.A(G22gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n280), .B(new_n303), .C1(new_n291), .C2(new_n300), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G78gat), .B(G106gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT31), .B(G50gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT85), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT89), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT86), .B1(new_n289), .B2(new_n290), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n299), .A2(new_n292), .A3(new_n265), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n313), .A2(new_n314), .B1(new_n264), .B2(new_n279), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(KEYINPUT89), .A3(new_n303), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT88), .B1(new_n315), .B2(new_n303), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT88), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n319), .A3(G22gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n320), .A3(new_n308), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n310), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT28), .ZN(new_n323));
  INV_X1    g122(.A(G190gat), .ZN(new_n324));
  AND2_X1   g123(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n323), .B(new_n324), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G183gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(new_n324), .ZN(new_n329));
  INV_X1    g128(.A(G169gat), .ZN(new_n330));
  INV_X1    g129(.A(G176gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n331), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT26), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT26), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT27), .B(G183gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n323), .B1(new_n338), .B2(new_n324), .ZN(new_n339));
  NOR3_X1   g138(.A1(new_n329), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT65), .ZN(new_n341));
  NAND3_X1  g140(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(G183gat), .B2(G190gat), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n341), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n344), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n324), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT65), .A4(new_n342), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT66), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(G176gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n331), .A2(KEYINPUT66), .ZN(new_n351));
  OAI211_X1 g150(.A(KEYINPUT23), .B(new_n330), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n332), .B1(new_n353), .B2(new_n333), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n345), .A2(new_n348), .A3(new_n352), .A4(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT23), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n358), .A2(KEYINPUT25), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(KEYINPUT67), .A2(G183gat), .A3(G190gat), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT24), .B1(new_n361), .B2(KEYINPUT68), .ZN(new_n362));
  NAND2_X1  g161(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n363), .A2(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n347), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n340), .B1(new_n357), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT1), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n368), .B1(G113gat), .B2(G120gat), .ZN(new_n369));
  XOR2_X1   g168(.A(KEYINPUT71), .B(G113gat), .Z(new_n370));
  AOI21_X1  g169(.A(new_n369), .B1(new_n370), .B2(G120gat), .ZN(new_n371));
  INV_X1    g170(.A(G134gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G127gat), .ZN(new_n373));
  INV_X1    g172(.A(G127gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G134gat), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT72), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n375), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT72), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n371), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT69), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(new_n372), .A3(G127gat), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT69), .B1(new_n374), .B2(G134gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n372), .A2(G127gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT70), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n369), .B1(G113gat), .B2(G120gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT70), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n389), .B(new_n382), .C1(new_n383), .C2(new_n384), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n380), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n367), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n355), .A2(new_n356), .B1(new_n360), .B2(new_n365), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n392), .B1(new_n395), .B2(new_n340), .ZN(new_n396));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n394), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(KEYINPUT34), .ZN(new_n399));
  XOR2_X1   g198(.A(G15gat), .B(G43gat), .Z(new_n400));
  XNOR2_X1  g199(.A(G71gat), .B(G99gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n397), .B1(new_n394), .B2(new_n396), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(KEYINPUT33), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT32), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n394), .A2(new_n396), .ZN(new_n408));
  INV_X1    g207(.A(new_n397), .ZN(new_n409));
  AOI221_X4 g208(.A(new_n405), .B1(KEYINPUT33), .B2(new_n402), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n399), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT73), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n367), .A2(new_n393), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n395), .A2(new_n392), .A3(new_n340), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n409), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT32), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n418), .A3(new_n402), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n406), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT34), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n398), .B(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n411), .A2(new_n412), .A3(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(KEYINPUT73), .B(new_n399), .C1(new_n407), .C2(new_n410), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(G226gat), .A2(G233gat), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n367), .B2(KEYINPUT29), .ZN(new_n428));
  OAI211_X1 g227(.A(G226gat), .B(G233gat), .C1(new_n395), .C2(new_n340), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n278), .ZN(new_n431));
  XNOR2_X1  g230(.A(G8gat), .B(G36gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(G64gat), .B(G92gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n428), .A2(new_n257), .A3(new_n429), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n431), .A2(KEYINPUT30), .A3(new_n436), .A4(new_n435), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n428), .A2(new_n257), .A3(new_n429), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n257), .B1(new_n428), .B2(new_n429), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n441), .B1(new_n444), .B2(new_n435), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT78), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n440), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449));
  INV_X1    g248(.A(G85gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT0), .B(G57gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n451), .B(new_n452), .Z(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n224), .A2(KEYINPUT3), .B1(new_n380), .B2(new_n391), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n455), .B1(new_n275), .B2(new_n276), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n393), .B(KEYINPUT4), .C1(new_n282), .C2(new_n284), .ZN(new_n457));
  NAND2_X1  g256(.A1(G225gat), .A2(G233gat), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n272), .A2(new_n380), .A3(new_n391), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT4), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n456), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n392), .A2(new_n224), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n460), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n392), .A2(KEYINPUT84), .A3(new_n224), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n459), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n463), .A2(KEYINPUT5), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n296), .A2(new_n297), .ZN(new_n470));
  INV_X1    g269(.A(new_n460), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n470), .A2(new_n455), .B1(new_n471), .B2(KEYINPUT4), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n461), .B1(new_n285), .B2(new_n392), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n459), .A2(KEYINPUT5), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n454), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT6), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n469), .A2(new_n475), .A3(new_n454), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n477), .B1(new_n480), .B2(new_n476), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n445), .A2(KEYINPUT78), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n448), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n322), .A2(new_n426), .A3(new_n483), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n484), .A2(KEYINPUT35), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n478), .A2(new_n479), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n476), .A2(KEYINPUT92), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT92), .ZN(new_n488));
  AOI211_X1 g287(.A(new_n488), .B(new_n454), .C1(new_n469), .C2(new_n475), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n486), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n477), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n439), .B(new_n441), .C1(new_n435), .C2(new_n444), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT93), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(KEYINPUT93), .A3(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n411), .A2(new_n423), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n322), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n322), .A2(KEYINPUT90), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT90), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n504), .B(new_n310), .C1(new_n317), .C2(new_n321), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n483), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n426), .A2(KEYINPUT36), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT36), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n499), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n309), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n511), .B1(new_n302), .B2(new_n304), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n318), .A2(new_n308), .A3(new_n320), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n312), .A2(new_n316), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT37), .B1(new_n442), .B2(new_n443), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT37), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n431), .A2(new_n517), .A3(new_n436), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT38), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n516), .A2(new_n518), .A3(new_n519), .A4(new_n434), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n520), .A2(new_n437), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(new_n518), .A3(new_n434), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT38), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n490), .A2(new_n521), .A3(new_n477), .A4(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n476), .B(KEYINPUT92), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n472), .A2(new_n473), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n459), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n466), .A2(new_n467), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n528), .B(KEYINPUT39), .C1(new_n529), .C2(new_n459), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT39), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT91), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n527), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n458), .B1(new_n472), .B2(new_n473), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n453), .B1(new_n535), .B2(new_n532), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT40), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n534), .A2(new_n536), .A3(KEYINPUT40), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n525), .A2(new_n539), .A3(new_n492), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n510), .B1(new_n515), .B2(new_n542), .ZN(new_n543));
  OAI22_X1  g342(.A1(new_n485), .A2(new_n502), .B1(new_n506), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT95), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(KEYINPUT96), .ZN(new_n548));
  OAI22_X1  g347(.A1(new_n548), .A2(G1gat), .B1(KEYINPUT16), .B2(new_n547), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n548), .A2(G1gat), .ZN(new_n550));
  OR3_X1    g349(.A1(new_n549), .A2(new_n550), .A3(G8gat), .ZN(new_n551));
  OAI21_X1  g350(.A(G8gat), .B1(new_n549), .B2(new_n550), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OR3_X1    g352(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n554), .A2(new_n555), .B1(G29gat), .B2(G36gat), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n556), .A2(KEYINPUT15), .ZN(new_n557));
  XNOR2_X1  g356(.A(G43gat), .B(G50gat), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n556), .A2(KEYINPUT15), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n553), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT13), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n562), .B(KEYINPUT17), .Z(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(new_n552), .A3(new_n551), .ZN(new_n568));
  INV_X1    g367(.A(new_n562), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n568), .A2(KEYINPUT18), .A3(new_n570), .A4(new_n564), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n564), .A3(new_n570), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT18), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n566), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(G197gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT11), .B(G169gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(KEYINPUT94), .B(KEYINPUT12), .Z(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n581), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n566), .A2(new_n574), .A3(new_n583), .A4(new_n571), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G57gat), .B(G64gat), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT97), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G71gat), .B(G78gat), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n590), .B(KEYINPUT98), .Z(new_n594));
  OAI21_X1  g393(.A(new_n593), .B1(new_n594), .B2(new_n592), .ZN(new_n595));
  MUX2_X1   g394(.A(new_n595), .B(new_n593), .S(new_n553), .Z(new_n596));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(new_n328), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G211gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n596), .B(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G127gat), .B(G155gat), .Z(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  OR2_X1    g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n600), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n607), .B1(new_n450), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT99), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT7), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G99gat), .B(G106gat), .Z(new_n614));
  OR2_X1    g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT100), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n613), .A2(new_n614), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n567), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n616), .B(new_n617), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n569), .ZN(new_n621));
  XOR2_X1   g420(.A(G190gat), .B(G218gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT101), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n623), .A2(KEYINPUT102), .ZN(new_n624));
  AND2_X1   g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n624), .B1(KEYINPUT41), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n619), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n623), .A2(KEYINPUT102), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n627), .A2(new_n628), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n632), .B1(new_n629), .B2(new_n633), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n606), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(G230gat), .ZN(new_n639));
  INV_X1    g438(.A(G233gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT104), .B(KEYINPUT10), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n620), .A2(new_n591), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n615), .A2(KEYINPUT103), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n645), .A2(new_n617), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n617), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(new_n590), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n643), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n618), .A2(new_n650), .A3(new_n594), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n642), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n644), .A2(new_n648), .A3(new_n641), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(G176gat), .B(G204gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT105), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n652), .A2(new_n653), .A3(new_n658), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n638), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n544), .A2(new_n585), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n481), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g466(.A1(new_n664), .A2(new_n492), .ZN(new_n668));
  INV_X1    g467(.A(G8gat), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT42), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT106), .B(KEYINPUT16), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G8gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  MUX2_X1   g472(.A(KEYINPUT42), .B(new_n670), .S(new_n673), .Z(G1325gat));
  INV_X1    g473(.A(new_n499), .ZN(new_n675));
  AOI21_X1  g474(.A(G15gat), .B1(new_n664), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n510), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n677), .A2(G15gat), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n676), .B1(new_n664), .B2(new_n678), .ZN(G1326gat));
  NAND2_X1  g478(.A1(new_n503), .A2(new_n505), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  INV_X1    g482(.A(new_n483), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n543), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n484), .A2(KEYINPUT35), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(new_n498), .B2(new_n501), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n637), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n606), .ZN(new_n691));
  INV_X1    g490(.A(new_n585), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n662), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n690), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(G29gat), .A3(new_n481), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT45), .Z(new_n696));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n543), .B1(new_n680), .B2(new_n684), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n322), .A2(new_n500), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT93), .B1(new_n491), .B2(new_n493), .ZN(new_n700));
  AOI211_X1 g499(.A(new_n495), .B(new_n492), .C1(new_n490), .C2(new_n477), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI22_X1  g501(.A1(new_n699), .A2(new_n702), .B1(new_n484), .B2(KEYINPUT35), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n697), .B(new_n636), .C1(new_n698), .C2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT44), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n544), .A2(new_n697), .A3(new_n706), .A4(new_n636), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n691), .A3(new_n693), .ZN(new_n709));
  OAI21_X1  g508(.A(G29gat), .B1(new_n709), .B2(new_n481), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n696), .A2(new_n710), .ZN(G1328gat));
  NOR3_X1   g510(.A1(new_n694), .A2(G36gat), .A3(new_n493), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT46), .ZN(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n709), .B2(new_n493), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1329gat));
  INV_X1    g514(.A(G43gat), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n709), .A2(new_n716), .A3(new_n510), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n694), .B2(new_n499), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n717), .B2(new_n718), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(G1330gat));
  NAND4_X1  g521(.A1(new_n708), .A2(new_n680), .A3(new_n691), .A4(new_n693), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G50gat), .ZN(new_n724));
  INV_X1    g523(.A(new_n680), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n694), .A2(G50gat), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT109), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n726), .B1(new_n723), .B2(G50gat), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n731), .A2(new_n732), .A3(KEYINPUT48), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n708), .A2(new_n515), .A3(new_n691), .A4(new_n693), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G50gat), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n726), .A2(new_n729), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n736), .A2(new_n737), .A3(new_n734), .ZN(new_n739));
  OAI22_X1  g538(.A1(new_n730), .A2(new_n733), .B1(new_n738), .B2(new_n739), .ZN(G1331gat));
  NAND2_X1  g539(.A1(new_n692), .A2(new_n662), .ZN(new_n741));
  AOI211_X1 g540(.A(new_n638), .B(new_n741), .C1(new_n687), .C2(new_n689), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n481), .B(KEYINPUT111), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G57gat), .ZN(G1332gat));
  INV_X1    g544(.A(new_n742), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n493), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  AND2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n747), .B2(new_n748), .ZN(G1333gat));
  NAND3_X1  g550(.A1(new_n742), .A2(G71gat), .A3(new_n677), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n746), .A2(new_n499), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(G71gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n742), .A2(new_n680), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  INV_X1    g556(.A(new_n662), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n544), .A2(new_n691), .A3(new_n636), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(new_n585), .ZN(new_n763));
  INV_X1    g562(.A(new_n761), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n690), .A2(new_n692), .A3(new_n691), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n759), .A2(new_n760), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n758), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n450), .A3(new_n665), .ZN(new_n769));
  INV_X1    g568(.A(new_n741), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n708), .A2(new_n691), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(G85gat), .B1(new_n771), .B2(new_n481), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(G1336gat));
  NOR2_X1   g572(.A1(new_n493), .A2(G92gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(G92gat), .B1(new_n771), .B2(new_n493), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n777), .B1(new_n775), .B2(new_n778), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(G1337gat));
  INV_X1    g580(.A(G99gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n768), .A2(new_n782), .A3(new_n675), .ZN(new_n783));
  OAI21_X1  g582(.A(G99gat), .B1(new_n771), .B2(new_n510), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1338gat));
  OR2_X1    g584(.A1(new_n322), .A2(G106gat), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n768), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(G106gat), .B1(new_n771), .B2(new_n322), .ZN(new_n789));
  XOR2_X1   g588(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n790));
  NAND3_X1  g589(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n708), .A2(new_n680), .A3(new_n691), .A4(new_n770), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n768), .A2(new_n787), .B1(G106gat), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n791), .B1(new_n792), .B2(new_n794), .ZN(G1339gat));
  OR2_X1    g594(.A1(new_n652), .A2(KEYINPUT54), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n644), .A2(new_n648), .ZN(new_n797));
  INV_X1    g596(.A(new_n643), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OR3_X1    g598(.A1(new_n618), .A2(new_n650), .A3(new_n594), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n800), .A3(new_n641), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n801), .A2(KEYINPUT54), .A3(new_n652), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n796), .A2(new_n659), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n796), .A2(new_n802), .A3(KEYINPUT55), .A4(new_n659), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n805), .A2(new_n585), .A3(new_n661), .A4(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n584), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n564), .B1(new_n568), .B2(new_n570), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n809), .A2(new_n810), .B1(new_n563), .B2(new_n565), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n579), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n636), .B1(new_n814), .B2(new_n662), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n606), .B1(new_n807), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n805), .A2(new_n814), .A3(new_n661), .A4(new_n806), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n636), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n816), .A2(new_n818), .B1(new_n663), .B2(new_n692), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n819), .A2(new_n499), .A3(new_n680), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n481), .A2(new_n492), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G113gat), .B1(new_n822), .B2(new_n692), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT116), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n815), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n818), .A3(new_n691), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n663), .A2(new_n692), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n743), .A2(new_n493), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n322), .A2(new_n426), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n692), .A2(new_n370), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n824), .B1(new_n833), .B2(new_n834), .ZN(G1340gat));
  OAI21_X1  g634(.A(G120gat), .B1(new_n822), .B2(new_n758), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n758), .A2(G120gat), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n833), .B2(new_n837), .ZN(G1341gat));
  NAND4_X1  g637(.A1(new_n820), .A2(G127gat), .A3(new_n606), .A4(new_n821), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n839), .A2(KEYINPUT117), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n374), .B1(new_n833), .B2(new_n691), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(KEYINPUT117), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(G1342gat));
  NAND4_X1  g642(.A1(new_n831), .A2(new_n372), .A3(new_n832), .A4(new_n636), .ZN(new_n844));
  XOR2_X1   g643(.A(new_n844), .B(KEYINPUT56), .Z(new_n845));
  OAI21_X1  g644(.A(G134gat), .B1(new_n822), .B2(new_n637), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n845), .A2(new_n848), .A3(new_n849), .ZN(G1343gat));
  NAND2_X1  g649(.A1(new_n510), .A2(new_n821), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n322), .B1(new_n826), .B2(new_n827), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT57), .B1(new_n819), .B2(new_n725), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n585), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT119), .B1(new_n856), .B2(G141gat), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n677), .A2(new_n322), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n585), .A2(new_n202), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n830), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n861), .B1(new_n856), .B2(G141gat), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n857), .A2(new_n862), .A3(KEYINPUT58), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864));
  AOI221_X4 g663(.A(new_n861), .B1(KEYINPUT119), .B2(new_n864), .C1(new_n856), .C2(G141gat), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n863), .A2(new_n865), .ZN(G1344gat));
  NOR2_X1   g665(.A1(new_n830), .A2(new_n859), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n204), .A3(new_n662), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT57), .B1(new_n819), .B2(new_n322), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n828), .A2(new_n853), .A3(new_n680), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n872), .A2(new_n510), .A3(new_n662), .A4(new_n821), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n869), .B1(new_n873), .B2(G148gat), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n854), .A2(new_n855), .ZN(new_n875));
  AOI211_X1 g674(.A(KEYINPUT59), .B(new_n204), .C1(new_n875), .C2(new_n662), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n868), .B1(new_n874), .B2(new_n876), .ZN(G1345gat));
  AOI21_X1  g676(.A(KEYINPUT120), .B1(new_n867), .B2(new_n606), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(G155gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n867), .A2(KEYINPUT120), .A3(new_n606), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n606), .A2(G155gat), .ZN(new_n881));
  AOI22_X1  g680(.A1(new_n879), .A2(new_n880), .B1(new_n875), .B2(new_n881), .ZN(G1346gat));
  INV_X1    g681(.A(G162gat), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n883), .A3(new_n636), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n875), .A2(new_n636), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n883), .ZN(G1347gat));
  NOR3_X1   g685(.A1(new_n819), .A2(new_n665), .A3(new_n493), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n887), .A2(new_n832), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n330), .A3(new_n585), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n743), .A2(new_n493), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n820), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n692), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n889), .B1(new_n330), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT122), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n889), .B(new_n900), .C1(new_n330), .C2(new_n897), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1348gat));
  AOI21_X1  g701(.A(G176gat), .B1(new_n888), .B2(new_n662), .ZN(new_n903));
  INV_X1    g702(.A(new_n896), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n758), .A2(new_n350), .A3(new_n351), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(G1349gat));
  NAND3_X1  g705(.A1(new_n888), .A2(new_n338), .A3(new_n606), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n896), .A2(new_n691), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n328), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT60), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n907), .B(new_n911), .C1(new_n328), .C2(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1350gat));
  NAND3_X1  g712(.A1(new_n888), .A2(new_n324), .A3(new_n636), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n914), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G190gat), .B1(new_n896), .B2(new_n637), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT61), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1351gat));
  NAND3_X1  g718(.A1(new_n892), .A2(new_n510), .A3(new_n893), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n921), .A2(KEYINPUT124), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(KEYINPUT124), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n870), .A2(new_n871), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(G197gat), .B1(new_n924), .B2(new_n692), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n887), .A2(new_n858), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n239), .A3(new_n585), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1352gat));
  NOR2_X1   g727(.A1(new_n665), .A2(new_n493), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n758), .A2(G204gat), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n828), .A2(new_n858), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n931), .B(KEYINPUT62), .Z(new_n932));
  OAI21_X1  g731(.A(G204gat), .B1(new_n924), .B2(new_n758), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT125), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n932), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(G1353gat));
  NAND3_X1  g737(.A1(new_n926), .A2(new_n230), .A3(new_n606), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n872), .A2(new_n606), .A3(new_n921), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n940), .B2(G211gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1354gat));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n637), .B1(new_n924), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n945), .B1(new_n944), .B2(new_n924), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G218gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n926), .A2(new_n231), .A3(new_n636), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1355gat));
endmodule


