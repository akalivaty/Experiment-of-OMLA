//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT83), .Z(new_n203));
  XOR2_X1   g002(.A(G141gat), .B(G148gat), .Z(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n204), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G141gat), .B(G148gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n208), .B(new_n207), .C1(new_n212), .C2(KEYINPUT2), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT82), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT82), .B1(new_n211), .B2(new_n213), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217));
  XNOR2_X1  g016(.A(G211gat), .B(G218gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G218gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT76), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT76), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G218gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT22), .B1(new_n224), .B2(G211gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(G197gat), .B(G204gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n219), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G211gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n229), .B1(new_n221), .B2(new_n223), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n218), .B(new_n226), .C1(new_n230), .C2(KEYINPUT22), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT29), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT84), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n217), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI211_X1 g033(.A(KEYINPUT84), .B(KEYINPUT29), .C1(new_n228), .C2(new_n231), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n216), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n211), .A2(new_n213), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n217), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT29), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT77), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n228), .A2(new_n241), .A3(new_n231), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT22), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT76), .B(G218gat), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n243), .B1(new_n244), .B2(new_n229), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n218), .B1(new_n245), .B2(new_n226), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT77), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n239), .A2(new_n240), .B1(new_n242), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n203), .B1(new_n236), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n242), .A2(new_n240), .A3(new_n247), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n238), .B1(new_n251), .B2(new_n217), .ZN(new_n252));
  NOR3_X1   g051(.A1(new_n252), .A2(new_n248), .A3(new_n202), .ZN(new_n253));
  OAI21_X1  g052(.A(G22gat), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT85), .ZN(new_n255));
  XNOR2_X1  g054(.A(G78gat), .B(G106gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT31), .B(G50gat), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n256), .B(new_n257), .Z(new_n258));
  NOR2_X1   g057(.A1(new_n248), .A2(new_n202), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n251), .A2(new_n217), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n237), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G22gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n231), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n240), .B1(new_n264), .B2(new_n246), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT84), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n232), .A2(new_n233), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n267), .A3(new_n217), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n248), .B1(new_n268), .B2(new_n216), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n262), .B(new_n263), .C1(new_n269), .C2(new_n203), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n255), .A2(new_n258), .B1(new_n254), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT85), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n254), .A2(new_n270), .A3(new_n272), .A4(new_n258), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G1gat), .B(G29gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT0), .ZN(new_n277));
  XNOR2_X1  g076(.A(G57gat), .B(G85gat), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n277), .B(new_n278), .Z(new_n279));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n280));
  INV_X1    g079(.A(G127gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G134gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n281), .A2(KEYINPUT71), .A3(G134gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT70), .B(G134gat), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n284), .B(new_n285), .C1(new_n286), .C2(new_n281), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n288));
  INV_X1    g087(.A(G113gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(G120gat), .ZN(new_n290));
  INV_X1    g089(.A(G120gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(G113gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n288), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n289), .B2(G120gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n291), .A2(KEYINPUT72), .A3(G113gat), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n296), .B(new_n297), .C1(G113gat), .C2(new_n291), .ZN(new_n298));
  INV_X1    g097(.A(G134gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G127gat), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n282), .A2(new_n300), .A3(new_n288), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n294), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n237), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n287), .A2(new_n293), .B1(new_n301), .B2(new_n298), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n238), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n280), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n305), .B1(KEYINPUT3), .B2(new_n237), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n239), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n308), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n305), .B1(new_n214), .B2(new_n215), .ZN(new_n314));
  XOR2_X1   g113(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n303), .A2(new_n237), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT4), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n314), .A2(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n310), .B1(new_n313), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n306), .A2(KEYINPUT4), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n305), .B(new_n315), .C1(new_n214), .C2(new_n215), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n321), .A2(new_n322), .B1(new_n311), .B2(new_n239), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(new_n280), .A3(new_n308), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n279), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n325), .A2(KEYINPUT86), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n320), .A2(new_n279), .A3(new_n324), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT6), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n325), .A2(KEYINPUT86), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n326), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G226gat), .ZN(new_n333));
  INV_X1    g132(.A(G233gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n337));
  NOR2_X1   g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT23), .ZN(new_n339));
  NAND2_X1  g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(G169gat), .B2(G176gat), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT65), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT65), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n346), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(G183gat), .A2(G190gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT24), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G183gat), .ZN(new_n351));
  INV_X1    g150(.A(G190gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n345), .A2(new_n347), .A3(new_n350), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n343), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT67), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(new_n351), .A3(new_n352), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT66), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n350), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT66), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n360), .A2(new_n362), .A3(new_n344), .A4(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n339), .A2(KEYINPUT25), .A3(new_n342), .A4(new_n340), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n355), .A2(new_n356), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n348), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT68), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT68), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n372), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n340), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT26), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(new_n338), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n369), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n351), .A2(KEYINPUT27), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT27), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G183gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n381), .A3(new_n352), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT28), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT27), .B(G183gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n385), .A2(KEYINPUT28), .A3(new_n352), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n378), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n337), .B1(new_n368), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n378), .A2(new_n387), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT25), .B1(new_n343), .B2(new_n354), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n363), .B(new_n361), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n349), .A2(new_n351), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n359), .A2(new_n358), .B1(new_n393), .B2(G190gat), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n366), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n390), .B(KEYINPUT78), .C1(new_n391), .C2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n336), .B1(new_n389), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n335), .A2(KEYINPUT29), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n390), .A2(KEYINPUT69), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT69), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n378), .A2(new_n387), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n355), .A2(new_n356), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n365), .A2(new_n367), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n399), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n242), .A2(new_n247), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n397), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n389), .A2(new_n396), .A3(new_n398), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n403), .A2(new_n406), .A3(new_n335), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT37), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n411), .A2(new_n412), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n408), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT78), .B1(new_n406), .B2(new_n390), .ZN(new_n419));
  INV_X1    g218(.A(new_n396), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n335), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n378), .A2(new_n387), .A3(new_n401), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n401), .B1(new_n378), .B2(new_n387), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n406), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n398), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(new_n409), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n418), .A2(new_n426), .A3(KEYINPUT37), .ZN(new_n427));
  XOR2_X1   g226(.A(G8gat), .B(G36gat), .Z(new_n428));
  XNOR2_X1  g227(.A(G64gat), .B(G92gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n430), .B(KEYINPUT79), .Z(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(KEYINPUT38), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n427), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n325), .A2(KEYINPUT6), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n409), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n421), .A2(new_n408), .A3(new_n425), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(new_n430), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n332), .A2(new_n433), .A3(new_n434), .A4(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n430), .B1(new_n414), .B2(new_n415), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n439), .B1(new_n415), .B2(new_n414), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n440), .A2(KEYINPUT38), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n414), .A2(KEYINPUT80), .A3(KEYINPUT30), .A4(new_n430), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT30), .A4(new_n430), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT80), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT30), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n437), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n323), .A2(new_n308), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT39), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT39), .B1(new_n307), .B2(new_n309), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n454), .B(new_n279), .C1(new_n452), .C2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT40), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n325), .B(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n451), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n460), .A2(KEYINPUT87), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(KEYINPUT87), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n275), .B(new_n442), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT73), .B(G71gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(G99gat), .ZN(new_n465));
  XOR2_X1   g264(.A(G15gat), .B(G43gat), .Z(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n424), .A2(new_n305), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n403), .A2(new_n303), .A3(new_n406), .ZN(new_n469));
  NAND2_X1  g268(.A1(G227gat), .A2(G233gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT64), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT33), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(KEYINPUT32), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n472), .B(KEYINPUT32), .C1(new_n473), .C2(new_n467), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n468), .A2(new_n469), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n480), .B1(new_n481), .B2(new_n471), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n471), .B1(new_n468), .B2(new_n469), .ZN(new_n483));
  NAND2_X1  g282(.A1(KEYINPUT74), .A2(KEYINPUT34), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n478), .A2(KEYINPUT75), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT36), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n478), .A2(new_n486), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n476), .A2(new_n477), .A3(new_n482), .A4(new_n485), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n487), .B(new_n488), .C1(new_n491), .C2(KEYINPUT75), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n489), .A2(new_n490), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT36), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n254), .A2(new_n270), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n262), .B1(new_n269), .B2(new_n203), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n272), .B1(new_n496), .B2(G22gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n258), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n273), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n434), .B1(new_n329), .B2(new_n325), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n447), .A2(new_n501), .A3(new_n450), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n492), .A2(new_n494), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n499), .A2(new_n273), .A3(new_n490), .A4(new_n489), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT35), .B1(new_n504), .B2(new_n502), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT89), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(KEYINPUT89), .B(KEYINPUT35), .C1(new_n504), .C2(new_n502), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n459), .A2(new_n330), .B1(KEYINPUT6), .B2(new_n325), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT88), .B1(new_n510), .B2(new_n451), .ZN(new_n511));
  INV_X1    g310(.A(new_n451), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n332), .A2(new_n434), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT88), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n487), .B1(new_n491), .B2(KEYINPUT75), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n511), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n463), .A2(new_n503), .B1(new_n509), .B2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT91), .ZN(new_n521));
  XOR2_X1   g320(.A(G113gat), .B(G141gat), .Z(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G169gat), .B(G197gat), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n523), .B(new_n524), .Z(new_n525));
  INV_X1    g324(.A(KEYINPUT12), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT92), .ZN(new_n528));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT16), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(G1gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n531), .B1(G1gat), .B2(new_n529), .ZN(new_n532));
  INV_X1    g331(.A(G8gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(G36gat), .ZN(new_n535));
  AND2_X1   g334(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n536));
  NOR2_X1   g335(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(G29gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n541), .A2(KEYINPUT15), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(KEYINPUT15), .ZN(new_n543));
  XNOR2_X1  g342(.A(G43gat), .B(G50gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n543), .A2(new_n544), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(KEYINPUT17), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n549), .B1(new_n545), .B2(new_n546), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n528), .B(new_n534), .C1(new_n548), .C2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n534), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n545), .A2(new_n546), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n549), .ZN(new_n554));
  INV_X1    g353(.A(new_n550), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n552), .A2(new_n547), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT92), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n551), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT18), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n559), .A2(KEYINPUT93), .A3(new_n560), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n559), .A2(KEYINPUT18), .A3(new_n560), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n553), .A2(new_n534), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n557), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n560), .B(KEYINPUT13), .Z(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n527), .B1(new_n565), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT95), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n561), .A2(new_n562), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT18), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n574), .A2(KEYINPUT94), .A3(new_n575), .A4(new_n564), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n527), .A2(new_n570), .A3(new_n566), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT94), .B1(new_n563), .B2(new_n564), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n573), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT94), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n582), .A2(KEYINPUT95), .A3(new_n576), .A4(new_n577), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n572), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n519), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G127gat), .B(G155gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G57gat), .B(G64gat), .Z(new_n589));
  XOR2_X1   g388(.A(G71gat), .B(G78gat), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT9), .ZN(new_n592));
  INV_X1    g391(.A(G71gat), .ZN(new_n593));
  INV_X1    g392(.A(G78gat), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n589), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n589), .A2(new_n595), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n590), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n598), .A3(KEYINPUT96), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT96), .B1(new_n596), .B2(new_n598), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT21), .ZN(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n604), .B1(new_n602), .B2(new_n603), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n588), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n606), .A2(new_n607), .A3(new_n588), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n586), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  INV_X1    g411(.A(new_n586), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(new_n613), .A3(new_n608), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G183gat), .B(G211gat), .Z(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n611), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n534), .B1(new_n602), .B2(new_n603), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT97), .B(KEYINPUT98), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n617), .A2(new_n623), .A3(new_n619), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT99), .B(G85gat), .ZN(new_n629));
  INV_X1    g428(.A(G92gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G85gat), .A2(G92gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT7), .ZN(new_n633));
  INV_X1    g432(.A(G99gat), .ZN(new_n634));
  INV_X1    g433(.A(G106gat), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT8), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n631), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G99gat), .B(G106gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(new_n548), .B2(new_n550), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n642));
  AND2_X1   g441(.A1(G232gat), .A2(G233gat), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n547), .A2(new_n639), .B1(KEYINPUT41), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n642), .B1(new_n641), .B2(new_n644), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G134gat), .B(G162gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n645), .B2(new_n646), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n643), .A2(KEYINPUT41), .ZN(new_n653));
  XNOR2_X1  g452(.A(G190gat), .B(G218gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n650), .A2(new_n655), .A3(new_n651), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT10), .ZN(new_n661));
  INV_X1    g460(.A(new_n601), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n639), .B1(new_n599), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n596), .A2(new_n598), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n639), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n661), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(new_n599), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n667), .A2(KEYINPUT101), .A3(KEYINPUT10), .A4(new_n639), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT10), .B1(new_n600), .B2(new_n601), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n669), .B1(new_n670), .B2(new_n640), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n666), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(G230gat), .A2(G233gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OR3_X1    g473(.A1(new_n663), .A2(new_n665), .A3(new_n673), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(G120gat), .B(G148gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT102), .ZN(new_n678));
  XOR2_X1   g477(.A(G176gat), .B(G204gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n680), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n628), .A2(new_n660), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n585), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n501), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g490(.A1(new_n687), .A2(new_n512), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT16), .B(G8gat), .Z(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n533), .B2(new_n692), .ZN(new_n695));
  MUX2_X1   g494(.A(new_n694), .B(new_n695), .S(KEYINPUT42), .Z(G1325gat));
  AOI21_X1  g495(.A(G15gat), .B1(new_n688), .B2(new_n516), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n492), .A2(new_n494), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G15gat), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT103), .Z(new_n701));
  AOI21_X1  g500(.A(new_n697), .B1(new_n688), .B2(new_n701), .ZN(G1326gat));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n275), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT43), .B(G22gat), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  NOR2_X1   g504(.A1(new_n628), .A2(new_n683), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n585), .A2(new_n659), .A3(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n707), .A2(G29gat), .A3(new_n501), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT45), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT44), .B1(new_n519), .B2(new_n660), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n447), .A2(new_n501), .A3(new_n450), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(new_n275), .A3(new_n493), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT89), .B1(new_n712), .B2(KEYINPUT35), .ZN(new_n713));
  INV_X1    g512(.A(new_n508), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n518), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n509), .A2(KEYINPUT104), .A3(new_n518), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n717), .A2(new_n718), .B1(new_n463), .B2(new_n503), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n720));
  NOR2_X1   g519(.A1(new_n660), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n710), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n580), .A2(new_n583), .ZN(new_n724));
  INV_X1    g523(.A(new_n572), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n723), .A2(new_n726), .A3(new_n706), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n539), .B1(new_n727), .B2(new_n689), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n709), .A2(new_n728), .ZN(G1328gat));
  AND2_X1   g528(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n707), .A2(G36gat), .A3(new_n512), .ZN(new_n733));
  MUX2_X1   g532(.A(new_n732), .B(new_n730), .S(new_n733), .Z(new_n734));
  AND2_X1   g533(.A1(new_n727), .A2(new_n451), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n535), .B2(new_n735), .ZN(G1329gat));
  INV_X1    g535(.A(new_n516), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n707), .A2(G43gat), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n727), .A2(new_n699), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(G43gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g540(.A1(new_n707), .A2(G50gat), .A3(new_n275), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n500), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(G50gat), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g544(.A1(new_n717), .A2(new_n718), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n463), .A2(new_n503), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR4_X1   g547(.A1(new_n726), .A2(new_n627), .A3(new_n659), .A4(new_n684), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n501), .B(KEYINPUT107), .Z(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G57gat), .ZN(G1332gat));
  INV_X1    g552(.A(new_n750), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n512), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  AND2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n755), .B2(new_n756), .ZN(G1333gat));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n754), .B2(new_n737), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n750), .A2(KEYINPUT108), .A3(new_n516), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(new_n593), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n750), .A2(G71gat), .A3(new_n699), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n500), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g567(.A1(new_n584), .A2(new_n627), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(KEYINPUT109), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(KEYINPUT109), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n684), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n723), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n774), .A2(new_n689), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n775), .A2(KEYINPUT110), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(KEYINPUT110), .ZN(new_n777));
  OR3_X1    g576(.A1(new_n776), .A2(new_n777), .A3(new_n629), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  INV_X1    g578(.A(new_n772), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n659), .B1(new_n780), .B2(new_n770), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n781), .B2(new_n719), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n660), .B1(new_n771), .B2(new_n772), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n783), .A2(KEYINPUT51), .A3(new_n748), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n683), .A2(new_n689), .A3(new_n629), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT111), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n778), .B1(new_n785), .B2(new_n787), .ZN(G1336gat));
  AOI21_X1  g587(.A(new_n630), .B1(new_n774), .B2(new_n451), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n782), .A2(new_n784), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n684), .A2(new_n512), .A3(G92gat), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  XOR2_X1   g591(.A(new_n792), .B(KEYINPUT52), .Z(G1337gat));
  AND2_X1   g592(.A1(new_n774), .A2(new_n699), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n516), .A2(new_n634), .A3(new_n683), .ZN(new_n795));
  XOR2_X1   g594(.A(new_n795), .B(KEYINPUT112), .Z(new_n796));
  OAI22_X1  g595(.A1(new_n794), .A2(new_n634), .B1(new_n785), .B2(new_n796), .ZN(G1338gat));
  NOR3_X1   g596(.A1(new_n684), .A2(new_n275), .A3(G106gat), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n790), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n722), .B1(new_n746), .B2(new_n747), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n747), .A2(new_n715), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(new_n659), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n500), .B(new_n773), .C1(new_n800), .C2(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n804), .A2(G106gat), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT53), .B1(new_n799), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n723), .A2(KEYINPUT113), .A3(new_n500), .A4(new_n773), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(G106gat), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT53), .B1(new_n790), .B2(new_n798), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n810), .A2(KEYINPUT114), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT114), .B1(new_n810), .B2(new_n811), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n806), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g615(.A(KEYINPUT115), .B(new_n806), .C1(new_n812), .C2(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1339gat));
  INV_X1    g617(.A(new_n673), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n666), .A2(new_n671), .A3(new_n819), .A4(new_n668), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n674), .A2(KEYINPUT54), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n672), .A2(new_n822), .A3(new_n673), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n821), .A2(KEYINPUT55), .A3(new_n680), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n681), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n823), .A2(new_n680), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT55), .B1(new_n826), .B2(new_n821), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT116), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n821), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n831), .A2(new_n832), .A3(new_n681), .A4(new_n824), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n828), .A2(new_n833), .A3(new_n659), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n568), .A2(new_n569), .ZN(new_n835));
  INV_X1    g634(.A(new_n559), .ZN(new_n836));
  INV_X1    g635(.A(new_n560), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n525), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n580), .B2(new_n583), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n834), .A2(new_n840), .A3(KEYINPUT117), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT117), .B1(new_n834), .B2(new_n840), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n833), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n726), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n840), .A2(new_n683), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n659), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n627), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n685), .A2(new_n726), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n500), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n451), .A2(new_n501), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n516), .A3(new_n853), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(new_n289), .A3(new_n584), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n849), .A2(new_n851), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n856), .A2(new_n751), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n504), .A2(new_n451), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n726), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n855), .B1(new_n861), .B2(new_n289), .ZN(G1340gat));
  OAI21_X1  g661(.A(G120gat), .B1(new_n854), .B2(new_n684), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n683), .A2(new_n291), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT118), .Z(G1341gat));
  NOR3_X1   g665(.A1(new_n854), .A2(new_n281), .A3(new_n627), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n859), .A2(KEYINPUT119), .A3(new_n627), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(G127gat), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT119), .B1(new_n859), .B2(new_n627), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(G1342gat));
  OR3_X1    g670(.A1(new_n859), .A2(new_n286), .A3(new_n660), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n873));
  OAI21_X1  g672(.A(G134gat), .B1(new_n854), .B2(new_n660), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(G1343gat));
  AND2_X1   g675(.A1(new_n698), .A2(new_n853), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n275), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n834), .A2(new_n840), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n834), .A2(new_n840), .A3(KEYINPUT117), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n825), .B1(new_n829), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n584), .A2(new_n888), .ZN(new_n889));
  AOI211_X1 g688(.A(new_n684), .B(new_n839), .C1(new_n580), .C2(new_n583), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n660), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n628), .B1(new_n885), .B2(new_n891), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n878), .B(new_n880), .C1(new_n892), .C2(new_n850), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n275), .B1(new_n849), .B2(new_n851), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(KEYINPUT57), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n726), .A2(new_n887), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n659), .B1(new_n896), .B2(new_n847), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n627), .B1(new_n843), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n851), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n878), .B1(new_n899), .B2(new_n880), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n877), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G141gat), .B1(new_n901), .B2(new_n584), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n698), .A2(new_n500), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(new_n451), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n857), .A2(new_n904), .ZN(new_n905));
  OR3_X1    g704(.A1(new_n905), .A2(G141gat), .A3(new_n584), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT58), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n902), .A2(new_n909), .A3(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1344gat));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n584), .A2(new_n844), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n660), .B1(new_n913), .B2(new_n890), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n628), .B1(new_n885), .B2(new_n914), .ZN(new_n915));
  OAI211_X1 g714(.A(KEYINPUT57), .B(new_n500), .C1(new_n915), .C2(new_n850), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n825), .A2(new_n827), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n840), .A2(new_n659), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n847), .B1(new_n584), .B2(new_n888), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n920), .B2(new_n660), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n851), .B1(new_n921), .B2(new_n628), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT57), .B1(new_n922), .B2(new_n500), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n683), .B(new_n877), .C1(new_n917), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G148gat), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n683), .B(new_n877), .C1(new_n895), .C2(new_n900), .ZN(new_n926));
  INV_X1    g725(.A(G148gat), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(KEYINPUT59), .ZN(new_n928));
  AOI22_X1  g727(.A1(new_n925), .A2(KEYINPUT59), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n905), .A2(G148gat), .A3(new_n684), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n912), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n930), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n926), .A2(new_n928), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n934), .B1(new_n924), .B2(G148gat), .ZN(new_n935));
  OAI211_X1 g734(.A(KEYINPUT122), .B(new_n932), .C1(new_n933), .C2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n931), .A2(new_n936), .ZN(G1345gat));
  OAI21_X1  g736(.A(G155gat), .B1(new_n901), .B2(new_n627), .ZN(new_n938));
  INV_X1    g737(.A(new_n905), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n205), .A3(new_n628), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1346gat));
  OAI21_X1  g740(.A(G162gat), .B1(new_n901), .B2(new_n660), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n939), .A2(new_n206), .A3(new_n659), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1347gat));
  AOI21_X1  g743(.A(new_n689), .B1(new_n849), .B2(new_n851), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n504), .A2(new_n512), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n947), .A2(G169gat), .A3(new_n584), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT123), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n751), .A2(new_n512), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n516), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT124), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n852), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(G169gat), .B1(new_n953), .B2(new_n584), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n949), .A2(new_n954), .ZN(G1348gat));
  OAI21_X1  g754(.A(G176gat), .B1(new_n953), .B2(new_n684), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n684), .A2(G176gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n947), .B2(new_n957), .ZN(G1349gat));
  OAI21_X1  g757(.A(G183gat), .B1(new_n953), .B2(new_n627), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n628), .A2(new_n385), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n947), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g761(.A(G190gat), .B1(new_n953), .B2(new_n660), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT125), .ZN(new_n964));
  XOR2_X1   g763(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n945), .A2(new_n352), .A3(new_n659), .A4(new_n946), .ZN(new_n967));
  OR2_X1    g766(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n966), .B(new_n967), .C1(new_n964), .C2(new_n968), .ZN(G1351gat));
  NOR2_X1   g768(.A1(new_n903), .A2(new_n512), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n945), .A2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g771(.A(G197gat), .B1(new_n972), .B2(new_n726), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n917), .A2(new_n923), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n950), .A2(new_n698), .ZN(new_n975));
  XOR2_X1   g774(.A(new_n975), .B(KEYINPUT127), .Z(new_n976));
  INV_X1    g775(.A(G197gat), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n976), .A2(new_n977), .A3(new_n584), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n973), .B1(new_n974), .B2(new_n978), .ZN(G1352gat));
  NAND2_X1  g778(.A1(new_n974), .A2(new_n683), .ZN(new_n980));
  OAI21_X1  g779(.A(G204gat), .B1(new_n980), .B2(new_n976), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n971), .A2(G204gat), .A3(new_n684), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT62), .ZN(new_n983));
  OR2_X1    g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(G1353gat));
  NOR2_X1   g785(.A1(new_n975), .A2(new_n627), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n229), .B1(new_n974), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT63), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n229), .A3(new_n628), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1354gat));
  AOI21_X1  g790(.A(G218gat), .B1(new_n972), .B2(new_n659), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n976), .A2(new_n244), .A3(new_n660), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n992), .B1(new_n974), .B2(new_n993), .ZN(G1355gat));
endmodule


