

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U321 ( .A(n446), .B(n445), .ZN(n450) );
  NOR2_X1 U322 ( .A1(n474), .A2(n473), .ZN(n560) );
  XOR2_X1 U323 ( .A(n377), .B(n306), .Z(n524) );
  AND2_X1 U324 ( .A1(G230GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U325 ( .A(n435), .B(n289), .ZN(n437) );
  XOR2_X1 U326 ( .A(G120GAT), .B(G71GAT), .Z(n435) );
  XNOR2_X1 U327 ( .A(n437), .B(n436), .ZN(n439) );
  INV_X1 U328 ( .A(n326), .ZN(n300) );
  XNOR2_X1 U329 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U330 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U331 ( .A(KEYINPUT99), .B(KEYINPUT26), .ZN(n404) );
  XNOR2_X1 U332 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n466) );
  XNOR2_X1 U333 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U334 ( .A(n405), .B(n404), .ZN(n568) );
  XNOR2_X1 U335 ( .A(n467), .B(n466), .ZN(n538) );
  OR2_X1 U336 ( .A1(n513), .A2(n483), .ZN(n452) );
  XNOR2_X1 U337 ( .A(n575), .B(KEYINPUT41), .ZN(n546) );
  INV_X1 U338 ( .A(G43GAT), .ZN(n453) );
  XNOR2_X1 U339 ( .A(n452), .B(KEYINPUT38), .ZN(n499) );
  XNOR2_X1 U340 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U341 ( .A(n453), .B(KEYINPUT40), .ZN(n454) );
  XNOR2_X1 U342 ( .A(n478), .B(n477), .ZN(G1349GAT) );
  XNOR2_X1 U343 ( .A(n455), .B(n454), .ZN(G1330GAT) );
  XOR2_X1 U344 ( .A(KEYINPUT83), .B(KEYINPUT17), .Z(n291) );
  XNOR2_X1 U345 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n290) );
  XNOR2_X1 U346 ( .A(n291), .B(n290), .ZN(n292) );
  XNOR2_X1 U347 ( .A(KEYINPUT19), .B(n292), .ZN(n377) );
  XOR2_X1 U348 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n294) );
  XNOR2_X1 U349 ( .A(G169GAT), .B(G113GAT), .ZN(n293) );
  XNOR2_X1 U350 ( .A(n294), .B(n293), .ZN(n305) );
  XOR2_X1 U351 ( .A(KEYINPUT0), .B(KEYINPUT81), .Z(n362) );
  XOR2_X1 U352 ( .A(G99GAT), .B(n362), .Z(n296) );
  XNOR2_X1 U353 ( .A(G43GAT), .B(n435), .ZN(n295) );
  XNOR2_X1 U354 ( .A(n296), .B(n295), .ZN(n303) );
  XOR2_X1 U355 ( .A(G190GAT), .B(G134GAT), .Z(n309) );
  XOR2_X1 U356 ( .A(KEYINPUT82), .B(G176GAT), .Z(n298) );
  NAND2_X1 U357 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U358 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U359 ( .A(n309), .B(n299), .ZN(n301) );
  XOR2_X1 U360 ( .A(G15GAT), .B(G127GAT), .Z(n326) );
  XOR2_X1 U361 ( .A(n305), .B(n304), .Z(n306) );
  INV_X1 U362 ( .A(n524), .ZN(n474) );
  XOR2_X1 U363 ( .A(KEYINPUT73), .B(G92GAT), .Z(n308) );
  XNOR2_X1 U364 ( .A(G99GAT), .B(G85GAT), .ZN(n307) );
  XNOR2_X1 U365 ( .A(n308), .B(n307), .ZN(n440) );
  XOR2_X1 U366 ( .A(n440), .B(n309), .Z(n311) );
  NAND2_X1 U367 ( .A1(G232GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U369 ( .A(KEYINPUT11), .B(KEYINPUT76), .Z(n313) );
  XNOR2_X1 U370 ( .A(G162GAT), .B(G106GAT), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U372 ( .A(n315), .B(n314), .Z(n325) );
  XOR2_X1 U373 ( .A(G43GAT), .B(G29GAT), .Z(n317) );
  XNOR2_X1 U374 ( .A(KEYINPUT8), .B(G50GAT), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U376 ( .A(n318), .B(KEYINPUT69), .Z(n320) );
  XNOR2_X1 U377 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n434) );
  XOR2_X1 U379 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n322) );
  XNOR2_X1 U380 ( .A(G218GAT), .B(KEYINPUT64), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n434), .B(n323), .ZN(n324) );
  XNOR2_X1 U383 ( .A(n325), .B(n324), .ZN(n559) );
  XOR2_X1 U384 ( .A(KEYINPUT36), .B(n559), .Z(n582) );
  XOR2_X1 U385 ( .A(G57GAT), .B(KEYINPUT13), .Z(n447) );
  XOR2_X1 U386 ( .A(n447), .B(G78GAT), .Z(n328) );
  XNOR2_X1 U387 ( .A(n326), .B(G211GAT), .ZN(n327) );
  XNOR2_X1 U388 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U389 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n330) );
  XNOR2_X1 U390 ( .A(G8GAT), .B(KEYINPUT14), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U392 ( .A(n332), .B(n331), .Z(n334) );
  XNOR2_X1 U393 ( .A(G22GAT), .B(G155GAT), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U395 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n336) );
  NAND2_X1 U396 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U397 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U398 ( .A(n338), .B(n337), .Z(n343) );
  XOR2_X1 U399 ( .A(G64GAT), .B(G71GAT), .Z(n340) );
  XNOR2_X1 U400 ( .A(G1GAT), .B(G183GAT), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n341), .B(KEYINPUT77), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n579) );
  XOR2_X1 U404 ( .A(KEYINPUT88), .B(G162GAT), .Z(n345) );
  XNOR2_X1 U405 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U407 ( .A(KEYINPUT3), .B(n346), .Z(n398) );
  XOR2_X1 U408 ( .A(G148GAT), .B(G127GAT), .Z(n348) );
  XNOR2_X1 U409 ( .A(G141GAT), .B(G134GAT), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U411 ( .A(n349), .B(G85GAT), .Z(n351) );
  XOR2_X1 U412 ( .A(G113GAT), .B(G1GAT), .Z(n417) );
  XNOR2_X1 U413 ( .A(G29GAT), .B(n417), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n398), .B(n352), .ZN(n366) );
  XOR2_X1 U416 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n354) );
  XNOR2_X1 U417 ( .A(G120GAT), .B(KEYINPUT93), .ZN(n353) );
  XNOR2_X1 U418 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U419 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n356) );
  XNOR2_X1 U420 ( .A(KEYINPUT90), .B(G57GAT), .ZN(n355) );
  XNOR2_X1 U421 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U422 ( .A(n358), .B(n357), .Z(n364) );
  XOR2_X1 U423 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n360) );
  NAND2_X1 U424 ( .A1(G225GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U425 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n366), .B(n365), .ZN(n493) );
  XOR2_X1 U429 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n368) );
  XNOR2_X1 U430 ( .A(G190GAT), .B(KEYINPUT96), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U432 ( .A(n369), .B(G92GAT), .Z(n371) );
  XOR2_X1 U433 ( .A(G176GAT), .B(G64GAT), .Z(n448) );
  XNOR2_X1 U434 ( .A(G36GAT), .B(n448), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n376) );
  XNOR2_X1 U436 ( .A(G169GAT), .B(G197GAT), .ZN(n372) );
  XNOR2_X1 U437 ( .A(n372), .B(G8GAT), .ZN(n430) );
  XOR2_X1 U438 ( .A(n430), .B(KEYINPUT97), .Z(n374) );
  NAND2_X1 U439 ( .A1(G226GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U440 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U441 ( .A(n376), .B(n375), .Z(n383) );
  INV_X1 U442 ( .A(n377), .ZN(n381) );
  XOR2_X1 U443 ( .A(KEYINPUT87), .B(G218GAT), .Z(n379) );
  XNOR2_X1 U444 ( .A(G211GAT), .B(G204GAT), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U446 ( .A(KEYINPUT21), .B(n380), .Z(n394) );
  XNOR2_X1 U447 ( .A(n381), .B(n394), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n496) );
  XOR2_X1 U449 ( .A(n496), .B(KEYINPUT27), .Z(n406) );
  XOR2_X1 U450 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n385) );
  XNOR2_X1 U451 ( .A(G50GAT), .B(KEYINPUT85), .ZN(n384) );
  XNOR2_X1 U452 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U453 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n387) );
  XNOR2_X1 U454 ( .A(G197GAT), .B(KEYINPUT86), .ZN(n386) );
  XNOR2_X1 U455 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U456 ( .A(n389), .B(n388), .Z(n396) );
  XOR2_X1 U457 ( .A(G141GAT), .B(G22GAT), .Z(n418) );
  XNOR2_X1 U458 ( .A(G106GAT), .B(G78GAT), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n390), .B(G148GAT), .ZN(n436) );
  XOR2_X1 U460 ( .A(n418), .B(n436), .Z(n392) );
  NAND2_X1 U461 ( .A1(G228GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U462 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U463 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U464 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U465 ( .A(n398), .B(n397), .ZN(n471) );
  XOR2_X1 U466 ( .A(KEYINPUT28), .B(n471), .Z(n498) );
  NAND2_X1 U467 ( .A1(n406), .A2(n498), .ZN(n399) );
  NOR2_X1 U468 ( .A1(n493), .A2(n399), .ZN(n525) );
  XNOR2_X1 U469 ( .A(n525), .B(KEYINPUT98), .ZN(n400) );
  NAND2_X1 U470 ( .A1(n400), .A2(n474), .ZN(n411) );
  NOR2_X1 U471 ( .A1(n474), .A2(n496), .ZN(n401) );
  XNOR2_X1 U472 ( .A(n401), .B(KEYINPUT100), .ZN(n402) );
  NOR2_X1 U473 ( .A1(n471), .A2(n402), .ZN(n403) );
  XNOR2_X1 U474 ( .A(KEYINPUT25), .B(n403), .ZN(n407) );
  NAND2_X1 U475 ( .A1(n471), .A2(n474), .ZN(n405) );
  NAND2_X1 U476 ( .A1(n406), .A2(n568), .ZN(n537) );
  NAND2_X1 U477 ( .A1(n407), .A2(n537), .ZN(n408) );
  NAND2_X1 U478 ( .A1(n408), .A2(n493), .ZN(n409) );
  XOR2_X1 U479 ( .A(KEYINPUT101), .B(n409), .Z(n410) );
  NAND2_X1 U480 ( .A1(n411), .A2(n410), .ZN(n481) );
  NAND2_X1 U481 ( .A1(n579), .A2(n481), .ZN(n412) );
  NOR2_X1 U482 ( .A1(n582), .A2(n412), .ZN(n414) );
  XNOR2_X1 U483 ( .A(KEYINPUT37), .B(KEYINPUT104), .ZN(n413) );
  XNOR2_X1 U484 ( .A(n414), .B(n413), .ZN(n513) );
  XOR2_X1 U485 ( .A(KEYINPUT70), .B(KEYINPUT68), .Z(n416) );
  XNOR2_X1 U486 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n415) );
  XNOR2_X1 U487 ( .A(n416), .B(n415), .ZN(n422) );
  XNOR2_X1 U488 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U489 ( .A(KEYINPUT66), .B(G15GAT), .Z(n419) );
  XNOR2_X1 U490 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U491 ( .A(n422), .B(n421), .ZN(n423) );
  AND2_X1 U492 ( .A1(G229GAT), .A2(G233GAT), .ZN(n424) );
  NAND2_X1 U493 ( .A1(n423), .A2(n424), .ZN(n428) );
  INV_X1 U494 ( .A(n423), .ZN(n426) );
  INV_X1 U495 ( .A(n424), .ZN(n425) );
  NAND2_X1 U496 ( .A1(n426), .A2(n425), .ZN(n427) );
  NAND2_X1 U497 ( .A1(n428), .A2(n427), .ZN(n429) );
  XOR2_X1 U498 ( .A(n429), .B(KEYINPUT30), .Z(n432) );
  XNOR2_X1 U499 ( .A(n430), .B(KEYINPUT65), .ZN(n431) );
  XNOR2_X1 U500 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U501 ( .A(n434), .B(n433), .Z(n570) );
  XNOR2_X1 U502 ( .A(KEYINPUT71), .B(n570), .ZN(n554) );
  INV_X1 U503 ( .A(KEYINPUT32), .ZN(n438) );
  XNOR2_X1 U504 ( .A(n439), .B(n438), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n440), .B(KEYINPUT31), .ZN(n444) );
  XOR2_X1 U506 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n442) );
  XNOR2_X1 U507 ( .A(G204GAT), .B(KEYINPUT74), .ZN(n441) );
  XOR2_X1 U508 ( .A(n442), .B(n441), .Z(n443) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U510 ( .A(n450), .B(n449), .ZN(n575) );
  NAND2_X1 U511 ( .A1(n554), .A2(n575), .ZN(n451) );
  XOR2_X1 U512 ( .A(KEYINPUT75), .B(n451), .Z(n483) );
  NOR2_X1 U513 ( .A1(n474), .A2(n499), .ZN(n455) );
  NOR2_X1 U514 ( .A1(n582), .A2(n579), .ZN(n456) );
  XOR2_X1 U515 ( .A(KEYINPUT45), .B(n456), .Z(n457) );
  NOR2_X1 U516 ( .A1(n554), .A2(n457), .ZN(n458) );
  NAND2_X1 U517 ( .A1(n458), .A2(n575), .ZN(n465) );
  INV_X1 U518 ( .A(n570), .ZN(n542) );
  NAND2_X1 U519 ( .A1(n542), .A2(n546), .ZN(n459) );
  XNOR2_X1 U520 ( .A(KEYINPUT46), .B(n459), .ZN(n460) );
  NAND2_X1 U521 ( .A1(n460), .A2(n579), .ZN(n461) );
  NOR2_X1 U522 ( .A1(n559), .A2(n461), .ZN(n463) );
  XNOR2_X1 U523 ( .A(KEYINPUT110), .B(KEYINPUT47), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n463), .B(n462), .ZN(n464) );
  NAND2_X1 U525 ( .A1(n465), .A2(n464), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n496), .A2(n538), .ZN(n469) );
  XNOR2_X1 U527 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U529 ( .A1(n470), .A2(n493), .ZN(n567) );
  NOR2_X1 U530 ( .A1(n471), .A2(n567), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n472), .B(KEYINPUT55), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n560), .A2(n546), .ZN(n478) );
  XOR2_X1 U533 ( .A(KEYINPUT57), .B(KEYINPUT119), .Z(n476) );
  XOR2_X1 U534 ( .A(G176GAT), .B(KEYINPUT56), .Z(n475) );
  INV_X1 U535 ( .A(n493), .ZN(n540) );
  XNOR2_X1 U536 ( .A(KEYINPUT80), .B(KEYINPUT16), .ZN(n480) );
  NOR2_X1 U537 ( .A1(n559), .A2(n579), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(n482) );
  NAND2_X1 U539 ( .A1(n482), .A2(n481), .ZN(n502) );
  NOR2_X1 U540 ( .A1(n483), .A2(n502), .ZN(n491) );
  NAND2_X1 U541 ( .A1(n540), .A2(n491), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n484), .B(KEYINPUT34), .ZN(n485) );
  XOR2_X1 U543 ( .A(n485), .B(KEYINPUT103), .Z(n487) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(KEYINPUT102), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(G1324GAT) );
  INV_X1 U546 ( .A(n496), .ZN(n515) );
  NAND2_X1 U547 ( .A1(n515), .A2(n491), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U550 ( .A1(n491), .A2(n524), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  INV_X1 U552 ( .A(n498), .ZN(n520) );
  NAND2_X1 U553 ( .A1(n491), .A2(n520), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n495) );
  NOR2_X1 U556 ( .A1(n493), .A2(n499), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U558 ( .A1(n496), .A2(n499), .ZN(n497) );
  XOR2_X1 U559 ( .A(G36GAT), .B(n497), .Z(G1329GAT) );
  NOR2_X1 U560 ( .A1(n499), .A2(n498), .ZN(n500) );
  XOR2_X1 U561 ( .A(G50GAT), .B(n500), .Z(G1331GAT) );
  XNOR2_X1 U562 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  NAND2_X1 U563 ( .A1(n546), .A2(n570), .ZN(n501) );
  XOR2_X1 U564 ( .A(KEYINPUT105), .B(n501), .Z(n512) );
  NOR2_X1 U565 ( .A1(n512), .A2(n502), .ZN(n508) );
  NAND2_X1 U566 ( .A1(n508), .A2(n540), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U568 ( .A1(n515), .A2(n508), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(KEYINPUT106), .ZN(n506) );
  XNOR2_X1 U570 ( .A(G64GAT), .B(n506), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n524), .A2(n508), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U574 ( .A1(n508), .A2(n520), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U576 ( .A(G78GAT), .B(n511), .Z(G1335GAT) );
  NOR2_X1 U577 ( .A1(n513), .A2(n512), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n540), .A2(n521), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(G85GAT), .ZN(G1336GAT) );
  XNOR2_X1 U580 ( .A(G92GAT), .B(KEYINPUT108), .ZN(n517) );
  NAND2_X1 U581 ( .A1(n521), .A2(n515), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1337GAT) );
  XOR2_X1 U583 ( .A(G99GAT), .B(KEYINPUT109), .Z(n519) );
  NAND2_X1 U584 ( .A1(n521), .A2(n524), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1338GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(KEYINPUT44), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U590 ( .A1(n538), .A2(n526), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n554), .A2(n534), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n529) );
  NAND2_X1 U594 ( .A1(n534), .A2(n546), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(G120GAT), .B(n530), .ZN(G1341GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT113), .B(KEYINPUT50), .Z(n532) );
  INV_X1 U598 ( .A(n579), .ZN(n556) );
  NAND2_X1 U599 ( .A1(n534), .A2(n556), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U603 ( .A1(n534), .A2(n559), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(G1343GAT) );
  NOR2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U607 ( .A(KEYINPUT114), .B(n541), .Z(n552) );
  NAND2_X1 U608 ( .A1(n552), .A2(n542), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT117), .B(KEYINPUT116), .Z(n545) );
  XNOR2_X1 U611 ( .A(KEYINPUT52), .B(KEYINPUT53), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n550) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT115), .ZN(n548) );
  NAND2_X1 U614 ( .A1(n546), .A2(n552), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n552), .A2(n556), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n559), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n560), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n556), .A2(n560), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(KEYINPUT120), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G183GAT), .B(n558), .ZN(G1350GAT) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(KEYINPUT121), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n562) );
  XOR2_X1 U628 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1351GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n566) );
  XNOR2_X1 U632 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n574) );
  INV_X1 U634 ( .A(n567), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n581) );
  NOR2_X1 U636 ( .A1(n570), .A2(n581), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(n574), .B(n573), .Z(G1352GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n581), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n581), .ZN(n580) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

