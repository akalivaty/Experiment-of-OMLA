//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n578, new_n579, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1258, new_n1259, new_n1260;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n461), .A2(G137), .B1(G101), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(G2105), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n470), .B(KEYINPUT66), .ZN(G160));
  NAND2_X1  g046(.A1(new_n461), .A2(G136), .ZN(new_n472));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n472), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  OAI211_X1 g055(.A(G126), .B(G2105), .C1(new_n458), .C2(new_n459), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  INV_X1    g057(.A(G114), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(KEYINPUT67), .A2(G114), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n462), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n481), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n481), .B(KEYINPUT68), .C1(new_n486), .C2(new_n487), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n462), .C1(new_n458), .C2(new_n459), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT3), .B(G2104), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n494), .A2(new_n495), .A3(G138), .A4(new_n462), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n490), .A2(new_n491), .B1(new_n493), .B2(new_n496), .ZN(G164));
  AND2_X1   g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  NOR2_X1   g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  OAI211_X1 g074(.A(G50), .B(G543), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  OAI22_X1  g077(.A1(new_n501), .A2(new_n502), .B1(new_n498), .B2(new_n499), .ZN(new_n503));
  XOR2_X1   g078(.A(KEYINPUT69), .B(G88), .Z(new_n504));
  OAI21_X1  g079(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT70), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT69), .B(G88), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(new_n500), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n502), .A2(new_n501), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n506), .A2(new_n514), .B1(G651), .B2(new_n518), .ZN(G166));
  OAI21_X1  g094(.A(G89), .B1(new_n498), .B2(new_n499), .ZN(new_n520));
  NAND2_X1  g095(.A1(G63), .A2(G651), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n516), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g102(.A(G51), .B(G543), .C1(new_n498), .C2(new_n499), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n522), .A2(new_n529), .ZN(G168));
  NAND3_X1  g105(.A1(new_n509), .A2(new_n510), .A3(G90), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n510), .A2(G52), .A3(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  OAI21_X1  g109(.A(G64), .B1(new_n502), .B2(new_n501), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n533), .A2(new_n537), .ZN(G171));
  AOI22_X1  g113(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n534), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n510), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n541), .A2(new_n542), .B1(new_n503), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  INV_X1    g125(.A(G65), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT71), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G65), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n552), .B(new_n554), .C1(new_n502), .C2(new_n501), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  OAI211_X1 g133(.A(G53), .B(G543), .C1(new_n498), .C2(new_n499), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n510), .A2(new_n561), .A3(G53), .A4(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  OR2_X1    g138(.A1(KEYINPUT6), .A2(G651), .ZN(new_n564));
  NAND2_X1  g139(.A1(KEYINPUT6), .A2(G651), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n507), .A2(new_n508), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G91), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n558), .A2(new_n563), .A3(new_n567), .ZN(G299));
  OAI21_X1  g143(.A(KEYINPUT72), .B1(new_n533), .B2(new_n537), .ZN(new_n569));
  INV_X1    g144(.A(G64), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n507), .B2(new_n508), .ZN(new_n571));
  INV_X1    g146(.A(new_n536), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT72), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n573), .A2(new_n574), .A3(new_n532), .A4(new_n531), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G301));
  INV_X1    g152(.A(new_n522), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n527), .A2(new_n528), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G286));
  NAND2_X1  g155(.A1(new_n518), .A2(G651), .ZN(new_n581));
  INV_X1    g156(.A(new_n514), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n513), .B1(new_n512), .B2(new_n500), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(G303));
  NAND2_X1  g159(.A1(new_n566), .A2(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n586));
  INV_X1    g161(.A(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n564), .B2(new_n565), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G49), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n585), .A2(new_n586), .A3(new_n589), .ZN(G288));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n516), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n566), .A2(G86), .B1(new_n588), .B2(G48), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G305));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n516), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(G651), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n566), .A2(G85), .B1(new_n588), .B2(G47), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n503), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT10), .A4(G92), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(KEYINPUT74), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT74), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G66), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n611), .B(new_n613), .C1(new_n502), .C2(new_n501), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(G54), .B2(new_n588), .ZN(new_n617));
  AND2_X1   g192(.A1(new_n609), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT73), .B1(new_n618), .B2(G868), .ZN(new_n619));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n576), .A2(new_n620), .ZN(new_n621));
  MUX2_X1   g196(.A(new_n619), .B(KEYINPUT73), .S(new_n621), .Z(G321));
  XNOR2_X1  g197(.A(G321), .B(KEYINPUT75), .ZN(G284));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  AND3_X1   g199(.A1(new_n558), .A2(new_n563), .A3(new_n567), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G297));
  XOR2_X1   g201(.A(G297), .B(KEYINPUT76), .Z(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n618), .B1(new_n628), .B2(G860), .ZN(G148));
  OAI21_X1  g204(.A(KEYINPUT78), .B1(new_n545), .B2(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n618), .A2(new_n628), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT77), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  MUX2_X1   g208(.A(KEYINPUT78), .B(new_n630), .S(new_n633), .Z(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n494), .A2(new_n463), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n461), .A2(G135), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT80), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n475), .A2(G123), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n462), .A2(G111), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n643), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n647), .A2(G2096), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n640), .A2(G2100), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(G2096), .ZN(new_n650));
  NAND4_X1  g225(.A1(new_n641), .A2(new_n648), .A3(new_n649), .A4(new_n650), .ZN(G156));
  INV_X1    g226(.A(G14), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT82), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2427), .B(G2430), .Z(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(KEYINPUT14), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2443), .B(G2446), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2451), .B(G2454), .Z(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT83), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT84), .ZN(new_n669));
  AOI211_X1 g244(.A(new_n652), .B(new_n669), .C1(new_n667), .C2(new_n665), .ZN(G401));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT18), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT85), .B(KEYINPUT17), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n671), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n674), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n678), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n672), .B2(new_n673), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n678), .B2(new_n673), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n676), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2096), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n690), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT20), .Z(new_n694));
  AOI211_X1 g269(.A(new_n692), .B(new_n694), .C1(new_n687), .C2(new_n691), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT86), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n698), .A2(new_n699), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n698), .A2(new_n699), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n704), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(G229));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G23), .ZN(new_n710));
  INV_X1    g285(.A(G288), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT33), .B(G1976), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT89), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n712), .B(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(G6), .A2(G16), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G305), .B2(new_n709), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT32), .B(G1981), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT88), .B(G16), .Z(new_n720));
  NOR2_X1   g295(.A1(G166), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G22), .B2(new_n720), .ZN(new_n722));
  INV_X1    g297(.A(G1971), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n715), .B(new_n719), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n723), .B2(new_n722), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT34), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT87), .B(G29), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(G25), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n461), .A2(G131), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n475), .A2(G119), .ZN(new_n732));
  OR2_X1    g307(.A1(G95), .A2(G2105), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n733), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n734));
  AND3_X1   g309(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n730), .B1(new_n735), .B2(new_n729), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT35), .B(G1991), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n720), .ZN(new_n739));
  MUX2_X1   g314(.A(G24), .B(G290), .S(new_n739), .Z(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(G1986), .Z(new_n741));
  NAND3_X1  g316(.A1(new_n727), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n742), .A2(KEYINPUT90), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(KEYINPUT90), .ZN(new_n744));
  OAI22_X1  g319(.A1(new_n743), .A2(new_n744), .B1(new_n726), .B2(new_n725), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT31), .B(G11), .ZN(new_n748));
  NOR2_X1   g323(.A1(KEYINPUT96), .A2(G28), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(KEYINPUT96), .A2(G28), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n750), .A2(new_n751), .B1(KEYINPUT97), .B2(KEYINPUT30), .ZN(new_n752));
  NOR2_X1   g327(.A1(KEYINPUT97), .A2(KEYINPUT30), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n752), .B2(new_n753), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n748), .B1(new_n755), .B2(new_n757), .C1(new_n647), .C2(new_n728), .ZN(new_n758));
  INV_X1    g333(.A(G1961), .ZN(new_n759));
  NOR2_X1   g334(.A1(G5), .A2(G16), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT98), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n573), .A2(new_n532), .A3(new_n531), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(new_n709), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n758), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n739), .A2(G19), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n545), .B2(new_n739), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G1341), .Z(new_n767));
  NOR2_X1   g342(.A1(G29), .A2(G33), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT25), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n461), .A2(G139), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n494), .A2(G127), .ZN(new_n775));
  NAND2_X1  g350(.A1(G115), .A2(G2104), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n462), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n768), .B1(new_n778), .B2(G29), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(G2072), .Z(new_n780));
  NAND3_X1  g355(.A1(new_n764), .A2(new_n767), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n756), .A2(G32), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT92), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G141), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n494), .A2(new_n462), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n475), .A2(G129), .ZN(new_n789));
  NAND3_X1  g364(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(KEYINPUT26), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(KEYINPUT26), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n789), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n794));
  OR3_X1    g369(.A1(new_n788), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n788), .B2(new_n793), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n782), .B1(new_n797), .B2(new_n756), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT27), .B(G1996), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT94), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n763), .A2(new_n759), .ZN(new_n802));
  NOR2_X1   g377(.A1(G168), .A2(new_n709), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n709), .B2(G21), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT95), .B(G1966), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n804), .B2(new_n805), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n781), .A2(new_n801), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n729), .A2(G27), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G164), .B2(new_n729), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT99), .B(G2078), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n728), .A2(G26), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT28), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n475), .A2(G128), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n462), .A2(G116), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n817));
  INV_X1    g392(.A(G140), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n815), .B1(new_n816), .B2(new_n817), .C1(new_n818), .C2(new_n787), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(KEYINPUT91), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(KEYINPUT91), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n814), .B1(new_n822), .B2(G29), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G2067), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n808), .A2(new_n812), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(G160), .A2(G29), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT24), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(G34), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(G34), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n728), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G2084), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n720), .A2(G20), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT23), .Z(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G299), .B2(G16), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(G1956), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n709), .A2(G4), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n618), .B2(new_n709), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G1348), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n729), .A2(G35), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G162), .B2(new_n729), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT29), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(G2090), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n800), .A2(new_n798), .B1(new_n843), .B2(G2090), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n832), .A2(new_n840), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n747), .A2(new_n825), .A3(new_n846), .ZN(G311));
  INV_X1    g422(.A(G311), .ZN(G150));
  NAND2_X1  g423(.A1(new_n618), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT38), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n509), .A2(new_n510), .A3(G93), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n510), .A2(G55), .A3(G543), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT101), .ZN(new_n853));
  AOI21_X1  g428(.A(KEYINPUT101), .B1(new_n851), .B2(new_n852), .ZN(new_n854));
  OAI21_X1  g429(.A(G67), .B1(new_n502), .B2(new_n501), .ZN(new_n855));
  NAND2_X1  g430(.A1(G80), .A2(G543), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT100), .B1(new_n857), .B2(G651), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n859));
  AOI211_X1 g434(.A(new_n859), .B(new_n534), .C1(new_n855), .C2(new_n856), .ZN(new_n860));
  OAI22_X1  g435(.A1(new_n853), .A2(new_n854), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n540), .A2(new_n544), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n851), .A2(new_n852), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT101), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n857), .A2(G651), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n859), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n857), .A2(KEYINPUT100), .A3(G651), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n868), .A2(new_n872), .A3(new_n545), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n863), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n850), .B(new_n874), .Z(new_n875));
  AND2_X1   g450(.A1(new_n875), .A2(KEYINPUT39), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(KEYINPUT39), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n876), .A2(new_n877), .A3(G860), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n861), .A2(G860), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT37), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n878), .A2(new_n880), .ZN(G145));
  XNOR2_X1  g456(.A(new_n797), .B(new_n822), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n493), .A2(new_n496), .ZN(new_n883));
  INV_X1    g458(.A(new_n485), .ZN(new_n884));
  NOR2_X1   g459(.A1(KEYINPUT67), .A2(G114), .ZN(new_n885));
  OAI21_X1  g460(.A(G2105), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n487), .ZN(new_n887));
  AOI22_X1  g462(.A1(G126), .A2(new_n475), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n882), .B(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n778), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n882), .A2(new_n889), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n882), .A2(new_n889), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n778), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n475), .A2(G130), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n462), .A2(G118), .ZN(new_n898));
  OAI21_X1  g473(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(G142), .B2(new_n461), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n637), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n735), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT103), .B1(new_n896), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n906));
  AOI211_X1 g481(.A(new_n906), .B(new_n903), .C1(new_n892), .C2(new_n895), .ZN(new_n907));
  OAI22_X1  g482(.A1(new_n905), .A2(new_n907), .B1(new_n896), .B2(new_n904), .ZN(new_n908));
  XNOR2_X1  g483(.A(G160), .B(KEYINPUT102), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(G162), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(new_n647), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n904), .B1(new_n896), .B2(KEYINPUT104), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(KEYINPUT104), .B2(new_n896), .ZN(new_n914));
  INV_X1    g489(.A(new_n911), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n914), .B(new_n915), .C1(new_n905), .C2(new_n907), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n912), .A2(KEYINPUT40), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT40), .B1(new_n912), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(G395));
  NAND2_X1  g494(.A1(new_n861), .A2(new_n620), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n632), .B(new_n874), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n618), .A2(G299), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n609), .A2(new_n617), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n625), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n625), .A2(new_n923), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n924), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n625), .A2(new_n923), .A3(KEYINPUT105), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT105), .B1(new_n625), .B2(new_n923), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n932), .A2(new_n933), .A3(new_n928), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n931), .B1(new_n934), .B2(KEYINPUT41), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n927), .B1(new_n921), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G48), .ZN(new_n937));
  INV_X1    g512(.A(G86), .ZN(new_n938));
  OAI22_X1  g513(.A1(new_n541), .A2(new_n937), .B1(new_n503), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n509), .A2(G61), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n534), .B1(new_n940), .B2(new_n593), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n602), .B(new_n603), .C1(new_n939), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n509), .A2(G60), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n534), .B1(new_n943), .B2(new_n600), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n510), .A2(G47), .A3(G543), .ZN(new_n945));
  INV_X1    g520(.A(G85), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(new_n503), .B2(new_n946), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n595), .B(new_n596), .C1(new_n944), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n581), .B(G288), .C1(new_n582), .C2(new_n583), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n506), .A2(new_n514), .ZN(new_n952));
  AOI21_X1  g527(.A(G288), .B1(new_n952), .B2(new_n581), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n949), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(G303), .A2(new_n711), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n955), .A2(new_n950), .A3(new_n942), .A4(new_n948), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT42), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n951), .A2(new_n953), .A3(new_n949), .ZN(new_n959));
  AOI22_X1  g534(.A1(new_n955), .A2(new_n950), .B1(new_n942), .B2(new_n948), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n954), .A2(new_n956), .A3(KEYINPUT106), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n957), .B1(new_n963), .B2(KEYINPUT42), .ZN(new_n964));
  XOR2_X1   g539(.A(new_n936), .B(new_n964), .Z(new_n965));
  OAI21_X1  g540(.A(new_n920), .B1(new_n965), .B2(new_n620), .ZN(G295));
  OAI21_X1  g541(.A(new_n920), .B1(new_n965), .B2(new_n620), .ZN(G331));
  INV_X1    g542(.A(new_n963), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n569), .A2(G168), .A3(new_n575), .ZN(new_n969));
  NAND3_X1  g544(.A1(G171), .A2(G286), .A3(KEYINPUT107), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n762), .B2(G168), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n874), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(new_n863), .A3(new_n873), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n974), .A2(new_n925), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n974), .A2(KEYINPUT109), .A3(new_n976), .A4(new_n925), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n974), .A2(new_n976), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT105), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n618), .B2(G299), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n625), .A2(new_n923), .A3(KEYINPUT105), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n922), .A3(new_n985), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n986), .A2(new_n929), .B1(new_n924), .B2(new_n930), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n982), .A2(new_n987), .A3(KEYINPUT108), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n974), .A2(new_n976), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n935), .B2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n968), .B(new_n981), .C1(new_n988), .C2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G37), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT108), .B1(new_n982), .B2(new_n987), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n935), .A2(new_n989), .A3(new_n990), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n968), .B1(new_n997), .B2(new_n981), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n994), .A2(new_n998), .A3(KEYINPUT43), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n929), .B1(new_n974), .B2(new_n976), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n986), .A2(new_n1002), .B1(new_n961), .B2(new_n962), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n926), .B1(new_n982), .B2(new_n929), .ZN(new_n1004));
  AOI21_X1  g579(.A(G37), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1001), .B1(new_n992), .B2(new_n1005), .ZN(new_n1006));
  OR3_X1    g581(.A1(new_n999), .A2(new_n1000), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT43), .B1(new_n994), .B2(new_n998), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n992), .A2(new_n1005), .A3(new_n1009), .A4(new_n1001), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n992), .A2(new_n1005), .A3(new_n1001), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1008), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n1000), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1014), .B1(new_n1013), .B2(new_n1000), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1007), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT112), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1019), .B(new_n1007), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(G397));
  XNOR2_X1  g596(.A(new_n822), .B(G2067), .ZN(new_n1022));
  INV_X1    g597(.A(G1996), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n797), .A2(new_n1023), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n889), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n463), .A2(G101), .ZN(new_n1028));
  INV_X1    g603(.A(G137), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1028), .B1(new_n787), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n494), .A2(G125), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n462), .B1(new_n1031), .B2(new_n467), .ZN(new_n1032));
  INV_X1    g607(.A(G40), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1027), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT113), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(G1996), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1025), .A2(new_n1037), .B1(new_n797), .B2(new_n1038), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n735), .A2(new_n737), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n735), .A2(new_n737), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1036), .ZN(new_n1044));
  XNOR2_X1  g619(.A(G290), .B(G1986), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT63), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  NOR2_X1   g624(.A1(G166), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1050), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n490), .A2(new_n491), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n883), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n1026), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n464), .A2(new_n469), .A3(G40), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G2090), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1384), .B1(new_n883), .B2(new_n888), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1063), .B1(KEYINPUT45), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(G1384), .B1(new_n1059), .B2(new_n883), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1068), .B1(KEYINPUT45), .B2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1065), .A2(new_n1066), .B1(new_n1070), .B2(new_n723), .ZN(new_n1071));
  OAI211_X1 g646(.A(KEYINPUT119), .B(new_n1058), .C1(new_n1071), .C2(new_n1049), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT45), .B1(new_n1060), .B2(new_n1026), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1067), .A2(KEYINPUT45), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n1034), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n723), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1062), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1049), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1073), .B1(new_n1079), .B2(new_n1057), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1049), .B1(new_n1034), .B2(new_n1067), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n711), .A2(G1976), .ZN(new_n1082));
  INV_X1    g657(.A(G1976), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT52), .B1(G288), .B2(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT52), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT116), .A4(G1981), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT117), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n595), .A2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1093), .A2(G1981), .B1(new_n595), .B2(new_n596), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT49), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(G1981), .B1(new_n941), .B2(KEYINPUT116), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G305), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT49), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1097), .A2(KEYINPUT117), .A3(new_n1098), .A4(new_n1090), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1095), .A2(new_n1081), .A3(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1081), .A2(new_n1088), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1089), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1077), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1063), .B1(new_n1061), .B2(new_n1067), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(G2090), .ZN(new_n1108));
  OAI211_X1 g683(.A(G8), .B(new_n1057), .C1(new_n1104), .C2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1072), .A2(new_n1080), .A3(new_n1103), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G2084), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1107), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1060), .A2(KEYINPUT45), .A3(new_n1026), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1063), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1114));
  AOI21_X1  g689(.A(G1966), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1111), .A2(new_n1112), .B1(new_n1115), .B2(KEYINPUT120), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1115), .A2(KEYINPUT120), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1049), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(G168), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1048), .B1(new_n1110), .B2(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1121));
  OAI21_X1  g696(.A(G8), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1048), .B1(new_n1122), .B2(new_n1058), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1121), .A2(G168), .A3(new_n1118), .A4(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1100), .A2(new_n1083), .A3(new_n711), .ZN(new_n1126));
  NOR2_X1   g701(.A1(G305), .A2(G1981), .ZN(new_n1127));
  XOR2_X1   g702(.A(new_n1127), .B(KEYINPUT118), .Z(new_n1128));
  OR2_X1    g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1109), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1081), .A2(new_n1129), .B1(new_n1130), .B2(new_n1103), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1125), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n625), .B(KEYINPUT57), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT56), .B(G2072), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1074), .A2(new_n1076), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(G1956), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1134), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1137), .A2(new_n1134), .A3(new_n1138), .ZN(new_n1140));
  AOI21_X1  g715(.A(G1348), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1034), .A2(new_n1067), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(G2067), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n618), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1139), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(KEYINPUT121), .B(new_n1139), .C1(new_n1140), .C2(new_n1144), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1068), .B(new_n1135), .C1(KEYINPUT45), .C2(new_n1069), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1133), .B(new_n1150), .C1(new_n1065), .C2(G1956), .ZN(new_n1151));
  AOI21_X1  g726(.A(KEYINPUT61), .B1(new_n1139), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1152), .A2(KEYINPUT123), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n1154));
  AOI211_X1 g729(.A(new_n1154), .B(KEYINPUT61), .C1(new_n1139), .C2(new_n1151), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1139), .A2(new_n1151), .A3(KEYINPUT61), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1141), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1143), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1158), .A2(new_n1159), .A3(new_n618), .A4(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1158), .A2(new_n923), .A3(new_n1160), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1159), .B1(new_n1163), .B2(new_n1144), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1068), .B(new_n1023), .C1(KEYINPUT45), .C2(new_n1069), .ZN(new_n1165));
  XOR2_X1   g740(.A(KEYINPUT58), .B(G1341), .Z(new_n1166));
  NAND2_X1  g741(.A1(new_n1142), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT59), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n545), .B1(KEYINPUT122), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1168), .A2(new_n1171), .B1(KEYINPUT122), .B2(new_n1169), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1169), .A2(KEYINPUT122), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n1170), .B(new_n1173), .C1(new_n1165), .C2(new_n1167), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1162), .A2(new_n1164), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1149), .B1(new_n1156), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(G2078), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1068), .B(new_n1178), .C1(KEYINPUT45), .C2(new_n1069), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT53), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1113), .A2(new_n1114), .A3(KEYINPUT53), .A4(new_n1178), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1061), .B1(new_n1060), .B2(new_n1026), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1034), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n759), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1181), .A2(G301), .A3(new_n1182), .A4(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(KEYINPUT54), .ZN(new_n1187));
  AOI211_X1 g762(.A(new_n1180), .B(G2078), .C1(new_n1067), .C2(KEYINPUT45), .ZN(new_n1188));
  AOI22_X1  g763(.A1(new_n1179), .A2(new_n1180), .B1(new_n1114), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1185), .A2(KEYINPUT126), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1107), .A2(new_n1191), .A3(new_n759), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1187), .B1(G171), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1194), .A2(new_n1110), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1185), .A2(new_n1182), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n576), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI211_X1 g775(.A(KEYINPUT125), .B(new_n576), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1189), .A2(new_n1190), .A3(G301), .A4(new_n1192), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT54), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1195), .A2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1177), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1209));
  OAI211_X1 g784(.A(new_n1208), .B(G8), .C1(new_n1209), .C2(G286), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT51), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g787(.A1(G168), .A2(new_n1049), .ZN(new_n1213));
  OAI211_X1 g788(.A(new_n1208), .B(KEYINPUT51), .C1(new_n1118), .C2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1209), .A2(new_n1213), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1132), .B1(new_n1207), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1217), .A2(KEYINPUT62), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1216), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1220), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1221));
  INV_X1    g796(.A(KEYINPUT62), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1110), .B1(new_n1201), .B2(new_n1200), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1219), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1047), .B1(new_n1218), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1227));
  OAI21_X1  g802(.A(new_n1227), .B1(G2067), .B2(new_n822), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1228), .A2(new_n1037), .ZN(new_n1229));
  INV_X1    g804(.A(new_n797), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1037), .B1(new_n1022), .B2(new_n1230), .ZN(new_n1231));
  XOR2_X1   g806(.A(new_n1038), .B(KEYINPUT46), .Z(new_n1232));
  NAND2_X1  g807(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  XNOR2_X1  g808(.A(new_n1233), .B(KEYINPUT47), .ZN(new_n1234));
  NOR3_X1   g809(.A1(new_n1036), .A2(G1986), .A3(G290), .ZN(new_n1235));
  XOR2_X1   g810(.A(new_n1235), .B(KEYINPUT48), .Z(new_n1236));
  NAND3_X1  g811(.A1(new_n1039), .A2(new_n1042), .A3(new_n1236), .ZN(new_n1237));
  NAND3_X1  g812(.A1(new_n1229), .A2(new_n1234), .A3(new_n1237), .ZN(new_n1238));
  OAI21_X1  g813(.A(KEYINPUT127), .B1(new_n1226), .B2(new_n1238), .ZN(new_n1239));
  AND2_X1   g814(.A1(new_n1125), .A2(new_n1131), .ZN(new_n1240));
  AND2_X1   g815(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1241));
  XNOR2_X1  g816(.A(new_n1152), .B(KEYINPUT123), .ZN(new_n1242));
  NOR2_X1   g817(.A1(new_n1175), .A2(new_n1164), .ZN(new_n1243));
  AND2_X1   g818(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1244));
  NAND2_X1  g819(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g820(.A(new_n1241), .B1(new_n1242), .B2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g821(.A1(new_n1246), .A2(new_n1205), .A3(new_n1195), .ZN(new_n1247));
  OAI21_X1  g822(.A(new_n1240), .B1(new_n1247), .B2(new_n1221), .ZN(new_n1248));
  OAI21_X1  g823(.A(new_n1224), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1249));
  AOI211_X1 g824(.A(KEYINPUT62), .B(new_n1220), .C1(new_n1212), .C2(new_n1214), .ZN(new_n1250));
  NOR2_X1   g825(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g826(.A(new_n1046), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1253));
  INV_X1    g828(.A(new_n1238), .ZN(new_n1254));
  NAND3_X1  g829(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g830(.A1(new_n1239), .A2(new_n1255), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g831(.A1(new_n912), .A2(new_n916), .ZN(new_n1258));
  INV_X1    g832(.A(G319), .ZN(new_n1259));
  NOR3_X1   g833(.A1(G401), .A2(new_n1259), .A3(G227), .ZN(new_n1260));
  AND4_X1   g834(.A1(new_n707), .A2(new_n1258), .A3(new_n1013), .A4(new_n1260), .ZN(G308));
  NAND4_X1  g835(.A1(new_n707), .A2(new_n1258), .A3(new_n1013), .A4(new_n1260), .ZN(G225));
endmodule


