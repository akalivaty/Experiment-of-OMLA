//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1306, new_n1307, new_n1308, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT65), .Z(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n203), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  INV_X1    g0026(.A(G77), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G107), .ZN(new_n229));
  INV_X1    g0029(.A(G264), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n211), .B1(new_n225), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  INV_X1    g0033(.A(KEYINPUT1), .ZN(new_n234));
  OR2_X1    g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  AND3_X1   g0036(.A1(new_n219), .A2(new_n235), .A3(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT67), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n255), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n254), .A2(new_n256), .A3(new_n215), .A4(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G1), .ZN(new_n260));
  OAI21_X1  g0060(.A(G97), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G97), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT74), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n261), .A2(KEYINPUT74), .A3(new_n263), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(new_n227), .ZN(new_n271));
  XNOR2_X1  g0071(.A(G97), .B(G107), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT6), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n273), .A2(new_n262), .A3(G107), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n271), .B1(new_n277), .B2(G20), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(KEYINPUT7), .B1(new_n282), .B2(new_n209), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT7), .ZN(new_n284));
  AOI211_X1 g0084(.A(new_n284), .B(G20), .C1(new_n279), .C2(new_n281), .ZN(new_n285));
  OAI21_X1  g0085(.A(G107), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n278), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n254), .A2(new_n215), .A3(new_n256), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n268), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G169), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G1), .A3(G13), .ZN(new_n293));
  AND2_X1   g0093(.A1(KEYINPUT4), .A2(G244), .ZN(new_n294));
  INV_X1    g0094(.A(G1698), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n279), .A2(new_n281), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G283), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT4), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT72), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n259), .B2(KEYINPUT3), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n280), .A2(KEYINPUT72), .A3(G33), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n228), .A2(G1698), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n301), .A2(new_n302), .A3(new_n303), .A4(new_n279), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n298), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n279), .A2(new_n281), .A3(G250), .A4(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT75), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT3), .B(G33), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n309), .A2(KEYINPUT75), .A3(G250), .A4(G1698), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n293), .B1(new_n305), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G45), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(G1), .ZN(new_n314));
  AND2_X1   g0114(.A1(KEYINPUT5), .A2(G41), .ZN(new_n315));
  NOR2_X1   g0115(.A1(KEYINPUT5), .A2(G41), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n317), .A2(G257), .A3(new_n293), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT5), .B(G41), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n319), .A2(G274), .A3(new_n293), .A4(new_n314), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT76), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n318), .A2(KEYINPUT76), .A3(new_n320), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n291), .B1(new_n312), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n304), .A2(new_n299), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n311), .A2(new_n327), .A3(new_n297), .A4(new_n296), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G179), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n318), .A2(KEYINPUT76), .A3(new_n320), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT76), .B1(new_n318), .B2(new_n320), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n330), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n290), .A2(new_n326), .A3(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(G200), .B1(new_n312), .B2(new_n325), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n267), .A2(new_n266), .B1(new_n287), .B2(new_n288), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n330), .A2(G190), .A3(new_n334), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT77), .ZN(new_n342));
  INV_X1    g0142(.A(G58), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(new_n221), .ZN(new_n344));
  OAI21_X1  g0144(.A(G20), .B1(new_n344), .B2(new_n202), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n269), .A2(G159), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n301), .A2(new_n279), .A3(new_n302), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(new_n284), .A3(new_n209), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G68), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n284), .B1(new_n349), .B2(new_n209), .ZN(new_n352));
  OAI211_X1 g0152(.A(KEYINPUT16), .B(new_n348), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT16), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n284), .B1(new_n309), .B2(G20), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n221), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n354), .B1(new_n357), .B2(new_n347), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(new_n288), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT8), .B(G58), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n257), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n209), .A2(G1), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n254), .A2(new_n215), .A3(new_n256), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(KEYINPUT69), .A3(new_n257), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT69), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n258), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n362), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n361), .B1(new_n367), .B2(new_n360), .ZN(new_n368));
  INV_X1    g0168(.A(G200), .ZN(new_n369));
  NOR2_X1   g0169(.A1(G223), .A2(G1698), .ZN(new_n370));
  INV_X1    g0170(.A(G226), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(G1698), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n372), .A2(new_n279), .A3(new_n301), .A4(new_n302), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G87), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n293), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G41), .ZN(new_n376));
  AOI21_X1  g0176(.A(G1), .B1(new_n376), .B2(new_n313), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(new_n293), .A3(G274), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n293), .A2(G232), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n369), .B1(new_n375), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n371), .A2(G1698), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(G223), .B2(G1698), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n374), .B1(new_n349), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n329), .ZN(new_n386));
  INV_X1    g0186(.A(G190), .ZN(new_n387));
  INV_X1    g0187(.A(new_n381), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n382), .A2(KEYINPUT73), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT73), .B1(new_n382), .B2(new_n389), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n359), .B(new_n368), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT17), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT73), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n375), .A2(G190), .A3(new_n381), .ZN(new_n396));
  AOI21_X1  g0196(.A(G200), .B1(new_n386), .B2(new_n388), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n382), .A2(KEYINPUT73), .A3(new_n389), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(G68), .B1(new_n283), .B2(new_n285), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n348), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n363), .B1(new_n402), .B2(new_n354), .ZN(new_n403));
  INV_X1    g0203(.A(new_n362), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n258), .A2(new_n365), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n258), .A2(new_n365), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n360), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n403), .A2(new_n353), .B1(new_n409), .B2(new_n361), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n400), .A2(new_n410), .A3(KEYINPUT17), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n394), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  OAI21_X1  g0213(.A(G169), .B1(new_n375), .B2(new_n381), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n386), .A2(G179), .A3(new_n388), .ZN(new_n415));
  AOI221_X4 g0215(.A(new_n413), .B1(new_n414), .B2(new_n415), .C1(new_n359), .C2(new_n368), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n359), .A2(new_n368), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n415), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT18), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n412), .A2(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n269), .A2(G50), .B1(G20), .B2(new_n221), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n259), .A2(G20), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n422), .B1(new_n424), .B2(new_n227), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n288), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT11), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n257), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n221), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT12), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n258), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(G68), .A3(new_n404), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n427), .B2(new_n426), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n371), .A2(new_n295), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n295), .A2(G232), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n309), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G97), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n329), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT13), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n293), .A2(new_n379), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G274), .ZN(new_n447));
  INV_X1    g0247(.A(new_n215), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n447), .B1(new_n448), .B2(new_n292), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n446), .A2(G238), .B1(new_n449), .B2(new_n377), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n443), .A2(new_n444), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n293), .B1(new_n440), .B2(new_n441), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n378), .B1(new_n222), .B2(new_n445), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT13), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT14), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(G169), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n451), .A2(G179), .A3(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n456), .B1(new_n455), .B2(G169), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n437), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n455), .A2(G200), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(new_n436), .C1(new_n387), .C2(new_n455), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G20), .A2(G77), .ZN(new_n464));
  XNOR2_X1  g0264(.A(KEYINPUT15), .B(G87), .ZN(new_n465));
  OAI221_X1 g0265(.A(new_n464), .B1(new_n360), .B2(new_n270), .C1(new_n465), .C2(new_n424), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n288), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n433), .A2(G77), .A3(new_n404), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n429), .A2(new_n227), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n378), .B1(new_n228), .B2(new_n445), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n309), .A2(G238), .A3(G1698), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n309), .A2(G232), .A3(new_n295), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n472), .B(new_n473), .C1(new_n229), .C2(new_n309), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(new_n474), .B2(new_n329), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n470), .B1(new_n476), .B2(G200), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(G190), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n475), .A2(new_n331), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n480), .B(new_n470), .C1(G169), .C2(new_n475), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n421), .A2(new_n461), .A3(new_n463), .A4(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(G50), .B(new_n404), .C1(new_n405), .C2(new_n406), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT68), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n269), .A2(G150), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n486), .C1(new_n360), .C2(new_n424), .ZN(new_n487));
  OAI21_X1  g0287(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n343), .A2(KEYINPUT8), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n343), .A2(KEYINPUT8), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n423), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n485), .B1(new_n492), .B2(new_n486), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n288), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G50), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n429), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n484), .A2(new_n494), .A3(KEYINPUT9), .A4(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT70), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n486), .B1(new_n360), .B2(new_n424), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT68), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(new_n488), .A3(new_n487), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(new_n288), .B1(new_n495), .B2(new_n429), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n503), .A2(KEYINPUT70), .A3(KEYINPUT9), .A4(new_n484), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n378), .B1(new_n371), .B2(new_n445), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n293), .B1(new_n282), .B2(new_n227), .ZN(new_n508));
  NOR2_X1   g0308(.A1(G222), .A2(G1698), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n295), .A2(G223), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n309), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n507), .A2(G190), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n506), .B1(new_n511), .B2(new_n508), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(new_n369), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n503), .A2(new_n484), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT9), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n505), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT10), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT71), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(KEYINPUT71), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n519), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT71), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n505), .A2(new_n518), .A3(new_n525), .A4(KEYINPUT10), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n514), .A2(new_n331), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n516), .B(new_n527), .C1(G169), .C2(new_n514), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n483), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT77), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n336), .A2(new_n340), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n224), .A2(new_n295), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(G257), .B2(new_n295), .ZN(new_n534));
  INV_X1    g0334(.A(G294), .ZN(new_n535));
  OAI22_X1  g0335(.A1(new_n349), .A2(new_n534), .B1(new_n259), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n329), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n329), .B1(new_n314), .B2(new_n319), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G264), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n320), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT85), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n536), .A2(new_n329), .B1(new_n538), .B2(G264), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(KEYINPUT85), .A3(new_n320), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(G169), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n540), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G179), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n229), .A2(G20), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT23), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n550), .A2(KEYINPUT82), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n549), .A2(KEYINPUT23), .ZN(new_n552));
  NAND2_X1  g0352(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G33), .A2(G116), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(G20), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n550), .A2(KEYINPUT82), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n551), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n301), .A2(new_n302), .A3(new_n209), .A4(new_n279), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT22), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n559), .A2(new_n560), .A3(new_n223), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n209), .A2(G87), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n560), .B1(new_n282), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n558), .A2(new_n562), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n551), .A2(new_n566), .A3(new_n556), .A4(new_n557), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n563), .B1(new_n568), .B2(new_n561), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n569), .A3(new_n288), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n258), .A2(new_n229), .A3(new_n260), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT84), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n208), .A2(new_n229), .A3(G13), .A4(G20), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n573), .B(KEYINPUT25), .ZN(new_n574));
  OR3_X1    g0374(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n572), .B1(new_n571), .B2(new_n574), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n570), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n548), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(G190), .B1(new_n542), .B2(new_n544), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n546), .A2(G200), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n577), .B(new_n570), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n532), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n258), .A2(new_n260), .ZN(new_n584));
  INV_X1    g0384(.A(new_n465), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT80), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT19), .B1(new_n423), .B2(G97), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n223), .A2(new_n262), .A3(new_n229), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT78), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT78), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n591), .A2(new_n223), .A3(new_n262), .A4(new_n229), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT19), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n441), .B2(new_n209), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n588), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n301), .A2(new_n279), .A3(new_n302), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT79), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n597), .A2(new_n598), .A3(new_n209), .A4(G68), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT79), .B1(new_n559), .B2(new_n221), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n288), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n585), .A2(new_n257), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n587), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  AOI211_X1 g0405(.A(KEYINPUT80), .B(new_n603), .C1(new_n601), .C2(new_n288), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n586), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n208), .A2(G45), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n293), .A2(G250), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n293), .A2(G274), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(new_n608), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n228), .A2(G1698), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(G238), .B2(G1698), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n554), .B1(new_n349), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n611), .B1(new_n329), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(G169), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n331), .B2(new_n615), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n607), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n387), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(G200), .B2(new_n615), .ZN(new_n620));
  INV_X1    g0420(.A(new_n584), .ZN(new_n621));
  OAI221_X1 g0421(.A(new_n620), .B1(new_n223), .B2(new_n621), .C1(new_n605), .C2(new_n606), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n317), .A2(G270), .A3(new_n293), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n320), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n282), .A2(G303), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n230), .A2(G1698), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(G257), .B2(G1698), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n349), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n625), .B1(new_n329), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n630), .A2(new_n291), .ZN(new_n631));
  AOI21_X1  g0431(.A(G20), .B1(G33), .B2(G283), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n259), .A2(G97), .ZN(new_n633));
  INV_X1    g0433(.A(G116), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n632), .A2(new_n633), .B1(G20), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n288), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT20), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n288), .A2(new_n635), .A3(KEYINPUT20), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n638), .A2(new_n639), .B1(new_n634), .B2(new_n429), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n584), .A2(G116), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT21), .B1(new_n631), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n642), .ZN(new_n645));
  INV_X1    g0445(.A(new_n625), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n629), .A2(new_n329), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G200), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n645), .B(new_n649), .C1(new_n387), .C2(new_n648), .ZN(new_n650));
  INV_X1    g0450(.A(new_n628), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n597), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n293), .B1(new_n652), .B2(new_n626), .ZN(new_n653));
  OAI211_X1 g0453(.A(KEYINPUT21), .B(G169), .C1(new_n653), .C2(new_n625), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n646), .A2(new_n647), .A3(G179), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n656), .A2(KEYINPUT81), .A3(new_n642), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT81), .B1(new_n656), .B2(new_n642), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n644), .B(new_n650), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n623), .A2(new_n659), .ZN(new_n660));
  AND4_X1   g0460(.A1(new_n342), .A2(new_n530), .A3(new_n583), .A4(new_n660), .ZN(G372));
  INV_X1    g0461(.A(new_n470), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n662), .B1(new_n291), .B2(new_n476), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n463), .A2(new_n480), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n412), .B1(new_n461), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g0465(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n416), .B2(new_n419), .ZN(new_n668));
  INV_X1    g0468(.A(new_n418), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n413), .B1(new_n410), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n417), .A2(KEYINPUT18), .A3(new_n418), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n671), .A3(new_n666), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n524), .B(new_n526), .C1(new_n665), .C2(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n674), .A2(new_n528), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n621), .A2(new_n223), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n602), .A2(new_n604), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT80), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n602), .A2(new_n587), .A3(new_n604), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n680), .A2(new_n620), .B1(new_n607), .B2(new_n617), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n656), .A2(new_n642), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n579), .A2(new_n682), .A3(new_n644), .ZN(new_n683));
  INV_X1    g0483(.A(new_n341), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n681), .A2(new_n683), .A3(new_n684), .A4(new_n582), .ZN(new_n685));
  INV_X1    g0485(.A(new_n336), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT26), .B1(new_n681), .B2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n618), .A2(new_n622), .A3(KEYINPUT26), .A4(new_n686), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n618), .B(new_n685), .C1(new_n687), .C2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n530), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n675), .A2(new_n691), .ZN(G369));
  NAND3_X1  g0492(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g0496(.A(KEYINPUT88), .B(G343), .Z(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n642), .B(new_n698), .C1(new_n643), .C2(new_n656), .ZN(new_n699));
  INV_X1    g0499(.A(new_n698), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n645), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n699), .B1(new_n659), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT89), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(KEYINPUT89), .A3(G330), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n579), .A2(new_n582), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n578), .A2(new_n698), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n548), .A2(new_n578), .A3(new_n698), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT81), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n682), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n656), .A2(KEYINPUT81), .A3(new_n642), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n643), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n698), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n709), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n579), .B2(new_n698), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n715), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT90), .Z(G399));
  NOR2_X1   g0524(.A1(new_n593), .A2(G116), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT91), .ZN(new_n726));
  INV_X1    g0526(.A(new_n212), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G41), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(G1), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n217), .B2(new_n729), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n660), .A2(new_n342), .A3(new_n583), .A4(new_n700), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT92), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n615), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n330), .A2(new_n334), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n630), .A2(G179), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n735), .A2(new_n736), .A3(new_n540), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n543), .A2(new_n615), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n655), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n740), .A2(KEYINPUT30), .A3(new_n330), .A4(new_n334), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT30), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n630), .A2(new_n615), .A3(G179), .A4(new_n543), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n742), .B1(new_n736), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n738), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n698), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT31), .B1(new_n745), .B2(new_n698), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT93), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n745), .A2(new_n698), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT31), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT93), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(new_n753), .A3(new_n746), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n733), .A2(new_n749), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT29), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n690), .A2(new_n757), .A3(new_n700), .ZN(new_n758));
  INV_X1    g0558(.A(new_n618), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n618), .A2(new_n622), .A3(new_n686), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT26), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n759), .B1(new_n762), .B2(new_n688), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n719), .A2(new_n579), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n764), .A2(new_n684), .A3(new_n582), .A4(new_n681), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n698), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n756), .B(new_n758), .C1(new_n757), .C2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n732), .B1(new_n768), .B2(G1), .ZN(G364));
  AND2_X1   g0569(.A1(new_n209), .A2(G13), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n208), .B1(new_n770), .B2(G45), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n728), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n708), .B(new_n774), .C1(G330), .C2(new_n702), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n212), .A2(new_n309), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n776), .A2(new_n206), .B1(G116), .B2(new_n212), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n727), .A2(new_n597), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n313), .B2(new_n218), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n248), .A2(G45), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n215), .B1(G20), .B2(new_n291), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n773), .B1(new_n782), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n209), .A2(new_n331), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G190), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n790), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n793), .A2(new_n387), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n309), .B1(new_n227), .B2(new_n792), .C1(new_n795), .C2(new_n343), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n793), .A2(new_n387), .A3(new_n369), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(KEYINPUT94), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n797), .A2(KEYINPUT94), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n796), .B1(new_n802), .B2(G50), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n209), .A2(G179), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n804), .A2(G190), .A3(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n223), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n804), .A2(new_n387), .A3(G200), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n806), .B1(G107), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n804), .A2(new_n791), .ZN(new_n810));
  INV_X1    g0610(.A(G159), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT32), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n803), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n387), .A2(G179), .A3(G200), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n209), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n262), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n793), .A2(new_n369), .A3(G190), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(G68), .B2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT95), .Z(new_n820));
  NAND2_X1  g0620(.A1(new_n802), .A2(G326), .ZN(new_n821));
  XNOR2_X1  g0621(.A(KEYINPUT33), .B(G317), .ZN(new_n822));
  INV_X1    g0622(.A(new_n792), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n818), .A2(new_n822), .B1(new_n823), .B2(G311), .ZN(new_n824));
  INV_X1    g0624(.A(new_n810), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n794), .A2(G322), .B1(G329), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n816), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n827), .A2(G294), .B1(new_n808), .B2(G283), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n821), .A2(new_n824), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G303), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n282), .B1(new_n805), .B2(new_n830), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT96), .Z(new_n832));
  OAI22_X1  g0632(.A1(new_n814), .A2(new_n820), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n833), .A2(KEYINPUT97), .ZN(new_n834));
  INV_X1    g0634(.A(new_n786), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n833), .B2(KEYINPUT97), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n789), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n785), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n837), .B1(new_n702), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n775), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G396));
  INV_X1    g0641(.A(KEYINPUT99), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n663), .A2(new_n842), .A3(new_n480), .A4(new_n698), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT99), .B1(new_n481), .B2(new_n700), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n479), .B(new_n481), .C1(new_n662), .C2(new_n700), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n690), .B2(new_n700), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n700), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n763), .B2(new_n685), .ZN(new_n850));
  OR2_X1    g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n756), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n773), .B1(new_n851), .B2(new_n756), .ZN(new_n854));
  INV_X1    g0654(.A(new_n847), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n783), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n786), .A2(new_n783), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n773), .B1(G77), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n794), .A2(G143), .B1(G159), .B2(new_n823), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n802), .A2(G137), .B1(G150), .B2(new_n818), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT98), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n862), .A2(KEYINPUT98), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n867), .A2(KEYINPUT34), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n816), .A2(new_n343), .B1(new_n807), .B2(new_n221), .ZN(new_n869));
  INV_X1    g0669(.A(G132), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n597), .B1(new_n870), .B2(new_n810), .ZN(new_n871));
  INV_X1    g0671(.A(new_n805), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n869), .B(new_n871), .C1(G50), .C2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n867), .B2(KEYINPUT34), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n309), .B(new_n817), .C1(G294), .C2(new_n794), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n875), .B1(new_n223), .B2(new_n807), .C1(new_n229), .C2(new_n805), .ZN(new_n876));
  AOI22_X1  g0676(.A1(G116), .A2(new_n823), .B1(new_n825), .B2(G311), .ZN(new_n877));
  INV_X1    g0677(.A(G283), .ZN(new_n878));
  INV_X1    g0678(.A(new_n818), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n877), .B1(new_n878), .B2(new_n879), .C1(new_n801), .C2(new_n830), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n868), .A2(new_n874), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n859), .B1(new_n881), .B2(new_n786), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n853), .A2(new_n854), .B1(new_n856), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(G384));
  OR2_X1    g0684(.A1(new_n277), .A2(KEYINPUT35), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n277), .A2(KEYINPUT35), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n885), .A2(G116), .A3(new_n216), .A4(new_n886), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT36), .Z(new_n888));
  OR3_X1    g0688(.A1(new_n217), .A2(new_n227), .A3(new_n344), .ZN(new_n889));
  INV_X1    g0689(.A(new_n201), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(G68), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n208), .B(G13), .C1(new_n889), .C2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n353), .A2(new_n288), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT7), .B1(new_n597), .B2(G20), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(G68), .A3(new_n350), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT16), .B1(new_n897), .B2(new_n348), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n368), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n696), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n400), .A2(new_n410), .A3(KEYINPUT17), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT17), .B1(new_n400), .B2(new_n410), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n670), .A2(new_n671), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n696), .B1(new_n359), .B2(new_n368), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n417), .A2(new_n418), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n392), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT37), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n899), .A2(new_n418), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n392), .A2(new_n901), .A3(new_n913), .A4(KEYINPUT37), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n894), .B1(new_n906), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n901), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n412), .B2(new_n420), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n392), .A2(KEYINPUT37), .A3(new_n901), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n919), .A2(new_n913), .B1(new_n910), .B2(new_n911), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(new_n920), .A3(KEYINPUT38), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n437), .A2(new_n698), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n461), .A2(new_n463), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n923), .B1(new_n461), .B2(new_n463), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n481), .A2(new_n698), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n922), .B(new_n927), .C1(new_n850), .C2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n673), .A2(new_n696), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n392), .A2(new_n908), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT37), .B1(new_n932), .B2(KEYINPUT86), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n907), .B1(new_n410), .B2(new_n400), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT102), .B1(new_n934), .B2(new_n909), .ZN(new_n935));
  AND4_X1   g0735(.A1(KEYINPUT102), .A2(new_n392), .A3(new_n909), .A4(new_n908), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT86), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n911), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT102), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n910), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(KEYINPUT102), .A3(new_n909), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n668), .A2(new_n672), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n908), .B1(new_n945), .B2(new_n904), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n894), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT39), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(new_n948), .A3(new_n921), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n906), .A2(new_n915), .A3(new_n894), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT38), .B1(new_n918), .B2(new_n920), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT39), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT101), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT101), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n922), .A2(new_n954), .A3(KEYINPUT39), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n949), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n461), .A2(new_n698), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT100), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n931), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n758), .B1(new_n766), .B2(new_n757), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n530), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n962), .A2(new_n675), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n960), .B(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(G330), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n947), .A2(new_n921), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT40), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n847), .B1(new_n924), .B2(new_n925), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n747), .A2(new_n748), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n967), .B(new_n968), .C1(new_n733), .C2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n968), .B1(new_n733), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n922), .A2(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n966), .A2(new_n970), .B1(new_n972), .B2(new_n967), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n733), .A2(new_n969), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n530), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n965), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n973), .B2(new_n975), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n964), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n208), .B2(new_n770), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n964), .A2(new_n977), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n893), .B1(new_n979), .B2(new_n980), .ZN(G367));
  NOR2_X1   g0781(.A1(new_n338), .A2(new_n700), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n341), .A2(new_n982), .B1(new_n336), .B2(new_n700), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT103), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n720), .A2(new_n709), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT42), .Z(new_n987));
  INV_X1    g0787(.A(new_n984), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n336), .B1(new_n988), .B2(new_n579), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n700), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n680), .A2(new_n700), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n759), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n623), .B2(new_n991), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n987), .A2(new_n990), .B1(KEYINPUT43), .B2(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n715), .A2(new_n984), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n998), .B(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n720), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n985), .B1(new_n714), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n707), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n721), .B1(new_n713), .B2(new_n720), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1005), .A2(new_n705), .A3(new_n706), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n961), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT105), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .A4(new_n756), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1011));
  OAI21_X1  g0811(.A(KEYINPUT105), .B1(new_n767), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n579), .A2(new_n698), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n985), .A2(new_n1013), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n1014), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT45), .B1(new_n1014), .B2(new_n984), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT44), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n1014), .A2(new_n1017), .A3(new_n984), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT44), .B1(new_n988), .B2(new_n722), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1015), .A2(new_n1016), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT104), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n715), .A2(new_n1021), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1010), .B(new_n1012), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n768), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n728), .B(KEYINPUT41), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n771), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1001), .A2(new_n1029), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n787), .B1(new_n212), .B2(new_n465), .C1(new_n779), .C2(new_n244), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n802), .A2(G143), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n309), .B1(new_n879), .B2(new_n811), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G58), .B2(new_n872), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n807), .A2(new_n227), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G68), .B2(new_n827), .ZN(new_n1036));
  INV_X1    g0836(.A(G150), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n795), .A2(new_n1037), .B1(new_n890), .B2(new_n792), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G137), .B2(new_n825), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1032), .A2(new_n1034), .A3(new_n1036), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(G311), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n801), .A2(new_n1041), .B1(new_n830), .B2(new_n795), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT106), .Z(new_n1043));
  NAND2_X1  g0843(.A1(new_n872), .A2(G116), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT46), .ZN(new_n1045));
  INV_X1    g0845(.A(G317), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n792), .A2(new_n878), .B1(new_n810), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G294), .B2(new_n818), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n808), .A2(G97), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n597), .B1(new_n827), .B2(G107), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1045), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1040), .B1(new_n1043), .B2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT47), .Z(new_n1053));
  OAI211_X1 g0853(.A(new_n773), .B(new_n1031), .C1(new_n1053), .C2(new_n835), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT107), .Z(new_n1055));
  OR2_X1    g0855(.A1(new_n993), .A2(new_n838), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1030), .A2(new_n1057), .ZN(G387));
  NAND2_X1  g0858(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n728), .B(KEYINPUT109), .Z(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n767), .B2(new_n1011), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n714), .A2(new_n785), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n778), .B1(new_n241), .B2(new_n313), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n726), .B2(new_n776), .ZN(new_n1066));
  OR3_X1    g0866(.A1(new_n360), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1067));
  OAI21_X1  g0867(.A(KEYINPUT50), .B1(new_n360), .B2(G50), .ZN(new_n1068));
  AOI21_X1  g0868(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n726), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1066), .A2(new_n1070), .B1(new_n229), .B2(new_n727), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n773), .B1(new_n1071), .B2(new_n788), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G311), .A2(new_n818), .B1(new_n794), .B2(G317), .ZN(new_n1073));
  INV_X1    g0873(.A(G322), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1073), .B1(new_n830), .B2(new_n792), .C1(new_n801), .C2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT48), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n827), .A2(G283), .B1(new_n872), .B2(G294), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT49), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n807), .A2(new_n634), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n597), .B(new_n1084), .C1(G326), .C2(new_n825), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n801), .A2(new_n811), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n827), .A2(new_n585), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n805), .A2(new_n227), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1088), .A2(new_n1090), .A3(new_n597), .A4(new_n1049), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n795), .A2(new_n495), .B1(new_n792), .B2(new_n221), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n879), .A2(new_n360), .B1(new_n810), .B2(new_n1037), .ZN(new_n1093));
  NOR4_X1   g0893(.A1(new_n1087), .A2(new_n1091), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT108), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1086), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1072), .B1(new_n1096), .B2(new_n786), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1007), .A2(new_n772), .B1(new_n1064), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1063), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT110), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1063), .A2(KEYINPUT110), .A3(new_n1098), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(G393));
  OAI22_X1  g0903(.A1(new_n801), .A2(new_n1037), .B1(new_n811), .B2(new_n795), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT51), .Z(new_n1105));
  AOI22_X1  g0905(.A1(new_n408), .A2(new_n823), .B1(new_n825), .B2(G143), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n890), .B2(new_n879), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n597), .B1(new_n223), .B2(new_n807), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n816), .A2(new_n227), .B1(new_n805), .B2(new_n221), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n801), .A2(new_n1046), .B1(new_n1041), .B2(new_n795), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT52), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n309), .B1(new_n825), .B2(G322), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n229), .B2(new_n807), .C1(new_n878), .C2(new_n805), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1114), .A2(KEYINPUT111), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n818), .A2(G303), .B1(G294), .B2(new_n823), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n634), .B2(new_n816), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT112), .Z(new_n1118));
  NAND2_X1  g0918(.A1(new_n1114), .A2(KEYINPUT111), .ZN(new_n1119));
  AND4_X1   g0919(.A1(new_n1112), .A2(new_n1115), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n786), .B1(new_n1110), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n778), .A2(new_n251), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n788), .B1(G97), .B2(new_n727), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n774), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1121), .B(new_n1124), .C1(new_n984), .C2(new_n838), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1020), .B(new_n715), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1025), .A2(new_n1060), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1126), .A2(new_n1059), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1125), .B1(new_n771), .B2(new_n1126), .C1(new_n1127), .C2(new_n1128), .ZN(G390));
  INV_X1    g0929(.A(new_n959), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n849), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n928), .B1(new_n690), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1130), .B1(new_n1132), .B2(new_n926), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1133), .A2(new_n949), .A3(new_n953), .A4(new_n955), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n755), .A2(G330), .A3(new_n847), .A4(new_n927), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n959), .B(KEYINPUT113), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n928), .B1(new_n766), .B2(new_n847), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1136), .B(new_n966), .C1(new_n1137), .C2(new_n926), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1134), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n974), .A2(G330), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1140), .A2(new_n968), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT114), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n926), .B1(new_n1140), .B2(new_n855), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1146), .A2(new_n1137), .A3(new_n1135), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n755), .A2(G330), .A3(new_n847), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1141), .B1(new_n926), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1147), .B1(new_n1149), .B2(new_n1132), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1140), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n530), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n962), .A2(new_n675), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1145), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1144), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1144), .A2(new_n1154), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1060), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1144), .A2(new_n772), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT54), .B(G143), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n818), .A2(G137), .B1(new_n823), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n870), .B2(new_n795), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n802), .B2(G128), .ZN(new_n1163));
  INV_X1    g0963(.A(G125), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n309), .B1(new_n810), .B2(new_n1164), .C1(new_n890), .C2(new_n807), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G159), .B2(new_n827), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n805), .A2(new_n1037), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1167), .B(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1163), .A2(new_n1166), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n802), .A2(G283), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n309), .B(new_n806), .C1(G116), .C2(new_n794), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n827), .A2(G77), .B1(new_n808), .B2(G68), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n879), .A2(new_n229), .B1(new_n810), .B2(new_n535), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G97), .B2(new_n823), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n835), .B1(new_n1170), .B2(new_n1176), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n774), .B(new_n1177), .C1(new_n360), .C2(new_n857), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n956), .B2(new_n784), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1158), .A2(KEYINPUT116), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT116), .B1(new_n1158), .B2(new_n1179), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1157), .B1(new_n1180), .B2(new_n1181), .ZN(G378));
  INV_X1    g0982(.A(KEYINPUT118), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n516), .A2(new_n900), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n529), .A2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n524), .A2(new_n526), .A3(new_n528), .A4(new_n1184), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1188), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1183), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1188), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(KEYINPUT118), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n783), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n801), .A2(new_n634), .B1(new_n221), .B2(new_n816), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT117), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n349), .A2(new_n376), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n794), .A2(G107), .B1(new_n585), .B2(new_n823), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n262), .B2(new_n879), .C1(new_n878), .C2(new_n810), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n807), .A2(new_n343), .ZN(new_n1204));
  OR3_X1    g1004(.A1(new_n1203), .A2(new_n1089), .A3(new_n1204), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1200), .A2(new_n1201), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1201), .B(new_n495), .C1(G33), .C2(G41), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(G128), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n1210), .A2(new_n795), .B1(new_n879), .B2(new_n870), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G137), .B2(new_n823), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n827), .A2(G150), .B1(new_n872), .B2(new_n1160), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n1164), .C2(new_n801), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n808), .A2(G159), .ZN(new_n1216));
  AOI211_X1 g1016(.A(G33), .B(G41), .C1(new_n825), .C2(G124), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n1206), .A2(KEYINPUT58), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n786), .B1(new_n1209), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n774), .B1(new_n890), .B2(new_n857), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1198), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n934), .A2(new_n938), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n941), .A2(new_n942), .B1(new_n1225), .B2(KEYINPUT37), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n907), .B1(new_n673), .B2(new_n412), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT38), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n970), .B1(new_n1229), .B2(new_n950), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n972), .A2(new_n967), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(G330), .A3(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(new_n1197), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n973), .B2(G330), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n954), .B1(new_n922), .B2(KEYINPUT39), .ZN(new_n1237));
  AOI211_X1 g1037(.A(KEYINPUT101), .B(new_n948), .C1(new_n916), .C2(new_n921), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1130), .B1(new_n1239), .B2(new_n949), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n1233), .A2(new_n1236), .B1(new_n1240), .B2(new_n931), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT119), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n973), .A2(new_n1244), .A3(G330), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n960), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1241), .A2(new_n1242), .A3(new_n1246), .ZN(new_n1247));
  OAI221_X1 g1047(.A(KEYINPUT119), .B1(new_n1240), .B2(new_n931), .C1(new_n1233), .C2(new_n1236), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1223), .B1(new_n1249), .B2(new_n771), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1153), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1144), .B2(new_n1150), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n960), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n956), .A2(new_n959), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n931), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1243), .A2(new_n1245), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(KEYINPUT57), .B1(new_n1253), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1060), .B1(new_n1252), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT120), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT57), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1141), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1134), .A2(new_n1138), .A3(new_n1135), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n1150), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1153), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1258), .A2(new_n1259), .B1(new_n1260), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1260), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1061), .B1(new_n1268), .B2(new_n1265), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT120), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1250), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(G375));
  NAND2_X1  g1072(.A1(new_n926), .A2(new_n783), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n773), .B1(G68), .B2(new_n858), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n794), .A2(G283), .B1(G303), .B2(new_n825), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n634), .B2(new_n879), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n309), .B(new_n1035), .C1(G107), .C2(new_n823), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1277), .B(new_n1088), .C1(new_n262), .C2(new_n805), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1276), .B(new_n1278), .C1(G294), .C2(new_n802), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT121), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n810), .A2(new_n1210), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n879), .A2(new_n1159), .B1(new_n792), .B2(new_n1037), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1283), .B(new_n1284), .C1(G137), .C2(new_n794), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1204), .A2(new_n349), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1286), .B(KEYINPUT122), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n802), .A2(G132), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n827), .A2(G50), .B1(new_n872), .B2(G159), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1285), .A2(new_n1287), .A3(new_n1288), .A4(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1281), .A2(new_n1282), .A3(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1274), .B1(new_n1291), .B2(new_n786), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1150), .A2(new_n772), .B1(new_n1273), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1027), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1293), .B1(new_n1295), .B2(new_n1296), .ZN(G381));
  NOR3_X1   g1097(.A1(G390), .A2(G381), .A3(G384), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1157), .A2(new_n1158), .A3(new_n1179), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n1001), .A2(new_n1029), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1101), .A2(new_n840), .A3(new_n1102), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1300), .A2(new_n1271), .A3(new_n1301), .A4(new_n1303), .ZN(new_n1304));
  XOR2_X1   g1104(.A(new_n1304), .B(KEYINPUT123), .Z(G407));
  NAND2_X1  g1105(.A1(new_n697), .A2(G213), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1271), .A2(new_n1299), .A3(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(G407), .A2(G213), .A3(new_n1308), .ZN(G409));
  NAND2_X1  g1109(.A1(new_n1296), .A2(KEYINPUT60), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT60), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1311), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1310), .A2(new_n1060), .A3(new_n1294), .A4(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(G384), .B1(new_n1313), .B2(new_n1293), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(G384), .A3(new_n1293), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1315), .A2(G2897), .A3(new_n1307), .A4(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1307), .A2(G2897), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1316), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1318), .B1(new_n1319), .B2(new_n1314), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1250), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1265), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1323));
  OAI22_X1  g1123(.A1(new_n1323), .A2(KEYINPUT57), .B1(new_n1269), .B2(KEYINPUT120), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1325));
  OAI211_X1 g1125(.A(G378), .B(new_n1322), .C1(new_n1324), .C2(new_n1325), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1265), .A2(new_n1247), .A3(new_n1027), .A4(new_n1248), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT124), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n771), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1223), .ZN(new_n1332));
  OAI21_X1  g1132(.A(KEYINPUT125), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n772), .B1(new_n1253), .B2(new_n1256), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT125), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1334), .A2(new_n1335), .A3(new_n1223), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1333), .B(new_n1336), .C1(new_n1327), .C2(new_n1328), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1299), .B1(new_n1330), .B2(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1307), .B1(new_n1326), .B2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT126), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1321), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1323), .A2(KEYINPUT124), .A3(new_n1027), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1342), .A2(new_n1329), .A3(new_n1333), .A4(new_n1336), .ZN(new_n1343));
  AOI22_X1  g1143(.A1(new_n1271), .A2(G378), .B1(new_n1343), .B2(new_n1299), .ZN(new_n1344));
  OAI21_X1  g1144(.A(KEYINPUT126), .B1(new_n1344), .B2(new_n1307), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1341), .A2(new_n1345), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1319), .A2(new_n1314), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1339), .A2(KEYINPUT63), .A3(new_n1347), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1125), .B1(new_n1126), .B2(new_n771), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n840), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1352));
  NOR3_X1   g1152(.A1(new_n1303), .A2(new_n1351), .A3(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(G393), .A2(G396), .ZN(new_n1354));
  AOI21_X1  g1154(.A(G390), .B1(new_n1354), .B2(new_n1302), .ZN(new_n1355));
  OAI21_X1  g1155(.A(G387), .B1(new_n1353), .B2(new_n1355), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1351), .B1(new_n1303), .B2(new_n1352), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1354), .A2(G390), .A3(new_n1302), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1357), .A2(new_n1301), .A3(new_n1358), .ZN(new_n1359));
  INV_X1    g1159(.A(KEYINPUT61), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1356), .A2(new_n1359), .A3(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1326), .A2(new_n1338), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1362), .A2(new_n1306), .A3(new_n1347), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT63), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1361), .B1(new_n1363), .B2(new_n1364), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1346), .A2(new_n1348), .A3(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT62), .ZN(new_n1367));
  AND3_X1   g1167(.A1(new_n1339), .A2(new_n1367), .A3(new_n1347), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1360), .B1(new_n1339), .B2(new_n1321), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1367), .B1(new_n1339), .B2(new_n1347), .ZN(new_n1370));
  NOR3_X1   g1170(.A1(new_n1368), .A2(new_n1369), .A3(new_n1370), .ZN(new_n1371));
  AND3_X1   g1171(.A1(new_n1356), .A2(KEYINPUT127), .A3(new_n1359), .ZN(new_n1372));
  AOI21_X1  g1172(.A(KEYINPUT127), .B1(new_n1356), .B2(new_n1359), .ZN(new_n1373));
  NOR2_X1   g1173(.A1(new_n1372), .A2(new_n1373), .ZN(new_n1374));
  INV_X1    g1174(.A(new_n1374), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1366), .B1(new_n1371), .B2(new_n1375), .ZN(G405));
  INV_X1    g1176(.A(new_n1299), .ZN(new_n1377));
  OAI21_X1  g1177(.A(new_n1326), .B1(new_n1271), .B2(new_n1377), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1378), .A2(new_n1347), .ZN(new_n1379));
  OR2_X1    g1179(.A1(new_n1378), .A2(new_n1347), .ZN(new_n1380));
  AND3_X1   g1180(.A1(new_n1374), .A2(new_n1379), .A3(new_n1380), .ZN(new_n1381));
  AOI21_X1  g1181(.A(new_n1374), .B1(new_n1379), .B2(new_n1380), .ZN(new_n1382));
  NOR2_X1   g1182(.A1(new_n1381), .A2(new_n1382), .ZN(G402));
endmodule


