//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n564, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT67), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT69), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n471), .B(G125), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n463), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n461), .B(new_n462), .C1(new_n473), .C2(new_n474), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n467), .A2(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n479), .A2(G137), .B1(G101), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n477), .A2(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n468), .A2(new_n469), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n463), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n460), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI22_X1  g062(.A1(G124), .A2(new_n485), .B1(new_n487), .B2(G136), .ZN(new_n488));
  INV_X1    g063(.A(new_n462), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI221_X1 g066(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n491), .C2(G112), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT4), .B1(new_n478), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n491), .A2(new_n483), .A3(new_n497), .A4(G138), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n502));
  AND2_X1   g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n503), .B1(new_n473), .B2(new_n474), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT71), .B1(new_n499), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  AOI211_X1 g083(.A(new_n508), .B(new_n505), .C1(new_n496), .C2(new_n498), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n507), .A2(new_n509), .ZN(G164));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT72), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n511), .A2(new_n515), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n514), .A2(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT74), .B(G89), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n511), .A2(new_n524), .B1(G63), .B2(G651), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT5), .B(G543), .Z(new_n526));
  OAI21_X1  g101(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n512), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n511), .A2(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT73), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n527), .B1(new_n532), .B2(G51), .ZN(G168));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n526), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G651), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n538), .B2(new_n518), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(new_n532), .B2(G52), .ZN(G171));
  AND2_X1   g115(.A1(new_n532), .A2(G43), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n517), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n544), .B2(new_n518), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n515), .B(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g130(.A1(G78), .A2(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OR3_X1    g133(.A1(new_n530), .A2(KEYINPUT9), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT9), .B1(new_n530), .B2(new_n558), .ZN(new_n560));
  INV_X1    g135(.A(new_n518), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n559), .A2(new_n560), .B1(G91), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n557), .A2(new_n562), .ZN(G299));
  NAND2_X1  g138(.A1(new_n532), .A2(G52), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n564), .B(new_n537), .C1(new_n538), .C2(new_n518), .ZN(G301));
  INV_X1    g140(.A(G168), .ZN(G286));
  INV_X1    g141(.A(G166), .ZN(G303));
  NAND2_X1  g142(.A1(new_n512), .A2(G49), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT76), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n515), .A2(G74), .ZN(new_n570));
  AOI22_X1  g145(.A1(G87), .A2(new_n561), .B1(new_n570), .B2(G651), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(new_n561), .A2(G86), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n512), .A2(G48), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n517), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G305));
  NAND2_X1  g154(.A1(G72), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G60), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n526), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(new_n561), .B2(G85), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n529), .A2(new_n531), .ZN(new_n584));
  INV_X1    g159(.A(G47), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(G290));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NOR2_X1   g162(.A1(G301), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n532), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G54), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n561), .A2(G92), .ZN(new_n592));
  XOR2_X1   g167(.A(KEYINPUT77), .B(KEYINPUT10), .Z(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT79), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n553), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n591), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT80), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n591), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n588), .B1(new_n605), .B2(new_n587), .ZN(G284));
  XNOR2_X1  g181(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  INV_X1    g183(.A(G299), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G297));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND3_X1  g188(.A1(new_n602), .A2(new_n612), .A3(new_n604), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n483), .A2(new_n480), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  INV_X1    g195(.A(G2100), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n485), .A2(G123), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n487), .A2(G135), .ZN(new_n625));
  OAI221_X1 g200(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n491), .C2(G111), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND3_X1  g203(.A1(new_n622), .A2(new_n623), .A3(new_n628), .ZN(G156));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2443), .B(G2446), .Z(new_n641));
  OAI21_X1  g216(.A(G14), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT82), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT17), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2084), .B(G2090), .ZN(new_n648));
  NOR3_X1   g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n645), .B2(new_n647), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n646), .B2(new_n647), .ZN(new_n651));
  INV_X1    g226(.A(new_n647), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n652), .A2(new_n648), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n645), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT18), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n649), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2096), .B(G2100), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1956), .B(G2474), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1961), .B(G1966), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n660), .A2(new_n663), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT20), .Z(new_n667));
  AOI211_X1 g242(.A(new_n665), .B(new_n667), .C1(new_n660), .C2(new_n664), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT84), .ZN(new_n669));
  XOR2_X1   g244(.A(G1981), .B(G1986), .Z(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT83), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n669), .B(new_n675), .ZN(G229));
  NOR2_X1   g251(.A1(G6), .A2(G16), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n578), .B2(G16), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT32), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G1981), .ZN(new_n680));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G23), .ZN(new_n682));
  INV_X1    g257(.A(G288), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT33), .B(G1976), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n684), .B(new_n685), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n681), .A2(G22), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G166), .B2(new_n681), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1971), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n680), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT34), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n485), .A2(G119), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n487), .A2(G131), .ZN(new_n695));
  OAI221_X1 g270(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n491), .C2(G107), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G25), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT35), .B(G1991), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT85), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT86), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n701), .A2(new_n703), .B1(new_n704), .B2(KEYINPUT36), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n703), .B2(new_n701), .ZN(new_n706));
  MUX2_X1   g281(.A(G24), .B(G290), .S(G16), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1986), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n692), .A2(new_n693), .A3(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n704), .A2(KEYINPUT36), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n681), .A2(G4), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n605), .B2(new_n681), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT87), .B(G1348), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n491), .A2(G103), .A3(G2104), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT25), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n487), .A2(G139), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n483), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n718), .B(new_n719), .C1(new_n491), .C2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(new_n699), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n699), .B2(G33), .ZN(new_n724));
  INV_X1    g299(.A(G2072), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT88), .ZN(new_n727));
  NOR2_X1   g302(.A1(G16), .A2(G21), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G168), .B2(G16), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT92), .B(G1966), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n724), .A2(new_n725), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NOR2_X1   g307(.A1(G16), .A2(G19), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n546), .B2(G16), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(G1341), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n727), .A2(new_n731), .A3(new_n732), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n480), .A2(G105), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT89), .ZN(new_n738));
  INV_X1    g313(.A(G141), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(new_n486), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT26), .Z(new_n742));
  INV_X1    g317(.A(G129), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n484), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT90), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G29), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT91), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n747), .B(new_n748), .C1(G29), .C2(G32), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n748), .B2(new_n747), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT27), .B(G1996), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n736), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n681), .A2(G20), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT95), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT23), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G299), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1956), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G27), .A2(G29), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G164), .B2(G29), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(G2078), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n761), .A2(G2078), .ZN(new_n763));
  NOR3_X1   g338(.A1(new_n759), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G171), .A2(new_n681), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G5), .B2(new_n681), .ZN(new_n766));
  INV_X1    g341(.A(G1961), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n699), .A2(G35), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G162), .B2(new_n699), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT29), .B(G2090), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n734), .A2(G1341), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n766), .A2(new_n767), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n768), .A2(new_n772), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT31), .B(G11), .ZN(new_n776));
  INV_X1    g351(.A(G28), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(KEYINPUT30), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n699), .B1(new_n779), .B2(G28), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n627), .A2(new_n699), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n776), .B1(new_n778), .B2(new_n780), .C1(new_n781), .C2(KEYINPUT93), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(KEYINPUT93), .B2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n699), .A2(G26), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT28), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n485), .A2(G128), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n487), .A2(G140), .ZN(new_n787));
  OAI221_X1 g362(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n491), .C2(G116), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n785), .B1(new_n789), .B2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2067), .ZN(new_n791));
  INV_X1    g366(.A(G2084), .ZN(new_n792));
  NAND2_X1  g367(.A1(G160), .A2(G29), .ZN(new_n793));
  INV_X1    g368(.A(G34), .ZN(new_n794));
  AOI21_X1  g369(.A(G29), .B1(new_n794), .B2(KEYINPUT24), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(KEYINPUT24), .B2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n783), .B(new_n791), .C1(new_n792), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n792), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT94), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n775), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  AND4_X1   g376(.A1(new_n716), .A2(new_n753), .A3(new_n764), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n712), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(G311));
  INV_X1    g379(.A(KEYINPUT96), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n803), .B(new_n805), .ZN(G150));
  INV_X1    g381(.A(KEYINPUT99), .ZN(new_n807));
  INV_X1    g382(.A(G860), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n605), .A2(G559), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(KEYINPUT38), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(KEYINPUT38), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n532), .A2(G55), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT97), .B(G93), .ZN(new_n815));
  OAI22_X1  g390(.A1(new_n814), .A2(new_n517), .B1(new_n518), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n546), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n817), .A2(new_n546), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n812), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n822), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n810), .A2(new_n824), .A3(new_n811), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n808), .B1(new_n826), .B2(KEYINPUT39), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n823), .A2(new_n825), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT98), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT98), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n826), .A2(new_n831), .A3(KEYINPUT39), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n827), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n818), .A2(G860), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT37), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n807), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n835), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n832), .A2(new_n830), .ZN(new_n838));
  OAI211_X1 g413(.A(KEYINPUT99), .B(new_n837), .C1(new_n838), .C2(new_n827), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n839), .ZN(G145));
  XNOR2_X1  g415(.A(G160), .B(new_n627), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G162), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT100), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n789), .B(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n505), .B1(new_n496), .B2(new_n498), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT101), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n499), .A2(new_n506), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n845), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n746), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n848), .A2(new_n852), .A3(new_n746), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n855), .A2(new_n722), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n722), .B1(new_n847), .B2(new_n745), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n745), .B2(new_n847), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n697), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AOI22_X1  g436(.A1(G130), .A2(new_n485), .B1(new_n487), .B2(G142), .ZN(new_n862));
  OAI221_X1 g437(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n491), .C2(G118), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n619), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n697), .B1(new_n857), .B2(new_n859), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n861), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n857), .A2(new_n859), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n698), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n865), .B1(new_n870), .B2(new_n860), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n843), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n866), .B1(new_n861), .B2(new_n867), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n870), .A2(new_n865), .A3(new_n860), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n842), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g453(.A(G166), .B(new_n578), .ZN(new_n879));
  XNOR2_X1  g454(.A(G288), .B(G290), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(new_n881), .B2(new_n880), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n881), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n884), .A2(new_n879), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT42), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n601), .A2(G299), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n591), .A2(new_n609), .A3(new_n600), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT41), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n889), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n614), .A2(new_n824), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n822), .A2(new_n602), .A3(new_n612), .A4(new_n604), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT102), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n897), .A3(new_n890), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n898), .A2(new_n902), .A3(new_n894), .A4(new_n891), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n900), .A2(KEYINPUT104), .A3(new_n901), .A4(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n901), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n902), .B1(new_n895), .B2(new_n898), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n887), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n908), .A2(new_n887), .ZN(new_n910));
  OAI21_X1  g485(.A(G868), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n818), .A2(new_n587), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(G331));
  NAND2_X1  g488(.A1(G331), .A2(KEYINPUT105), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(G295));
  NAND2_X1  g492(.A1(G301), .A2(G286), .ZN(new_n918));
  NAND2_X1  g493(.A1(G171), .A2(G168), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n822), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n918), .A2(new_n919), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(new_n820), .A3(new_n821), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n824), .A2(new_n922), .A3(KEYINPUT106), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n921), .A2(new_n923), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n822), .A2(KEYINPUT107), .A3(new_n920), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n892), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n895), .A2(new_n927), .B1(new_n931), .B2(KEYINPUT108), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n931), .A2(KEYINPUT108), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n886), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n873), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n886), .B1(new_n932), .B2(new_n933), .ZN(new_n936));
  OR3_X1    g511(.A1(new_n935), .A2(KEYINPUT43), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n892), .B1(new_n925), .B2(new_n926), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n891), .A2(new_n929), .A3(new_n894), .A4(new_n930), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n939), .B2(new_n940), .ZN(new_n943));
  OAI22_X1  g518(.A1(new_n941), .A2(new_n943), .B1(new_n883), .B2(new_n885), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n944), .A2(new_n934), .A3(new_n873), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n937), .B(KEYINPUT44), .C1(new_n938), .C2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n935), .B2(new_n936), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n944), .A2(new_n934), .A3(new_n938), .A4(new_n873), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI211_X1 g527(.A(KEYINPUT110), .B(KEYINPUT44), .C1(new_n948), .C2(new_n949), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n946), .B1(new_n952), .B2(new_n953), .ZN(G397));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n507), .B2(new_n509), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT50), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n477), .A2(G40), .A3(new_n481), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n849), .A2(new_n955), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(KEYINPUT50), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n959), .A2(new_n960), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n849), .A2(KEYINPUT45), .A3(new_n955), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n961), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n968), .B2(new_n956), .ZN(new_n969));
  OAI22_X1  g544(.A1(new_n965), .A2(G2090), .B1(G1971), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G8), .ZN(new_n971));
  NOR2_X1   g546(.A1(G166), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n972), .B1(new_n975), .B2(KEYINPUT55), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n970), .A2(G8), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n477), .A2(G40), .A3(new_n481), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n962), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(new_n971), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1976), .ZN(new_n983));
  NOR2_X1   g558(.A1(G288), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT52), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(G1981), .B1(new_n575), .B2(new_n577), .ZN(new_n986));
  INV_X1    g561(.A(new_n577), .ZN(new_n987));
  INV_X1    g562(.A(G1981), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n987), .A2(new_n988), .A3(new_n573), .A4(new_n574), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(KEYINPUT49), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT49), .B1(new_n986), .B2(new_n989), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(KEYINPUT113), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n993));
  AOI211_X1 g568(.A(new_n993), .B(KEYINPUT49), .C1(new_n986), .C2(new_n989), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n990), .B(new_n981), .C1(new_n992), .C2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT52), .B1(G288), .B2(new_n983), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n981), .B(new_n996), .C1(new_n983), .C2(G288), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n985), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n985), .A2(new_n995), .A3(KEYINPUT114), .A4(new_n997), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n978), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n995), .A2(new_n983), .A3(new_n683), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n989), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1004), .A2(KEYINPUT115), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n982), .B1(new_n1004), .B2(KEYINPUT115), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n965), .A2(new_n767), .ZN(new_n1008));
  INV_X1    g583(.A(G2078), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n846), .A2(G1384), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n979), .B1(new_n1010), .B2(KEYINPUT45), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n849), .A2(new_n508), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n846), .A2(KEYINPUT71), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1384), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1009), .B(new_n1011), .C1(new_n1014), .C2(KEYINPUT45), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT122), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT122), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1015), .A2(new_n1019), .A3(new_n1016), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1008), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT125), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n968), .B1(new_n846), .B2(G1384), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n961), .B(new_n1023), .C1(new_n956), .C2(new_n968), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1009), .A2(KEYINPUT53), .ZN(new_n1025));
  OR2_X1    g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1021), .A2(new_n1022), .A3(G301), .A4(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1008), .A2(new_n1018), .A3(new_n1026), .A4(new_n1020), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT125), .B1(new_n1028), .B2(G171), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n961), .A2(new_n1023), .A3(KEYINPUT123), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1025), .B1(new_n1010), .B2(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT123), .B1(new_n961), .B2(new_n1023), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT124), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1034), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT124), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1036), .A2(new_n1037), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1008), .A2(new_n1018), .A3(new_n1039), .A4(new_n1020), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1030), .B1(new_n1040), .B2(G171), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1027), .A2(new_n1029), .A3(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT58), .B(G1341), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n980), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1996), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n969), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT59), .B1(new_n1046), .B2(new_n819), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n956), .A2(new_n968), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1011), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1049), .A2(G1996), .B1(new_n980), .B2(new_n1043), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(new_n546), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n979), .B1(new_n962), .B2(KEYINPUT50), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1055), .B(new_n955), .C1(new_n507), .C2(new_n509), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n758), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n557), .A2(new_n562), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n557), .B2(new_n562), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT56), .B(G2072), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1011), .B(new_n1063), .C1(new_n1014), .C2(KEYINPUT45), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1058), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT61), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1058), .A2(new_n1064), .A3(new_n1062), .A4(KEYINPUT118), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1348), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n965), .A2(new_n1071), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n962), .A2(new_n979), .A3(G2067), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1072), .A2(KEYINPUT60), .A3(new_n601), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1058), .A2(new_n1064), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1062), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(KEYINPUT61), .A3(new_n1065), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1053), .A2(new_n1070), .A3(new_n1075), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT60), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n963), .B1(new_n957), .B2(new_n958), .ZN(new_n1082));
  AOI21_X1  g657(.A(G1348), .B1(new_n1082), .B2(new_n960), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1081), .B1(new_n1083), .B2(new_n1073), .ZN(new_n1084));
  INV_X1    g659(.A(new_n601), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n956), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT111), .B1(new_n956), .B2(KEYINPUT50), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n963), .ZN(new_n1088));
  OAI211_X1 g663(.A(KEYINPUT60), .B(new_n1074), .C1(new_n1088), .C2(G1348), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1084), .A2(new_n1085), .A3(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1080), .A2(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1078), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1085), .B1(new_n1083), .B2(new_n1073), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(KEYINPUT119), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1096), .B(new_n1085), .C1(new_n1083), .C2(new_n1073), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1092), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1042), .B1(new_n1091), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1028), .A2(G171), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n767), .A2(new_n965), .B1(new_n1017), .B2(KEYINPUT122), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1101), .A2(G301), .A3(new_n1020), .A4(new_n1039), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1971), .B1(new_n1048), .B2(new_n1011), .ZN(new_n1107));
  INV_X1    g682(.A(G2090), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1054), .A2(new_n1056), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1106), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(KEYINPUT116), .B(new_n1109), .C1(new_n969), .C2(G1971), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(new_n1112), .A3(G8), .ZN(new_n1113));
  INV_X1    g688(.A(new_n977), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n998), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1115), .A2(new_n978), .ZN(new_n1116));
  NOR2_X1   g691(.A1(G168), .A2(new_n971), .ZN(new_n1117));
  INV_X1    g692(.A(G1966), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1024), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n965), .B2(G2084), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1117), .B1(new_n1120), .B2(G8), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1117), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT51), .B1(new_n1122), .B2(KEYINPUT120), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(G8), .B(new_n1123), .C1(new_n1120), .C2(G286), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1120), .A2(new_n1117), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1105), .A2(new_n1116), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1007), .B1(new_n1099), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT63), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1120), .A2(G8), .A3(G168), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n970), .A2(G8), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n1114), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1132), .A2(new_n978), .A3(new_n1133), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT117), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1115), .A2(new_n1133), .A3(new_n1138), .A4(new_n978), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1139), .A2(new_n1131), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1115), .A2(new_n1133), .A3(new_n978), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT117), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1137), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT126), .B1(new_n1130), .B2(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1145), .A2(new_n1092), .B1(new_n1090), .B2(new_n1080), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1115), .A2(new_n978), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1121), .A2(new_n1124), .B1(new_n1120), .B2(new_n1117), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1147), .B1(new_n1148), .B2(new_n1126), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1146), .A2(new_n1105), .A3(new_n1149), .A4(new_n1042), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1141), .A2(KEYINPUT117), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1139), .A2(new_n1131), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1136), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1150), .A2(new_n1151), .A3(new_n1154), .A4(new_n1007), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1128), .A2(KEYINPUT62), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1128), .A2(KEYINPUT62), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1147), .A2(new_n1100), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1144), .A2(new_n1155), .A3(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1023), .A2(new_n979), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n746), .A2(new_n1045), .ZN(new_n1162));
  XOR2_X1   g737(.A(new_n789), .B(G2067), .Z(new_n1163));
  OAI21_X1  g738(.A(G1996), .B1(new_n740), .B2(new_n744), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n698), .A2(new_n703), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n698), .A2(new_n703), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(G290), .B(G1986), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1161), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1160), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1169), .A2(new_n1161), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1161), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1174), .A2(G1986), .A3(G290), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT127), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT48), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1176), .A2(KEYINPUT48), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1173), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1161), .A2(new_n1045), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT46), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1163), .A2(new_n745), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1181), .B1(new_n1174), .B2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT47), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n1165), .A2(new_n1168), .B1(G2067), .B2(new_n789), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n1161), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1179), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1172), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g764(.A(G319), .ZN(new_n1191));
  NOR4_X1   g765(.A1(G229), .A2(new_n1191), .A3(G227), .A4(G401), .ZN(new_n1192));
  NAND3_X1  g766(.A1(new_n877), .A2(new_n950), .A3(new_n1192), .ZN(G225));
  INV_X1    g767(.A(G225), .ZN(G308));
endmodule


