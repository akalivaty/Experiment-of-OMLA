

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798;

  NOR2_X1 U375 ( .A1(n740), .A2(G953), .ZN(n742) );
  NAND2_X1 U376 ( .A1(n355), .A2(n354), .ZN(n353) );
  INV_X1 U377 ( .A(n698), .ZN(n354) );
  NOR2_X1 U378 ( .A1(n405), .A2(n580), .ZN(n644) );
  INV_X1 U379 ( .A(n497), .ZN(n420) );
  NAND2_X2 U380 ( .A1(n504), .A2(G214), .ZN(n705) );
  XNOR2_X2 U381 ( .A(n357), .B(n414), .ZN(n700) );
  XNOR2_X2 U382 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X2 U383 ( .A(n688), .B(n691), .ZN(n692) );
  NAND2_X2 U384 ( .A1(n611), .A2(n460), .ZN(n371) );
  NAND2_X1 U385 ( .A1(n703), .A2(n353), .ZN(n738) );
  INV_X1 U386 ( .A(n699), .ZN(n355) );
  NOR2_X1 U387 ( .A1(n661), .A2(n590), .ZN(n453) );
  NOR2_X1 U388 ( .A1(G237), .A2(G953), .ZN(n483) );
  XNOR2_X1 U389 ( .A(G107), .B(G104), .ZN(n500) );
  BUF_X1 U390 ( .A(G116), .Z(n386) );
  BUF_X1 U391 ( .A(G146), .Z(n751) );
  XOR2_X1 U392 ( .A(n686), .B(KEYINPUT59), .Z(n356) );
  AND2_X2 U393 ( .A1(n362), .A2(n361), .ZN(n360) );
  XNOR2_X2 U394 ( .A(n772), .B(n416), .ZN(n687) );
  XNOR2_X2 U395 ( .A(n445), .B(G472), .ZN(n722) );
  XNOR2_X2 U396 ( .A(n668), .B(n667), .ZN(n670) );
  XNOR2_X1 U397 ( .A(n377), .B(n356), .ZN(n376) );
  INV_X1 U398 ( .A(KEYINPUT15), .ZN(n503) );
  NAND2_X1 U399 ( .A1(n376), .A2(n375), .ZN(n374) );
  NAND2_X1 U400 ( .A1(n400), .A2(G475), .ZN(n377) );
  XNOR2_X1 U401 ( .A(n632), .B(KEYINPUT109), .ZN(n361) );
  NOR2_X1 U402 ( .A1(n369), .A2(n367), .ZN(n366) );
  AND2_X1 U403 ( .A1(n629), .A2(n757), .ZN(n393) );
  XNOR2_X1 U404 ( .A(n446), .B(KEYINPUT39), .ZN(n662) );
  XNOR2_X1 U405 ( .A(n413), .B(n412), .ZN(n750) );
  NAND2_X1 U406 ( .A1(n382), .A2(n440), .ZN(n716) );
  NOR2_X1 U407 ( .A1(n591), .A2(n494), .ZN(n654) );
  XNOR2_X1 U408 ( .A(n600), .B(KEYINPUT38), .ZN(n655) );
  XNOR2_X1 U409 ( .A(n546), .B(n545), .ZN(n582) );
  INV_X1 U410 ( .A(n771), .ZN(n375) );
  NAND2_X1 U411 ( .A1(G953), .A2(G902), .ZN(n564) );
  XNOR2_X2 U412 ( .A(n786), .B(n558), .ZN(n389) );
  NAND2_X1 U413 ( .A1(n360), .A2(n358), .ZN(n357) );
  NAND2_X1 U414 ( .A1(n415), .A2(n359), .ZN(n358) );
  NAND2_X1 U415 ( .A1(n384), .A2(n619), .ZN(n359) );
  NAND2_X1 U416 ( .A1(n404), .A2(n620), .ZN(n362) );
  NAND2_X1 U417 ( .A1(n363), .A2(KEYINPUT35), .ZN(n370) );
  NAND2_X1 U418 ( .A1(n364), .A2(n457), .ZN(n363) );
  AND2_X2 U419 ( .A1(n371), .A2(n372), .ZN(n364) );
  NAND2_X1 U420 ( .A1(n370), .A2(n365), .ZN(n678) );
  NAND2_X1 U421 ( .A1(n366), .A2(n457), .ZN(n365) );
  NAND2_X1 U422 ( .A1(n371), .A2(n368), .ZN(n367) );
  INV_X1 U423 ( .A(KEYINPUT35), .ZN(n368) );
  INV_X1 U424 ( .A(n372), .ZN(n369) );
  AND2_X2 U425 ( .A1(n458), .A2(n615), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n374), .B(n373), .ZN(G60) );
  INV_X1 U427 ( .A(KEYINPUT60), .ZN(n373) );
  NOR2_X1 U428 ( .A1(n678), .A2(n616), .ZN(n617) );
  NAND2_X1 U429 ( .A1(n648), .A2(n410), .ZN(n649) );
  XNOR2_X1 U430 ( .A(n750), .B(n411), .ZN(n410) );
  INV_X1 U431 ( .A(KEYINPUT47), .ZN(n411) );
  NAND2_X1 U432 ( .A1(n582), .A2(KEYINPUT69), .ZN(n435) );
  INV_X1 U433 ( .A(n634), .ZN(n415) );
  AND2_X1 U434 ( .A1(n424), .A2(n385), .ZN(n422) );
  NAND2_X1 U435 ( .A1(n436), .A2(n429), .ZN(n423) );
  NAND2_X1 U436 ( .A1(n438), .A2(n437), .ZN(n436) );
  INV_X1 U437 ( .A(G469), .ZN(n438) );
  XNOR2_X1 U438 ( .A(n549), .B(n548), .ZN(n719) );
  XNOR2_X1 U439 ( .A(n462), .B(n657), .ZN(n461) );
  XNOR2_X1 U440 ( .A(G101), .B(KEYINPUT93), .ZN(n501) );
  INV_X1 U441 ( .A(G110), .ZN(n499) );
  XNOR2_X1 U442 ( .A(n523), .B(n409), .ZN(n535) );
  INV_X1 U443 ( .A(KEYINPUT8), .ZN(n409) );
  XNOR2_X1 U444 ( .A(KEYINPUT70), .B(KEYINPUT4), .ZN(n488) );
  XNOR2_X1 U445 ( .A(KEYINPUT80), .B(KEYINPUT18), .ZN(n466) );
  XNOR2_X1 U446 ( .A(KEYINPUT17), .B(KEYINPUT81), .ZN(n467) );
  XNOR2_X1 U447 ( .A(n387), .B(n495), .ZN(n421) );
  AND2_X1 U448 ( .A1(n776), .A2(G224), .ZN(n387) );
  NAND2_X1 U449 ( .A1(G237), .A2(G234), .ZN(n471) );
  NAND2_X1 U450 ( .A1(n671), .A2(n437), .ZN(n546) );
  XNOR2_X1 U451 ( .A(KEYINPUT71), .B(G137), .ZN(n552) );
  NAND2_X1 U452 ( .A1(n535), .A2(G221), .ZN(n408) );
  XNOR2_X1 U453 ( .A(G128), .B(KEYINPUT94), .ZN(n536) );
  XNOR2_X1 U454 ( .A(G104), .B(G122), .ZN(n508) );
  XOR2_X1 U455 ( .A(KEYINPUT12), .B(G143), .Z(n509) );
  XNOR2_X1 U456 ( .A(n515), .B(n512), .ZN(n455) );
  XNOR2_X1 U457 ( .A(n506), .B(KEYINPUT10), .ZN(n407) );
  INV_X1 U458 ( .A(G140), .ZN(n506) );
  XNOR2_X1 U459 ( .A(n469), .B(n468), .ZN(n734) );
  XNOR2_X1 U460 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n468) );
  NOR2_X1 U461 ( .A1(n709), .A2(n708), .ZN(n469) );
  NAND2_X1 U462 ( .A1(n654), .A2(n447), .ZN(n446) );
  NOR2_X1 U463 ( .A1(n655), .A2(n448), .ZN(n447) );
  XNOR2_X1 U464 ( .A(n521), .B(n520), .ZN(n628) );
  NAND2_X1 U465 ( .A1(n686), .A2(n437), .ZN(n521) );
  NAND2_X1 U466 ( .A1(n390), .A2(KEYINPUT34), .ZN(n457) );
  XNOR2_X1 U467 ( .A(n541), .B(KEYINPUT20), .ZN(n547) );
  NAND2_X1 U468 ( .A1(n540), .A2(G234), .ZN(n541) );
  XNOR2_X1 U469 ( .A(n453), .B(n452), .ZN(n710) );
  INV_X1 U470 ( .A(KEYINPUT107), .ZN(n452) );
  NAND2_X1 U471 ( .A1(G902), .A2(G469), .ZN(n439) );
  INV_X1 U472 ( .A(G237), .ZN(n491) );
  XOR2_X1 U473 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n482) );
  INV_X1 U474 ( .A(KEYINPUT45), .ZN(n414) );
  NAND2_X1 U475 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U476 ( .A1(n378), .A2(KEYINPUT1), .ZN(n425) );
  XNOR2_X1 U477 ( .A(n571), .B(KEYINPUT0), .ZN(n572) );
  NAND2_X1 U478 ( .A1(n718), .A2(n592), .ZN(n405) );
  BUF_X1 U479 ( .A(n700), .Z(n775) );
  XNOR2_X1 U480 ( .A(n467), .B(n466), .ZN(n465) );
  XNOR2_X1 U481 ( .A(n756), .B(KEYINPUT106), .ZN(n661) );
  NAND2_X1 U482 ( .A1(n442), .A2(n380), .ZN(n440) );
  NAND2_X1 U483 ( .A1(n575), .A2(KEYINPUT69), .ZN(n443) );
  INV_X2 U484 ( .A(G953), .ZN(n776) );
  XNOR2_X1 U485 ( .A(n444), .B(n406), .ZN(n671) );
  XNOR2_X1 U486 ( .A(n379), .B(n539), .ZN(n444) );
  XNOR2_X1 U487 ( .A(n408), .B(n785), .ZN(n406) );
  XNOR2_X1 U488 ( .A(n511), .B(n454), .ZN(n686) );
  XNOR2_X1 U489 ( .A(n455), .B(n517), .ZN(n454) );
  AND2_X1 U490 ( .A1(n674), .A2(G953), .ZN(n771) );
  AND2_X1 U491 ( .A1(n601), .A2(n464), .ZN(n664) );
  XNOR2_X1 U492 ( .A(n653), .B(n463), .ZN(n797) );
  INV_X1 U493 ( .A(KEYINPUT42), .ZN(n463) );
  INV_X1 U494 ( .A(KEYINPUT83), .ZN(n412) );
  NOR2_X1 U495 ( .A1(n652), .A2(n647), .ZN(n413) );
  AND2_X1 U496 ( .A1(n628), .A2(n627), .ZN(n756) );
  AND2_X1 U497 ( .A1(n586), .A2(n596), .ZN(n602) );
  INV_X1 U498 ( .A(G122), .ZN(n677) );
  NOR2_X1 U499 ( .A1(n760), .A2(n436), .ZN(n378) );
  XOR2_X1 U500 ( .A(n381), .B(n536), .Z(n379) );
  AND2_X1 U501 ( .A1(n550), .A2(n441), .ZN(n380) );
  XOR2_X1 U502 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n381) );
  AND2_X1 U503 ( .A1(n435), .A2(n443), .ZN(n382) );
  AND2_X1 U504 ( .A1(n504), .A2(G210), .ZN(n383) );
  OR2_X1 U505 ( .A1(n678), .A2(KEYINPUT44), .ZN(n384) );
  AND2_X1 U506 ( .A1(n423), .A2(n439), .ZN(n385) );
  INV_X1 U507 ( .A(G902), .ZN(n437) );
  BUF_X1 U508 ( .A(n582), .Z(n718) );
  AND2_X1 U509 ( .A1(n623), .A2(n580), .ZN(n744) );
  INV_X1 U510 ( .A(KEYINPUT1), .ZN(n429) );
  INV_X1 U511 ( .A(n600), .ZN(n464) );
  XOR2_X1 U512 ( .A(KEYINPUT5), .B(n386), .Z(n477) );
  BUF_X1 U513 ( .A(n715), .Z(n433) );
  NAND2_X1 U514 ( .A1(n715), .A2(n716), .ZN(n403) );
  NAND2_X1 U515 ( .A1(n426), .A2(n425), .ZN(n715) );
  NAND2_X1 U516 ( .A1(n716), .A2(n579), .ZN(n448) );
  BUF_X1 U517 ( .A(n522), .Z(n388) );
  XNOR2_X1 U518 ( .A(n786), .B(n558), .ZN(n760) );
  XNOR2_X1 U519 ( .A(n407), .B(n507), .ZN(n785) );
  XNOR2_X1 U520 ( .A(n751), .B(G137), .ZN(n481) );
  XNOR2_X1 U521 ( .A(n450), .B(n608), .ZN(n390) );
  BUF_X1 U522 ( .A(n631), .Z(n391) );
  AND2_X1 U523 ( .A1(n623), .A2(n394), .ZN(n392) );
  NOR2_X1 U524 ( .A1(n392), .A2(n393), .ZN(n630) );
  AND2_X1 U525 ( .A1(n580), .A2(n629), .ZN(n394) );
  XNOR2_X1 U526 ( .A(n395), .B(n396), .ZN(n605) );
  NOR2_X2 U527 ( .A1(n585), .A2(n584), .ZN(n395) );
  XOR2_X1 U528 ( .A(KEYINPUT66), .B(KEYINPUT32), .Z(n396) );
  NAND2_X1 U529 ( .A1(n459), .A2(KEYINPUT34), .ZN(n458) );
  NAND2_X1 U530 ( .A1(n586), .A2(n397), .ZN(n603) );
  AND2_X1 U531 ( .A1(n596), .A2(n580), .ZN(n397) );
  NAND2_X1 U532 ( .A1(n434), .A2(n718), .ZN(n606) );
  AND2_X1 U533 ( .A1(n610), .A2(n612), .ZN(n460) );
  XNOR2_X1 U534 ( .A(n578), .B(n577), .ZN(n398) );
  NOR2_X1 U535 ( .A1(n670), .A2(n669), .ZN(n399) );
  NOR2_X2 U536 ( .A1(n670), .A2(n669), .ZN(n400) );
  XNOR2_X1 U537 ( .A(n578), .B(n577), .ZN(n586) );
  NOR2_X2 U538 ( .A1(n670), .A2(n669), .ZN(n767) );
  BUF_X1 U539 ( .A(n553), .Z(n401) );
  BUF_X1 U540 ( .A(n678), .Z(n402) );
  XNOR2_X1 U541 ( .A(n450), .B(n449), .ZN(n611) );
  XNOR2_X1 U542 ( .A(n624), .B(KEYINPUT110), .ZN(n451) );
  XNOR2_X2 U543 ( .A(n403), .B(KEYINPUT75), .ZN(n624) );
  NAND2_X1 U544 ( .A1(n617), .A2(n618), .ZN(n404) );
  NOR2_X1 U545 ( .A1(n593), .A2(n405), .ZN(n594) );
  XNOR2_X1 U546 ( .A(n417), .B(n496), .ZN(n416) );
  XNOR2_X1 U547 ( .A(n421), .B(n465), .ZN(n417) );
  XNOR2_X2 U548 ( .A(n418), .B(n557), .ZN(n772) );
  XNOR2_X2 U549 ( .A(n502), .B(n501), .ZN(n557) );
  XNOR2_X2 U550 ( .A(n419), .B(n498), .ZN(n418) );
  XNOR2_X2 U551 ( .A(n522), .B(n420), .ZN(n419) );
  XNOR2_X2 U552 ( .A(n479), .B(n478), .ZN(n498) );
  NAND2_X1 U553 ( .A1(n431), .A2(n439), .ZN(n430) );
  NAND2_X1 U554 ( .A1(n422), .A2(n431), .ZN(n428) );
  NAND2_X1 U555 ( .A1(n760), .A2(n429), .ZN(n424) );
  NAND2_X1 U556 ( .A1(n428), .A2(n427), .ZN(n426) );
  NAND2_X1 U557 ( .A1(n430), .A2(n429), .ZN(n427) );
  OR2_X1 U558 ( .A1(n378), .A2(n430), .ZN(n579) );
  NAND2_X1 U559 ( .A1(n389), .A2(G469), .ZN(n431) );
  XNOR2_X1 U560 ( .A(n603), .B(KEYINPUT67), .ZN(n434) );
  NAND2_X1 U561 ( .A1(n630), .A2(n631), .ZN(n632) );
  INV_X2 U562 ( .A(G116), .ZN(n432) );
  XNOR2_X2 U563 ( .A(n432), .B(G122), .ZN(n522) );
  NAND2_X2 U564 ( .A1(n609), .A2(n576), .ZN(n578) );
  NAND2_X1 U565 ( .A1(n776), .A2(G234), .ZN(n523) );
  INV_X1 U566 ( .A(KEYINPUT69), .ZN(n441) );
  INV_X1 U567 ( .A(n582), .ZN(n442) );
  INV_X1 U568 ( .A(n722), .ZN(n580) );
  NAND2_X1 U569 ( .A1(n722), .A2(n705), .ZN(n492) );
  NAND2_X1 U570 ( .A1(n680), .A2(n437), .ZN(n445) );
  INV_X1 U571 ( .A(n608), .ZN(n449) );
  NAND2_X1 U572 ( .A1(n451), .A2(n607), .ZN(n450) );
  BUF_X2 U573 ( .A(n609), .Z(n610) );
  XNOR2_X2 U574 ( .A(n456), .B(G143), .ZN(n526) );
  XNOR2_X2 U575 ( .A(G128), .B(KEYINPUT84), .ZN(n456) );
  INV_X1 U576 ( .A(n610), .ZN(n459) );
  NAND2_X1 U577 ( .A1(n658), .A2(n461), .ZN(n660) );
  NAND2_X1 U578 ( .A1(n797), .A2(n798), .ZN(n462) );
  NAND2_X1 U579 ( .A1(n399), .A2(G217), .ZN(n673) );
  XNOR2_X2 U580 ( .A(n526), .B(n488), .ZN(n496) );
  INV_X1 U581 ( .A(n671), .ZN(n672) );
  NOR2_X1 U582 ( .A1(n713), .A2(n390), .ZN(n470) );
  INV_X1 U583 ( .A(KEYINPUT44), .ZN(n616) );
  INV_X1 U584 ( .A(KEYINPUT102), .ZN(n513) );
  XNOR2_X1 U585 ( .A(n514), .B(n513), .ZN(n515) );
  BUF_X1 U586 ( .A(n389), .Z(n763) );
  XNOR2_X1 U587 ( .A(KEYINPUT40), .B(n656), .ZN(n798) );
  XNOR2_X1 U588 ( .A(n471), .B(KEYINPUT14), .ZN(n731) );
  NOR2_X1 U589 ( .A1(G900), .A2(n564), .ZN(n472) );
  NAND2_X1 U590 ( .A1(n731), .A2(n472), .ZN(n473) );
  XNOR2_X1 U591 ( .A(n473), .B(KEYINPUT111), .ZN(n476) );
  INV_X1 U592 ( .A(n731), .ZN(n474) );
  NAND2_X1 U593 ( .A1(n776), .A2(G952), .ZN(n568) );
  NOR2_X1 U594 ( .A1(n474), .A2(n568), .ZN(n475) );
  NOR2_X1 U595 ( .A1(n476), .A2(n475), .ZN(n591) );
  XNOR2_X1 U596 ( .A(KEYINPUT30), .B(KEYINPUT113), .ZN(n493) );
  XNOR2_X1 U597 ( .A(n477), .B(G101), .ZN(n480) );
  XNOR2_X2 U598 ( .A(G119), .B(G113), .ZN(n479) );
  XNOR2_X2 U599 ( .A(KEYINPUT72), .B(KEYINPUT3), .ZN(n478) );
  XNOR2_X1 U600 ( .A(n480), .B(n498), .ZN(n487) );
  XNOR2_X1 U601 ( .A(n482), .B(n481), .ZN(n485) );
  XNOR2_X1 U602 ( .A(n483), .B(KEYINPUT78), .ZN(n516) );
  NAND2_X1 U603 ( .A1(n516), .A2(G210), .ZN(n484) );
  XNOR2_X1 U604 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U605 ( .A(n487), .B(n486), .ZN(n490) );
  XNOR2_X1 U606 ( .A(G134), .B(G131), .ZN(n489) );
  XNOR2_X2 U607 ( .A(n496), .B(n489), .ZN(n553) );
  XNOR2_X1 U608 ( .A(n401), .B(n490), .ZN(n680) );
  NAND2_X1 U609 ( .A1(n437), .A2(n491), .ZN(n504) );
  XOR2_X1 U610 ( .A(n493), .B(n492), .Z(n494) );
  XNOR2_X2 U611 ( .A(G125), .B(G146), .ZN(n507) );
  INV_X1 U612 ( .A(n507), .ZN(n495) );
  XNOR2_X2 U613 ( .A(KEYINPUT74), .B(KEYINPUT16), .ZN(n497) );
  XNOR2_X1 U614 ( .A(n500), .B(n499), .ZN(n502) );
  XNOR2_X2 U615 ( .A(n503), .B(G902), .ZN(n667) );
  INV_X1 U616 ( .A(n667), .ZN(n540) );
  NAND2_X1 U617 ( .A1(n687), .A2(n540), .ZN(n505) );
  XNOR2_X2 U618 ( .A(n505), .B(n383), .ZN(n561) );
  BUF_X1 U619 ( .A(n561), .Z(n600) );
  NAND2_X1 U620 ( .A1(n654), .A2(n600), .ZN(n534) );
  XOR2_X1 U621 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n512) );
  XNOR2_X1 U622 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U623 ( .A(n785), .B(n510), .ZN(n511) );
  XNOR2_X1 U624 ( .A(G113), .B(G131), .ZN(n514) );
  AND2_X1 U625 ( .A1(n516), .A2(G214), .ZN(n517) );
  XOR2_X1 U626 ( .A(KEYINPUT13), .B(KEYINPUT104), .Z(n519) );
  XNOR2_X1 U627 ( .A(KEYINPUT103), .B(G475), .ZN(n518) );
  XNOR2_X1 U628 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U629 ( .A(n388), .B(KEYINPUT9), .Z(n525) );
  NAND2_X1 U630 ( .A1(G217), .A2(n535), .ZN(n524) );
  XNOR2_X1 U631 ( .A(n525), .B(n524), .ZN(n532) );
  INV_X1 U632 ( .A(n526), .ZN(n530) );
  XOR2_X1 U633 ( .A(KEYINPUT7), .B(KEYINPUT105), .Z(n528) );
  XNOR2_X1 U634 ( .A(G107), .B(G134), .ZN(n527) );
  XNOR2_X1 U635 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U636 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U637 ( .A(n532), .B(n531), .ZN(n769) );
  NAND2_X1 U638 ( .A1(n769), .A2(n437), .ZN(n533) );
  XNOR2_X1 U639 ( .A(n533), .B(G478), .ZN(n627) );
  INV_X1 U640 ( .A(n627), .ZN(n574) );
  OR2_X1 U641 ( .A1(n628), .A2(n574), .ZN(n614) );
  NOR2_X1 U642 ( .A1(n534), .A2(n614), .ZN(n551) );
  INV_X1 U643 ( .A(G119), .ZN(n537) );
  XNOR2_X1 U644 ( .A(n537), .B(G110), .ZN(n538) );
  XNOR2_X1 U645 ( .A(n552), .B(n538), .ZN(n539) );
  XOR2_X1 U646 ( .A(KEYINPUT96), .B(KEYINPUT25), .Z(n543) );
  NAND2_X1 U647 ( .A1(n547), .A2(G217), .ZN(n542) );
  XNOR2_X1 U648 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U649 ( .A(n544), .B(KEYINPUT95), .ZN(n545) );
  NAND2_X1 U650 ( .A1(n547), .A2(G221), .ZN(n549) );
  XOR2_X1 U651 ( .A(KEYINPUT97), .B(KEYINPUT21), .Z(n548) );
  XNOR2_X1 U652 ( .A(n719), .B(KEYINPUT98), .ZN(n575) );
  INV_X1 U653 ( .A(n575), .ZN(n550) );
  AND2_X1 U654 ( .A1(n551), .A2(n716), .ZN(n559) );
  XNOR2_X2 U655 ( .A(n553), .B(n552), .ZN(n786) );
  XNOR2_X1 U656 ( .A(n751), .B(G140), .ZN(n555) );
  NAND2_X1 U657 ( .A1(n776), .A2(G227), .ZN(n554) );
  XNOR2_X1 U658 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U659 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U660 ( .A1(n559), .A2(n579), .ZN(n641) );
  XOR2_X1 U661 ( .A(G143), .B(KEYINPUT117), .Z(n560) );
  XNOR2_X1 U662 ( .A(n641), .B(n560), .ZN(G45) );
  NAND2_X1 U663 ( .A1(n561), .A2(n705), .ZN(n562) );
  XNOR2_X1 U664 ( .A(n562), .B(KEYINPUT90), .ZN(n635) );
  XNOR2_X1 U665 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n563) );
  XNOR2_X1 U666 ( .A(n635), .B(n563), .ZN(n646) );
  INV_X1 U667 ( .A(G898), .ZN(n566) );
  INV_X1 U668 ( .A(n564), .ZN(n565) );
  NAND2_X1 U669 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U670 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U671 ( .A1(n731), .A2(n569), .ZN(n570) );
  OR2_X2 U672 ( .A1(n646), .A2(n570), .ZN(n573) );
  INV_X1 U673 ( .A(KEYINPUT68), .ZN(n571) );
  XNOR2_X2 U674 ( .A(n573), .B(n572), .ZN(n609) );
  NAND2_X1 U675 ( .A1(n628), .A2(n574), .ZN(n708) );
  NOR2_X1 U676 ( .A1(n708), .A2(n575), .ZN(n576) );
  INV_X1 U677 ( .A(KEYINPUT22), .ZN(n577) );
  INV_X1 U678 ( .A(n398), .ZN(n585) );
  INV_X1 U679 ( .A(n433), .ZN(n596) );
  INV_X1 U680 ( .A(KEYINPUT6), .ZN(n581) );
  XNOR2_X1 U681 ( .A(n580), .B(n581), .ZN(n587) );
  NAND2_X1 U682 ( .A1(n587), .A2(n718), .ZN(n583) );
  OR2_X1 U683 ( .A1(n596), .A2(n583), .ZN(n584) );
  XNOR2_X1 U684 ( .A(n605), .B(G119), .ZN(G21) );
  INV_X1 U685 ( .A(n587), .ZN(n607) );
  NOR2_X1 U686 ( .A1(n607), .A2(n718), .ZN(n588) );
  NAND2_X1 U687 ( .A1(n602), .A2(n588), .ZN(n589) );
  XNOR2_X1 U688 ( .A(n589), .B(KEYINPUT108), .ZN(n631) );
  XNOR2_X1 U689 ( .A(n391), .B(G101), .ZN(G3) );
  NOR2_X1 U690 ( .A1(n628), .A2(n627), .ZN(n590) );
  INV_X1 U691 ( .A(n590), .ZN(n593) );
  NOR2_X1 U692 ( .A1(n719), .A2(n591), .ZN(n592) );
  NAND2_X1 U693 ( .A1(n594), .A2(n607), .ZN(n637) );
  INV_X1 U694 ( .A(n705), .ZN(n595) );
  NOR2_X1 U695 ( .A1(n637), .A2(n595), .ZN(n597) );
  NAND2_X1 U696 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U697 ( .A(n598), .B(KEYINPUT112), .ZN(n599) );
  XNOR2_X1 U698 ( .A(n599), .B(KEYINPUT43), .ZN(n601) );
  XOR2_X1 U699 ( .A(n664), .B(G140), .Z(G42) );
  XNOR2_X1 U700 ( .A(G110), .B(KEYINPUT116), .ZN(n604) );
  XNOR2_X1 U701 ( .A(n606), .B(n604), .ZN(G12) );
  NAND2_X1 U702 ( .A1(n606), .A2(n605), .ZN(n633) );
  INV_X1 U703 ( .A(KEYINPUT65), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n633), .A2(n619), .ZN(n618) );
  XNOR2_X1 U705 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n608) );
  INV_X1 U706 ( .A(KEYINPUT34), .ZN(n612) );
  INV_X1 U707 ( .A(KEYINPUT82), .ZN(n613) );
  XNOR2_X1 U708 ( .A(n614), .B(n613), .ZN(n615) );
  NAND2_X1 U709 ( .A1(n619), .A2(n616), .ZN(n620) );
  AND2_X1 U710 ( .A1(n716), .A2(n579), .ZN(n621) );
  NAND2_X1 U711 ( .A1(n610), .A2(n621), .ZN(n622) );
  XNOR2_X1 U712 ( .A(n622), .B(KEYINPUT99), .ZN(n623) );
  AND2_X1 U713 ( .A1(n624), .A2(n722), .ZN(n714) );
  NAND2_X1 U714 ( .A1(n610), .A2(n714), .ZN(n626) );
  XNOR2_X1 U715 ( .A(KEYINPUT100), .B(KEYINPUT31), .ZN(n625) );
  XNOR2_X1 U716 ( .A(n626), .B(n625), .ZN(n757) );
  INV_X1 U717 ( .A(n710), .ZN(n629) );
  BUF_X1 U718 ( .A(n633), .Z(n634) );
  BUF_X1 U719 ( .A(n635), .Z(n636) );
  NOR2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U721 ( .A(n638), .B(KEYINPUT36), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n639), .A2(n433), .ZN(n640) );
  XNOR2_X1 U723 ( .A(n640), .B(KEYINPUT115), .ZN(n795) );
  NAND2_X1 U724 ( .A1(n710), .A2(KEYINPUT47), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U726 ( .A(n643), .B(KEYINPUT85), .ZN(n650) );
  XNOR2_X1 U727 ( .A(KEYINPUT28), .B(n644), .ZN(n645) );
  NAND2_X1 U728 ( .A1(n645), .A2(n579), .ZN(n652) );
  BUF_X1 U729 ( .A(n646), .Z(n647) );
  NAND2_X1 U730 ( .A1(n750), .A2(n710), .ZN(n648) );
  NAND2_X1 U731 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U732 ( .A1(n795), .A2(n651), .ZN(n658) );
  XOR2_X1 U733 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n657) );
  INV_X1 U734 ( .A(n655), .ZN(n706) );
  NOR2_X1 U735 ( .A1(n734), .A2(n652), .ZN(n653) );
  NAND2_X1 U736 ( .A1(n590), .A2(n662), .ZN(n656) );
  XNOR2_X1 U737 ( .A(KEYINPUT48), .B(KEYINPUT89), .ZN(n659) );
  XNOR2_X1 U738 ( .A(n660), .B(n659), .ZN(n666) );
  NAND2_X1 U739 ( .A1(n662), .A2(n661), .ZN(n759) );
  INV_X1 U740 ( .A(n759), .ZN(n663) );
  NOR2_X1 U741 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U742 ( .A1(n666), .A2(n665), .ZN(n787) );
  NOR2_X2 U743 ( .A1(n700), .A2(n787), .ZN(n696) );
  NOR2_X2 U744 ( .A1(n696), .A2(KEYINPUT88), .ZN(n668) );
  XNOR2_X1 U745 ( .A(n696), .B(KEYINPUT2), .ZN(n669) );
  XNOR2_X1 U746 ( .A(n673), .B(n672), .ZN(n675) );
  INV_X1 U747 ( .A(G952), .ZN(n674) );
  NOR2_X2 U748 ( .A1(n675), .A2(n771), .ZN(n676) );
  XNOR2_X1 U749 ( .A(n676), .B(KEYINPUT124), .ZN(G66) );
  XNOR2_X1 U750 ( .A(n402), .B(n677), .ZN(G24) );
  NAND2_X1 U751 ( .A1(n767), .A2(G472), .ZN(n682) );
  XNOR2_X1 U752 ( .A(KEYINPUT91), .B(KEYINPUT62), .ZN(n679) );
  XNOR2_X1 U753 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X2 U754 ( .A1(n683), .A2(n771), .ZN(n685) );
  XOR2_X1 U755 ( .A(KEYINPUT92), .B(KEYINPUT63), .Z(n684) );
  XNOR2_X1 U756 ( .A(n685), .B(n684), .ZN(G57) );
  NAND2_X1 U757 ( .A1(n767), .A2(G210), .ZN(n693) );
  BUF_X1 U758 ( .A(n687), .Z(n688) );
  XOR2_X1 U759 ( .A(KEYINPUT86), .B(KEYINPUT55), .Z(n690) );
  XNOR2_X1 U760 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n689) );
  XOR2_X1 U761 ( .A(n690), .B(n689), .Z(n691) );
  XNOR2_X1 U762 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X2 U763 ( .A1(n694), .A2(n771), .ZN(n695) );
  XNOR2_X1 U764 ( .A(n695), .B(KEYINPUT56), .ZN(G51) );
  BUF_X1 U765 ( .A(n696), .Z(n697) );
  INV_X1 U766 ( .A(KEYINPUT2), .ZN(n701) );
  NOR2_X1 U767 ( .A1(n697), .A2(n701), .ZN(n699) );
  NOR2_X1 U768 ( .A1(n787), .A2(KEYINPUT2), .ZN(n698) );
  NAND2_X1 U769 ( .A1(n775), .A2(n701), .ZN(n702) );
  XOR2_X1 U770 ( .A(KEYINPUT87), .B(n702), .Z(n703) );
  NOR2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n712) );
  NOR2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U774 ( .A1(n712), .A2(n711), .ZN(n713) );
  INV_X1 U775 ( .A(n714), .ZN(n726) );
  OR2_X1 U776 ( .A1(n716), .A2(n433), .ZN(n717) );
  XNOR2_X1 U777 ( .A(n717), .B(KEYINPUT50), .ZN(n724) );
  NAND2_X1 U778 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U779 ( .A(KEYINPUT49), .B(n720), .ZN(n721) );
  NOR2_X1 U780 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U781 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U782 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U783 ( .A(KEYINPUT51), .B(n727), .ZN(n728) );
  NOR2_X1 U784 ( .A1(n734), .A2(n728), .ZN(n729) );
  NOR2_X1 U785 ( .A1(n470), .A2(n729), .ZN(n730) );
  XNOR2_X1 U786 ( .A(n730), .B(KEYINPUT52), .ZN(n733) );
  NAND2_X1 U787 ( .A1(n731), .A2(G952), .ZN(n732) );
  NOR2_X1 U788 ( .A1(n733), .A2(n732), .ZN(n736) );
  NOR2_X1 U789 ( .A1(n734), .A2(n390), .ZN(n735) );
  NOR2_X1 U790 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U791 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U792 ( .A(n739), .B(KEYINPUT120), .ZN(n740) );
  XOR2_X1 U793 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n741) );
  XNOR2_X1 U794 ( .A(n742), .B(n741), .ZN(G75) );
  NAND2_X1 U795 ( .A1(n744), .A2(n590), .ZN(n743) );
  XNOR2_X1 U796 ( .A(n743), .B(G104), .ZN(G6) );
  XOR2_X1 U797 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n746) );
  NAND2_X1 U798 ( .A1(n744), .A2(n756), .ZN(n745) );
  XNOR2_X1 U799 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U800 ( .A(G107), .B(n747), .ZN(G9) );
  XOR2_X1 U801 ( .A(G128), .B(KEYINPUT29), .Z(n749) );
  NAND2_X1 U802 ( .A1(n750), .A2(n756), .ZN(n748) );
  XNOR2_X1 U803 ( .A(n749), .B(n748), .ZN(G30) );
  NAND2_X1 U804 ( .A1(n750), .A2(n590), .ZN(n752) );
  XNOR2_X1 U805 ( .A(n752), .B(n751), .ZN(G48) );
  XOR2_X1 U806 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n754) );
  NAND2_X1 U807 ( .A1(n590), .A2(n757), .ZN(n753) );
  XNOR2_X1 U808 ( .A(n754), .B(n753), .ZN(n755) );
  XNOR2_X1 U809 ( .A(G113), .B(n755), .ZN(G15) );
  NAND2_X1 U810 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U811 ( .A(n758), .B(n386), .ZN(G18) );
  XNOR2_X1 U812 ( .A(G134), .B(n759), .ZN(G36) );
  NAND2_X1 U813 ( .A1(n400), .A2(G469), .ZN(n765) );
  XOR2_X1 U814 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n761) );
  XOR2_X1 U815 ( .A(n761), .B(KEYINPUT123), .Z(n762) );
  XNOR2_X1 U816 ( .A(n763), .B(n762), .ZN(n764) );
  XNOR2_X1 U817 ( .A(n765), .B(n764), .ZN(n766) );
  NOR2_X1 U818 ( .A1(n771), .A2(n766), .ZN(G54) );
  NAND2_X1 U819 ( .A1(n400), .A2(G478), .ZN(n768) );
  XOR2_X1 U820 ( .A(n769), .B(n768), .Z(n770) );
  NOR2_X1 U821 ( .A1(n771), .A2(n770), .ZN(G63) );
  XNOR2_X1 U822 ( .A(n772), .B(KEYINPUT126), .ZN(n774) );
  NOR2_X1 U823 ( .A1(G898), .A2(n776), .ZN(n773) );
  NOR2_X1 U824 ( .A1(n774), .A2(n773), .ZN(n784) );
  INV_X1 U825 ( .A(n775), .ZN(n777) );
  NAND2_X1 U826 ( .A1(n777), .A2(n776), .ZN(n782) );
  XOR2_X1 U827 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n779) );
  NAND2_X1 U828 ( .A1(G224), .A2(G953), .ZN(n778) );
  XNOR2_X1 U829 ( .A(n779), .B(n778), .ZN(n780) );
  NAND2_X1 U830 ( .A1(n780), .A2(G898), .ZN(n781) );
  NAND2_X1 U831 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U832 ( .A(n784), .B(n783), .ZN(G69) );
  XNOR2_X1 U833 ( .A(n786), .B(n785), .ZN(n790) );
  XNOR2_X1 U834 ( .A(n787), .B(n790), .ZN(n788) );
  NOR2_X1 U835 ( .A1(G953), .A2(n788), .ZN(n789) );
  XNOR2_X1 U836 ( .A(n789), .B(KEYINPUT127), .ZN(n794) );
  XOR2_X1 U837 ( .A(G227), .B(n790), .Z(n791) );
  NAND2_X1 U838 ( .A1(n791), .A2(G900), .ZN(n792) );
  NAND2_X1 U839 ( .A1(n792), .A2(G953), .ZN(n793) );
  NAND2_X1 U840 ( .A1(n794), .A2(n793), .ZN(G72) );
  XNOR2_X1 U841 ( .A(G125), .B(n795), .ZN(n796) );
  XNOR2_X1 U842 ( .A(n796), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U843 ( .A(G137), .B(n797), .ZN(G39) );
  XNOR2_X1 U844 ( .A(G131), .B(n798), .ZN(G33) );
endmodule

