//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT70), .B(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G234), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT24), .B(G110), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G110), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n199), .B1(new_n193), .B2(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(new_n194), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n198), .B1(new_n202), .B2(KEYINPUT72), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT72), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n200), .A2(new_n201), .A3(new_n204), .A4(new_n194), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n197), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G125), .B(G140), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT73), .A3(KEYINPUT16), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G125), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G140), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT16), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT73), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n211), .B2(KEYINPUT16), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n208), .B(new_n209), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n214), .B(new_n216), .C1(KEYINPUT16), .C2(new_n211), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n209), .B1(new_n220), .B2(new_n208), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n206), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n208), .B1(new_n215), .B2(new_n217), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n195), .A2(new_n196), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(G110), .B2(new_n202), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n207), .A2(new_n209), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT74), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT74), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n222), .A2(new_n231), .A3(new_n228), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT22), .B(G137), .ZN(new_n233));
  INV_X1    g047(.A(G953), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(G221), .A3(G234), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n233), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(KEYINPUT75), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n230), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n222), .A2(new_n228), .A3(new_n236), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n188), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT76), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n190), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(new_n241), .A3(KEYINPUT25), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n244), .A2(KEYINPUT77), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT77), .B1(new_n244), .B2(new_n245), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n238), .A2(new_n239), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n189), .A2(G902), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT32), .ZN(new_n254));
  XOR2_X1   g068(.A(G116), .B(G119), .Z(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT2), .B(G113), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT64), .B(G143), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(G146), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n209), .A2(G143), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n265));
  INV_X1    g079(.A(G134), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(G137), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(G137), .ZN(new_n268));
  INV_X1    g082(.A(G137), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT11), .A3(G134), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G131), .ZN(new_n272));
  INV_X1    g086(.A(G131), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n267), .A2(new_n270), .A3(new_n273), .A4(new_n268), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n209), .A2(G143), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n277), .B1(new_n261), .B2(G146), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n258), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n264), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n269), .A2(G134), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n266), .A2(G137), .ZN(new_n282));
  OAI21_X1  g096(.A(G131), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n191), .B1(new_n276), .B2(KEYINPUT1), .ZN(new_n285));
  INV_X1    g099(.A(G143), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT64), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT64), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G143), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n209), .ZN(new_n291));
  INV_X1    g105(.A(new_n263), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n285), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n287), .A2(new_n289), .A3(G146), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n294), .A2(new_n276), .A3(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n284), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT30), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n280), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n280), .B2(new_n297), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n257), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT65), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT65), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n303), .B(new_n257), .C1(new_n299), .C2(new_n300), .ZN(new_n304));
  INV_X1    g118(.A(new_n257), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n280), .A2(new_n297), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G237), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(new_n234), .A3(G210), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT27), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G101), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT66), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n280), .A2(new_n297), .A3(new_n305), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT66), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(new_n311), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n302), .A2(new_n304), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT31), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n305), .B1(new_n280), .B2(new_n297), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT28), .B1(new_n306), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT68), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n306), .B2(KEYINPUT28), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n314), .A2(KEYINPUT68), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n317), .A2(new_n318), .B1(new_n312), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n302), .A2(new_n304), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n313), .A2(new_n316), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT67), .A3(KEYINPUT31), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT67), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n317), .B2(new_n318), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n326), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(G472), .A2(G902), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n254), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n254), .A3(new_n334), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n327), .A2(new_n314), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n312), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n320), .A2(new_n322), .A3(new_n311), .A4(new_n324), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n188), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n280), .A2(new_n297), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n257), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n323), .B1(new_n347), .B2(new_n314), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n314), .A2(KEYINPUT68), .A3(new_n323), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT68), .B1(new_n314), .B2(new_n323), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n351), .A2(KEYINPUT69), .A3(KEYINPUT29), .A4(new_n311), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT69), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(new_n341), .B2(new_n342), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n345), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n344), .B1(new_n355), .B2(KEYINPUT71), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT71), .ZN(new_n357));
  AOI211_X1 g171(.A(new_n357), .B(new_n345), .C1(new_n352), .C2(new_n354), .ZN(new_n358));
  OAI21_X1  g172(.A(G472), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n253), .B1(new_n338), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT5), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n193), .A3(G116), .ZN(new_n362));
  OAI211_X1 g176(.A(G113), .B(new_n362), .C1(new_n255), .C2(new_n361), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n255), .B2(new_n256), .ZN(new_n364));
  INV_X1    g178(.A(G104), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G107), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n365), .A2(G107), .ZN(new_n368));
  OAI21_X1  g182(.A(G101), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT3), .B1(new_n365), .B2(G107), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n371));
  INV_X1    g185(.A(G107), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(G104), .ZN(new_n373));
  INV_X1    g187(.A(G101), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n370), .A2(new_n373), .A3(new_n374), .A4(new_n366), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n364), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n370), .A2(new_n373), .A3(new_n366), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G101), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT79), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n375), .A2(KEYINPUT4), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n382), .A3(G101), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT80), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n382), .B1(new_n378), .B2(G101), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n375), .A2(KEYINPUT4), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT80), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(new_n383), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n379), .A2(KEYINPUT4), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n305), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n377), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(G110), .B(G122), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT84), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n394), .B2(new_n395), .ZN(new_n398));
  AND4_X1   g212(.A1(new_n389), .A2(new_n380), .A3(new_n383), .A4(new_n381), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n389), .B1(new_n388), .B2(new_n383), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n393), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n377), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n404));
  INV_X1    g218(.A(new_n395), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n396), .A2(new_n398), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n392), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n257), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n385), .B2(new_n390), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n397), .B(new_n405), .C1(new_n410), .C2(new_n377), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT85), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT85), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n403), .A2(new_n413), .A3(new_n397), .A4(new_n405), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n264), .A2(new_n279), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(new_n212), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n293), .A2(new_n296), .A3(G125), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n234), .A2(G224), .ZN(new_n420));
  XOR2_X1   g234(.A(new_n420), .B(KEYINPUT86), .Z(new_n421));
  XNOR2_X1  g235(.A(new_n419), .B(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n407), .A2(new_n415), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n407), .A2(new_n415), .A3(KEYINPUT87), .A4(new_n422), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G210), .B1(G237), .B2(G902), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n419), .A2(KEYINPUT7), .A3(new_n420), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT88), .B(KEYINPUT8), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n395), .B(new_n430), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n364), .A2(new_n376), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n431), .B1(new_n432), .B2(new_n377), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n420), .A2(KEYINPUT7), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n417), .B2(new_n418), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n429), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n403), .A2(new_n405), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(G902), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n427), .A2(new_n428), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT89), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n428), .B1(new_n427), .B2(new_n439), .ZN(new_n443));
  INV_X1    g257(.A(new_n428), .ZN(new_n444));
  INV_X1    g258(.A(new_n439), .ZN(new_n445));
  AOI211_X1 g259(.A(new_n444), .B(new_n445), .C1(new_n425), .C2(new_n426), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n442), .B1(new_n447), .B2(new_n441), .ZN(new_n448));
  OAI21_X1  g262(.A(G214), .B1(G237), .B2(G902), .ZN(new_n449));
  INV_X1    g263(.A(G469), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n416), .B(new_n408), .C1(new_n399), .C2(new_n400), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n294), .A2(new_n276), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT1), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n290), .B2(new_n209), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n452), .B1(new_n454), .B2(new_n191), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n278), .A2(new_n295), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n376), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT10), .ZN(new_n460));
  INV_X1    g274(.A(new_n285), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n461), .B1(new_n262), .B2(new_n263), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n462), .B2(new_n456), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n459), .A2(new_n460), .B1(new_n463), .B2(new_n458), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n275), .B(KEYINPUT81), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n451), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G110), .B(G140), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT78), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n234), .A2(G227), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n468), .B(new_n469), .Z(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT82), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n458), .A2(new_n293), .A3(new_n296), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n376), .B1(new_n455), .B2(new_n456), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n472), .B(new_n275), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT83), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT12), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(KEYINPUT83), .B(new_n275), .C1(new_n474), .C2(new_n473), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n477), .B1(new_n475), .B2(new_n476), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n471), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n416), .A2(new_n408), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n390), .B2(new_n385), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n463), .A2(new_n458), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(KEYINPUT10), .B2(new_n474), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n275), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n470), .B1(new_n489), .B2(new_n466), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n450), .B(new_n188), .C1(new_n484), .C2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n466), .B1(new_n480), .B2(new_n482), .ZN(new_n492));
  INV_X1    g306(.A(new_n470), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n471), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n489), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(G469), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G902), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n450), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n491), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT9), .B(G234), .ZN(new_n502));
  OAI21_X1  g316(.A(G221), .B1(new_n502), .B2(G902), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n211), .A2(new_n213), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G146), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n227), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n307), .A2(new_n234), .A3(G143), .A4(G214), .ZN(new_n508));
  NAND2_X1  g322(.A1(KEYINPUT18), .A2(G131), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n307), .A2(new_n234), .A3(G214), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n508), .B(new_n509), .C1(new_n290), .C2(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n508), .B1(new_n290), .B2(new_n510), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(KEYINPUT18), .A3(G131), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(G113), .B(G122), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(new_n365), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(G131), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n224), .B(new_n218), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n273), .B(new_n508), .C1(new_n290), .C2(new_n510), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(KEYINPUT17), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n515), .B(new_n517), .C1(new_n520), .C2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n517), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT19), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n505), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n207), .A2(KEYINPUT19), .ZN(new_n528));
  AOI21_X1  g342(.A(G146), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(G146), .B2(new_n223), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n530), .A2(new_n522), .B1(new_n514), .B2(new_n512), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n525), .B1(new_n531), .B2(KEYINPUT90), .ZN(new_n532));
  INV_X1    g346(.A(new_n529), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n522), .A2(new_n224), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n515), .A3(KEYINPUT90), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n524), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT20), .ZN(new_n538));
  NOR2_X1   g352(.A1(G475), .A2(G902), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n539), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(KEYINPUT91), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT91), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n543), .B(new_n524), .C1(new_n532), .C2(new_n536), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n541), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n540), .B1(new_n545), .B2(new_n538), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n515), .B1(new_n520), .B2(new_n523), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n525), .A2(KEYINPUT92), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n548), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n498), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G475), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n191), .A2(G143), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n261), .B2(G128), .ZN(new_n556));
  INV_X1    g370(.A(G122), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G116), .ZN(new_n558));
  INV_X1    g372(.A(G116), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(G122), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G107), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n560), .A3(new_n372), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n556), .A2(new_n266), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n287), .A2(new_n289), .A3(G128), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n554), .A2(KEYINPUT13), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n261), .A2(KEYINPUT13), .A3(G128), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n567), .A2(new_n568), .A3(KEYINPUT93), .ZN(new_n569));
  OAI21_X1  g383(.A(G134), .B1(new_n567), .B2(KEYINPUT93), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n564), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT14), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(new_n559), .A3(G122), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT94), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT94), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n575), .A2(new_n572), .A3(new_n559), .A4(G122), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n560), .A2(KEYINPUT14), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n574), .A2(new_n558), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G107), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n565), .A2(new_n266), .A3(new_n554), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n266), .B1(new_n565), .B2(new_n554), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n579), .B(new_n563), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n571), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n502), .A2(new_n187), .A3(G953), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n571), .A2(new_n582), .A3(new_n584), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n188), .ZN(new_n589));
  INV_X1    g403(.A(G478), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(KEYINPUT15), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n589), .A2(new_n591), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(G234), .A2(G237), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n595), .A2(G952), .A3(new_n234), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n345), .A2(G953), .A3(new_n595), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT21), .B(G898), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n504), .A2(new_n553), .A3(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n360), .A2(new_n448), .A3(new_n449), .A4(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  NAND2_X1  g418(.A1(new_n242), .A2(new_n243), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n245), .A3(new_n189), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT77), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n244), .A2(KEYINPUT77), .A3(new_n245), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n608), .A2(new_n609), .A3(new_n252), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n333), .A2(new_n188), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n611), .A2(G472), .B1(new_n334), .B2(new_n333), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n588), .A2(new_n590), .A3(new_n188), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n571), .A2(new_n582), .A3(new_n584), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n584), .B1(new_n571), .B2(new_n582), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT33), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n586), .A2(new_n617), .A3(new_n587), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n345), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n613), .B1(new_n619), .B2(new_n590), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT95), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT95), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n622), .B(new_n613), .C1(new_n619), .C2(new_n590), .ZN(new_n623));
  AOI221_X4 g437(.A(new_n599), .B1(new_n621), .B2(new_n623), .C1(new_n546), .C2(new_n552), .ZN(new_n624));
  INV_X1    g438(.A(new_n503), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n470), .B(new_n466), .C1(new_n480), .C2(new_n482), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n489), .A2(new_n466), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n493), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n345), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n499), .B1(new_n629), .B2(new_n450), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n625), .B1(new_n630), .B2(new_n497), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n610), .A2(new_n612), .A3(new_n624), .A4(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n449), .B1(new_n443), .B2(new_n446), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT34), .B(G104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  INV_X1    g450(.A(new_n612), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n637), .A2(new_n253), .A3(new_n504), .ZN(new_n638));
  INV_X1    g452(.A(new_n633), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n552), .B1(new_n592), .B2(new_n593), .ZN(new_n640));
  INV_X1    g454(.A(new_n544), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n534), .A2(new_n515), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT90), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n535), .A3(new_n525), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n543), .B1(new_n645), .B2(new_n524), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n539), .B1(new_n641), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT20), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n545), .A2(new_n538), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n599), .B(new_n640), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n638), .A2(new_n639), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  AND2_X1   g467(.A1(new_n230), .A2(new_n232), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n237), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n251), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n608), .A2(new_n609), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n637), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n448), .A2(new_n659), .A3(new_n449), .A4(new_n602), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  INV_X1    g476(.A(KEYINPUT98), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n504), .B1(new_n248), .B2(new_n657), .ZN(new_n664));
  INV_X1    g478(.A(new_n337), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n359), .B1(new_n665), .B2(new_n335), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n597), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n596), .B1(new_n669), .B2(KEYINPUT96), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(KEYINPUT96), .B2(new_n669), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT97), .Z(new_n672));
  AOI211_X1 g486(.A(new_n672), .B(new_n640), .C1(new_n648), .C2(new_n649), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n449), .B(new_n673), .C1(new_n443), .C2(new_n446), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n663), .B1(new_n667), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n608), .A2(new_n609), .A3(new_n657), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n631), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n338), .B2(new_n359), .ZN(new_n678));
  INV_X1    g492(.A(new_n674), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n679), .A3(KEYINPUT98), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  XNOR2_X1  g496(.A(new_n448), .B(KEYINPUT38), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n672), .B(KEYINPUT39), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n504), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT40), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n594), .B1(new_n546), .B2(new_n552), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n658), .A2(new_n449), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n312), .B1(new_n306), .B2(new_n319), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n329), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n498), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n336), .A2(new_n337), .B1(G472), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n683), .A2(new_n686), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n290), .ZN(G45));
  NAND2_X1  g509(.A1(new_n621), .A2(new_n623), .ZN(new_n696));
  INV_X1    g510(.A(new_n672), .ZN(new_n697));
  INV_X1    g511(.A(new_n540), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n647), .B2(KEYINPUT20), .ZN(new_n699));
  INV_X1    g513(.A(new_n552), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n696), .B(new_n697), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT99), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n553), .A2(KEYINPUT99), .A3(new_n696), .A4(new_n697), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n678), .A2(new_n639), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  NAND2_X1  g522(.A1(new_n481), .A2(new_n483), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n490), .B1(new_n709), .B2(new_n495), .ZN(new_n710));
  OAI21_X1  g524(.A(G469), .B1(new_n710), .B2(new_n345), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n711), .A2(new_n503), .A3(new_n491), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n360), .A2(new_n639), .A3(new_n624), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND4_X1  g529(.A1(new_n360), .A2(new_n639), .A3(new_n650), .A4(new_n712), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  OAI211_X1 g531(.A(new_n449), .B(new_n712), .C1(new_n443), .C2(new_n446), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n658), .A2(new_n553), .A3(new_n601), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n666), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT100), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n317), .A2(new_n318), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n325), .A2(new_n312), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n317), .A2(new_n318), .ZN(new_n729));
  OAI211_X1 g543(.A(KEYINPUT100), .B(new_n726), .C1(new_n317), .C2(new_n318), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n611), .A2(G472), .B1(new_n731), .B2(new_n334), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n610), .A3(new_n600), .A4(new_n712), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n449), .B(new_n687), .C1(new_n443), .C2(new_n446), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT101), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  AOI211_X1 g551(.A(new_n723), .B(new_n733), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n734), .B(new_n735), .ZN(new_n739));
  INV_X1    g553(.A(new_n733), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT102), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT103), .B(G122), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G24));
  NAND2_X1  g558(.A1(new_n611), .A2(G472), .ZN(new_n745));
  INV_X1    g559(.A(new_n728), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n730), .A2(new_n729), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n334), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n676), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n705), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n719), .A3(KEYINPUT104), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT104), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n732), .A2(new_n703), .A3(new_n704), .A4(new_n676), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n752), .B1(new_n753), .B2(new_n718), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  INV_X1    g570(.A(new_n449), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n427), .A2(new_n439), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n444), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n441), .A3(new_n440), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n446), .A2(KEYINPUT89), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n499), .B(KEYINPUT105), .Z(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n629), .B2(new_n450), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n625), .B1(new_n765), .B2(new_n497), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n762), .A2(new_n360), .A3(new_n706), .A4(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n768), .A2(KEYINPUT106), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g584(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n771));
  NAND2_X1  g585(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G131), .ZN(G33));
  NAND4_X1  g588(.A1(new_n762), .A2(new_n360), .A3(new_n673), .A4(new_n766), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  AND2_X1   g590(.A1(new_n494), .A2(new_n496), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(KEYINPUT45), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(KEYINPUT45), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(G469), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT46), .B1(new_n780), .B2(new_n763), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n781), .B1(new_n450), .B2(new_n629), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(KEYINPUT46), .A3(new_n763), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n503), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n684), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n553), .B1(new_n621), .B2(new_n623), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT43), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n637), .A3(new_n676), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(KEYINPUT44), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(KEYINPUT44), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n786), .A2(new_n791), .A3(new_n762), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  XNOR2_X1  g608(.A(new_n785), .B(KEYINPUT47), .ZN(new_n795));
  INV_X1    g609(.A(new_n762), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n706), .A2(new_n338), .A3(new_n359), .A4(new_n253), .ZN(new_n797));
  OR3_X1    g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  AND2_X1   g613(.A1(new_n711), .A2(new_n491), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(KEYINPUT49), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(KEYINPUT49), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n449), .A3(new_n503), .A4(new_n787), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n692), .A2(new_n610), .ZN(new_n805));
  OR4_X1    g619(.A1(new_n683), .A2(new_n802), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n594), .B(KEYINPUT107), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n552), .A3(new_n697), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n648), .B2(new_n649), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(new_n666), .A3(new_n664), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n491), .A2(new_n497), .A3(new_n763), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n503), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n705), .A2(new_n749), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n762), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n775), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n770), .B2(new_n772), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n713), .A2(new_n716), .A3(new_n721), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n739), .A2(new_n740), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n723), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n739), .A2(KEYINPUT102), .A3(new_n740), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT108), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n807), .A2(new_n553), .A3(new_n599), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n448), .A2(new_n822), .A3(new_n449), .A4(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n760), .A2(new_n449), .A3(new_n823), .A4(new_n761), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT108), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n824), .A2(new_n826), .A3(new_n638), .ZN(new_n827));
  INV_X1    g641(.A(new_n632), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n448), .A3(new_n449), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n603), .A2(new_n660), .A3(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n827), .A2(new_n830), .A3(KEYINPUT109), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT109), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n760), .A2(new_n602), .A3(new_n449), .A4(new_n761), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n666), .A2(new_n610), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n760), .A2(new_n449), .A3(new_n761), .ZN(new_n835));
  OAI22_X1  g649(.A1(new_n833), .A2(new_n834), .B1(new_n835), .B2(new_n632), .ZN(new_n836));
  INV_X1    g650(.A(new_n659), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n833), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n824), .A2(new_n826), .A3(new_n638), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n832), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n816), .B(new_n821), .C1(new_n831), .C2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n658), .A2(KEYINPUT110), .A3(new_n697), .A4(new_n766), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT110), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n608), .A2(new_n609), .A3(new_n657), .A4(new_n697), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n845), .B1(new_n846), .B2(new_n812), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n692), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n734), .A2(new_n735), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n734), .A2(new_n735), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n681), .A2(new_n755), .A3(new_n851), .A4(new_n707), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n852), .A2(KEYINPUT52), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(KEYINPUT111), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n667), .A2(new_n633), .A3(new_n705), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n675), .B2(new_n680), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT111), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n857), .A3(new_n755), .A4(new_n851), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT52), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n853), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n843), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n859), .A2(new_n860), .ZN(new_n865));
  INV_X1    g679(.A(new_n817), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n741), .B2(new_n738), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n839), .A2(new_n832), .A3(new_n840), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT109), .B1(new_n827), .B2(new_n830), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n854), .A2(new_n858), .A3(KEYINPUT52), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n865), .A2(new_n870), .A3(new_n816), .A4(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n864), .B1(new_n863), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT54), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n843), .A2(KEYINPUT53), .A3(new_n861), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n854), .A2(KEYINPUT52), .A3(new_n858), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT52), .B1(new_n854), .B2(new_n858), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n842), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n875), .B1(new_n878), .B2(KEYINPUT53), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n874), .B1(KEYINPUT54), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n795), .B1(new_n503), .B2(new_n801), .ZN(new_n881));
  INV_X1    g695(.A(new_n732), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n253), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n788), .A2(new_n596), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n881), .A2(new_n883), .A3(new_n762), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n883), .ZN(new_n887));
  INV_X1    g701(.A(new_n712), .ZN(new_n888));
  NOR4_X1   g702(.A1(new_n887), .A2(new_n683), .A3(new_n449), .A4(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT50), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n796), .A2(new_n888), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n610), .A2(new_n891), .A3(new_n596), .A4(new_n692), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n553), .A2(new_n696), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n885), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n749), .ZN(new_n896));
  AOI22_X1  g710(.A1(new_n892), .A2(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n886), .A2(new_n890), .A3(new_n897), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT51), .Z(new_n899));
  NAND2_X1  g713(.A1(new_n895), .A2(new_n360), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT48), .ZN(new_n901));
  OAI211_X1 g715(.A(G952), .B(new_n234), .C1(new_n887), .C2(new_n718), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n553), .A2(new_n696), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n903), .B2(new_n892), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT112), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n880), .A2(new_n899), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(G952), .A2(G953), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n806), .B1(new_n907), .B2(new_n908), .ZN(G75));
  INV_X1    g723(.A(new_n879), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n188), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT56), .B1(new_n911), .B2(new_n444), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n407), .A2(new_n415), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n422), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n912), .B(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n234), .A2(G952), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT113), .Z(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n916), .A2(new_n919), .ZN(G51));
  XNOR2_X1  g734(.A(new_n879), .B(KEYINPUT54), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n763), .B(KEYINPUT114), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT57), .Z(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n710), .B(KEYINPUT115), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OR3_X1    g740(.A1(new_n910), .A2(new_n188), .A3(new_n780), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n917), .B1(new_n926), .B2(new_n927), .ZN(G54));
  NAND3_X1  g742(.A1(new_n911), .A2(KEYINPUT58), .A3(G475), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n542), .A2(new_n544), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n929), .A2(new_n931), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n932), .A2(new_n933), .A3(new_n917), .ZN(G60));
  NAND2_X1  g748(.A1(new_n616), .A2(new_n618), .ZN(new_n935));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT59), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n880), .B2(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n935), .A2(new_n937), .ZN(new_n939));
  AOI211_X1 g753(.A(new_n919), .B(new_n938), .C1(new_n921), .C2(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT60), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n876), .A2(new_n877), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT53), .B1(new_n944), .B2(new_n843), .ZN(new_n945));
  NOR4_X1   g759(.A1(new_n842), .A2(new_n877), .A3(new_n863), .A4(new_n853), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n249), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n872), .A2(new_n863), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n942), .B1(new_n949), .B2(new_n875), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n656), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n948), .A2(new_n951), .A3(KEYINPUT61), .A4(new_n918), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n953));
  OAI211_X1 g767(.A(KEYINPUT116), .B(new_n918), .C1(new_n950), .C2(new_n250), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n951), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT116), .B1(new_n948), .B2(new_n918), .ZN(new_n956));
  OAI211_X1 g770(.A(KEYINPUT117), .B(new_n953), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT116), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n250), .B1(new_n879), .B2(new_n943), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n960), .B2(new_n919), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n954), .A3(new_n951), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT117), .B1(new_n962), .B2(new_n953), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n952), .B1(new_n958), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT118), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT118), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n966), .B(new_n952), .C1(new_n958), .C2(new_n963), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n967), .ZN(G66));
  INV_X1    g782(.A(G224), .ZN(new_n969));
  OAI21_X1  g783(.A(G953), .B1(new_n598), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n870), .B2(G953), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n913), .B1(G898), .B2(new_n234), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(G69));
  NAND2_X1  g787(.A1(G900), .A2(G953), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n798), .A2(new_n793), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n856), .A2(new_n755), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT121), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n786), .A2(new_n360), .A3(new_n739), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n978), .A2(new_n775), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n975), .A2(new_n773), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n974), .B1(new_n980), .B2(G953), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n299), .A2(new_n300), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT119), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT120), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n527), .A2(new_n528), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n984), .B(new_n985), .Z(new_n986));
  NAND2_X1  g800(.A1(new_n981), .A2(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n977), .A2(new_n694), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT122), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n988), .A2(new_n989), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n796), .A2(new_n834), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n807), .A2(new_n553), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n993), .B(new_n685), .C1(new_n903), .C2(new_n994), .ZN(new_n995));
  AND4_X1   g809(.A1(new_n975), .A2(new_n991), .A3(new_n992), .A4(new_n995), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n986), .A2(G953), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n987), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n234), .B1(G227), .B2(G900), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT123), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n998), .B(new_n1000), .ZN(G72));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT63), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT124), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n870), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1005), .B1(new_n980), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n339), .A2(new_n311), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n917), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT126), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT127), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n317), .B1(new_n340), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n339), .A2(KEYINPUT127), .A3(new_n312), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1003), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n873), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1011), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1004), .B1(new_n996), .B2(new_n870), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT125), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n339), .A2(new_n311), .ZN(new_n1020));
  OR3_X1    g834(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1019), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1017), .B1(new_n1021), .B2(new_n1022), .ZN(G57));
endmodule


