//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(G50), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G13), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n216));
  XNOR2_X1  g0016(.A(new_n215), .B(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n203), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n210), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  INV_X1    g0025(.A(G97), .ZN(new_n226));
  INV_X1    g0026(.A(G257), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AND2_X1   g0028(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(G238), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n202), .ZN(new_n232));
  AOI22_X1  g0032(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n233));
  INV_X1    g0033(.A(G226), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n233), .B1(new_n205), .B2(new_n234), .ZN(new_n235));
  NOR4_X1   g0035(.A1(new_n229), .A2(new_n230), .A3(new_n232), .A4(new_n235), .ZN(new_n236));
  OR2_X1    g0036(.A1(new_n236), .A2(new_n211), .ZN(new_n237));
  OAI211_X1 g0037(.A(new_n217), .B(new_n222), .C1(new_n237), .C2(KEYINPUT1), .ZN(new_n238));
  AOI21_X1  g0038(.A(new_n238), .B1(KEYINPUT1), .B2(new_n237), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G264), .B(G270), .Z(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G358));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n249), .B(new_n250), .Z(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  NOR2_X1   g0055(.A1(new_n212), .A2(G1), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT70), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n212), .A2(new_n210), .A3(G1), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT70), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT12), .B1(new_n262), .B2(G68), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT12), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n256), .A2(new_n264), .A3(G20), .A4(new_n202), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n260), .B1(new_n256), .B2(G20), .ZN(new_n266));
  NOR4_X1   g0066(.A1(new_n212), .A2(new_n210), .A3(KEYINPUT70), .A4(G1), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n220), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n202), .B1(new_n209), .B2(G20), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n263), .A2(new_n265), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n210), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G77), .ZN(new_n275));
  OAI22_X1  g0075(.A1(new_n274), .A2(new_n275), .B1(new_n210), .B2(G68), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT73), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n210), .A2(new_n278), .ZN(new_n279));
  OAI22_X1  g0079(.A1(new_n276), .A2(new_n277), .B1(new_n205), .B2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n276), .A2(new_n277), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n270), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT11), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(KEYINPUT11), .B(new_n270), .C1(new_n280), .C2(new_n281), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n273), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n278), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n241), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n291), .A2(G1698), .B1(G33), .B2(G97), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT72), .ZN(new_n293));
  AOI21_X1  g0093(.A(G1698), .B1(new_n289), .B2(new_n290), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(G226), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  AND2_X1   g0096(.A1(KEYINPUT3), .A2(G33), .ZN(new_n297));
  NOR2_X1   g0097(.A1(KEYINPUT3), .A2(G33), .ZN(new_n298));
  OAI211_X1 g0098(.A(G226), .B(new_n296), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n292), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT13), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT67), .B(G45), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(G41), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n209), .A2(G274), .ZN(new_n307));
  INV_X1    g0107(.A(G41), .ZN(new_n308));
  OAI211_X1 g0108(.A(G1), .B(G13), .C1(new_n278), .C2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G238), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n306), .A2(new_n307), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n303), .A2(new_n304), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n289), .A2(new_n290), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n317), .A2(new_n293), .A3(G226), .A4(new_n296), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n309), .B1(new_n319), .B2(new_n292), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT13), .B1(new_n320), .B2(new_n313), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n315), .A2(new_n321), .A3(G190), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n287), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n315), .B2(new_n321), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n304), .B1(new_n303), .B2(new_n314), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n320), .A2(KEYINPUT13), .A3(new_n313), .ZN(new_n328));
  OAI21_X1  g0128(.A(G169), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT14), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n315), .A2(new_n321), .A3(G179), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT14), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n332), .B(G169), .C1(new_n327), .C2(new_n328), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n326), .B1(new_n334), .B2(new_n286), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT74), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT8), .B(G58), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(new_n209), .B2(G20), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n259), .A2(new_n270), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n339), .A2(new_n340), .B1(new_n259), .B2(new_n338), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n270), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n297), .A2(new_n298), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT7), .B1(new_n344), .B2(new_n210), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n289), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n290), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(G68), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G58), .A2(G68), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT76), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(KEYINPUT76), .A2(G58), .A3(G68), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n203), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT77), .ZN(new_n354));
  INV_X1    g0154(.A(G159), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n354), .B1(new_n279), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(G20), .A2(G33), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(KEYINPUT77), .A3(G159), .ZN(new_n358));
  AOI22_X1  g0158(.A1(G20), .A2(new_n353), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT16), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n343), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n348), .A2(KEYINPUT75), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n353), .A2(G20), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n356), .A2(new_n358), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT16), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n289), .A2(new_n210), .A3(new_n290), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT7), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n202), .B1(new_n370), .B2(new_n346), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT75), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n363), .A2(new_n367), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n342), .B1(new_n362), .B2(new_n374), .ZN(new_n375));
  OR2_X1    g0175(.A1(G223), .A2(G1698), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n234), .A2(G1698), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n376), .B(new_n377), .C1(new_n297), .C2(new_n298), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G33), .A2(G87), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT78), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT78), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n378), .A2(new_n382), .A3(new_n379), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n302), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G190), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n309), .A2(G232), .A3(new_n310), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n306), .B2(new_n307), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n384), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n309), .B1(new_n380), .B2(KEYINPUT78), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n387), .B1(new_n390), .B2(new_n383), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n389), .B1(G200), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n375), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT17), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n375), .A2(KEYINPUT17), .A3(new_n392), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G179), .ZN(new_n399));
  AOI211_X1 g0199(.A(new_n399), .B(new_n387), .C1(new_n390), .C2(new_n383), .ZN(new_n400));
  INV_X1    g0200(.A(G169), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(new_n384), .B2(new_n388), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT18), .B1(new_n375), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT79), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n370), .A2(new_n346), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n372), .B1(new_n406), .B2(G68), .ZN(new_n407));
  AOI211_X1 g0207(.A(KEYINPUT75), .B(new_n202), .C1(new_n370), .C2(new_n346), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n407), .A2(new_n408), .A3(new_n366), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n364), .A2(new_n365), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n361), .B1(new_n371), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n270), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n341), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n391), .A2(G179), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n401), .B2(new_n391), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n404), .A2(new_n405), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n405), .B1(new_n404), .B2(new_n417), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n398), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G244), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n306), .A2(new_n307), .B1(new_n311), .B2(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n291), .A2(new_n296), .B1(new_n344), .B2(G107), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n317), .A2(G1698), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n423), .B1(new_n231), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n422), .B1(new_n425), .B2(new_n302), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(KEYINPUT71), .A3(new_n399), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT71), .B1(new_n426), .B2(new_n399), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n338), .A2(new_n279), .B1(new_n210), .B2(new_n275), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n431), .A2(KEYINPUT69), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n278), .A2(G20), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT15), .B(G87), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n431), .A2(KEYINPUT69), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n343), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n262), .A2(new_n343), .ZN(new_n438));
  OAI21_X1  g0238(.A(G77), .B1(new_n210), .B2(G1), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n438), .A2(new_n439), .B1(G77), .B2(new_n262), .ZN(new_n440));
  OAI22_X1  g0240(.A1(G169), .A2(new_n426), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n430), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G150), .ZN(new_n444));
  OAI22_X1  g0244(.A1(new_n338), .A2(new_n274), .B1(new_n444), .B2(new_n279), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n210), .B1(new_n204), .B2(new_n205), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n270), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n205), .B1(new_n209), .B2(G20), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n340), .A2(new_n448), .B1(new_n205), .B2(new_n259), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n294), .A2(G222), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n317), .A2(G223), .A3(G1698), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n452), .B(new_n453), .C1(new_n275), .C2(new_n317), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n302), .ZN(new_n455));
  INV_X1    g0255(.A(new_n307), .ZN(new_n456));
  INV_X1    g0256(.A(new_n305), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n308), .ZN(new_n458));
  INV_X1    g0258(.A(new_n311), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n456), .A2(new_n458), .B1(new_n459), .B2(G226), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n451), .B1(new_n461), .B2(new_n401), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n455), .A2(new_n399), .A3(new_n460), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT68), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT68), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n462), .A2(new_n466), .A3(new_n463), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n437), .A2(new_n440), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n426), .A2(G190), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n469), .B(new_n470), .C1(new_n324), .C2(new_n426), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n461), .A2(G200), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n451), .A2(KEYINPUT9), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT9), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n450), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n455), .A2(G190), .A3(new_n460), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n472), .A2(new_n473), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT10), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n450), .B(KEYINPUT9), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT10), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n479), .A2(new_n480), .A3(new_n476), .A4(new_n472), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n443), .A2(new_n468), .A3(new_n471), .A4(new_n482), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n337), .A2(new_n420), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n335), .A2(new_n336), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G116), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n268), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n487), .B1(new_n209), .B2(G33), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n343), .B(new_n489), .C1(new_n266), .C2(new_n267), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n269), .A2(new_n220), .B1(G20), .B2(new_n487), .ZN(new_n491));
  AOI21_X1  g0291(.A(G20), .B1(G33), .B2(G283), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(G33), .B2(new_n226), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT20), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT20), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n488), .B(new_n490), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G45), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(G1), .ZN(new_n498));
  AND2_X1   g0298(.A1(KEYINPUT5), .A2(G41), .ZN(new_n499));
  NOR2_X1   g0299(.A1(KEYINPUT5), .A2(G41), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(G270), .A3(new_n309), .ZN(new_n502));
  OR2_X1    g0302(.A1(KEYINPUT5), .A2(G41), .ZN(new_n503));
  NAND2_X1  g0303(.A1(KEYINPUT5), .A2(G41), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G274), .A3(new_n498), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(G264), .B(G1698), .C1(new_n297), .C2(new_n298), .ZN(new_n508));
  OAI211_X1 g0308(.A(G257), .B(new_n296), .C1(new_n297), .C2(new_n298), .ZN(new_n509));
  INV_X1    g0309(.A(G303), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(new_n317), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n302), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n496), .A2(new_n513), .A3(G169), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT21), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n513), .A2(G200), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n488), .A2(new_n490), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n495), .A2(new_n494), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n507), .A2(new_n512), .A3(G190), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n513), .A2(new_n399), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n496), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n496), .A2(new_n513), .A3(KEYINPUT21), .A4(G169), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n516), .A2(new_n522), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G283), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n278), .A2(new_n527), .B1(KEYINPUT82), .B2(KEYINPUT4), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G250), .A2(G1698), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n296), .A2(G244), .ZN(new_n530));
  NAND2_X1  g0330(.A1(KEYINPUT82), .A2(KEYINPUT4), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n528), .B1(new_n532), .B2(new_n317), .ZN(new_n533));
  OAI211_X1 g0333(.A(G244), .B(new_n296), .C1(new_n297), .C2(new_n298), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n531), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n309), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n501), .A2(new_n309), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n506), .B1(new_n537), .B2(new_n227), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n399), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n401), .B1(new_n536), .B2(new_n538), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n357), .A2(G77), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT80), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n542), .B(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n406), .B2(G107), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT81), .ZN(new_n546));
  INV_X1    g0346(.A(G107), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT6), .A4(G97), .ZN(new_n548));
  NAND2_X1  g0348(.A1(KEYINPUT6), .A2(G97), .ZN(new_n549));
  OAI21_X1  g0349(.A(KEYINPUT81), .B1(new_n549), .B2(G107), .ZN(new_n550));
  AND2_X1   g0350(.A1(G97), .A2(G107), .ZN(new_n551));
  NOR2_X1   g0351(.A1(G97), .A2(G107), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n548), .B(new_n550), .C1(new_n553), .C2(KEYINPUT6), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G20), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n343), .B1(new_n545), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n259), .A2(new_n226), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n340), .B1(G1), .B2(new_n278), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n557), .B1(new_n558), .B2(new_n226), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n540), .B(new_n541), .C1(new_n556), .C2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n528), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n421), .A2(G1698), .ZN(new_n562));
  INV_X1    g0362(.A(new_n531), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n562), .A2(new_n563), .B1(G250), .B2(G1698), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n561), .B1(new_n564), .B2(new_n344), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n563), .B1(new_n294), .B2(G244), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n302), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n302), .B1(new_n505), .B2(new_n498), .ZN(new_n568));
  INV_X1    g0368(.A(new_n501), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n568), .A2(G257), .B1(new_n569), .B2(G274), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n385), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n324), .B1(new_n536), .B2(new_n538), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(G107), .B1(new_n345), .B2(new_n347), .ZN(new_n574));
  INV_X1    g0374(.A(new_n544), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n575), .A3(new_n555), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n559), .B1(new_n576), .B2(new_n270), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT19), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n433), .A2(new_n579), .A3(G97), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G97), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n552), .A2(new_n224), .B1(new_n581), .B2(new_n210), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n580), .B1(new_n582), .B2(new_n579), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n317), .A2(KEYINPUT83), .A3(new_n210), .A4(G68), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n210), .B(G68), .C1(new_n297), .C2(new_n298), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT83), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n583), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n270), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n268), .A2(new_n434), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n558), .C2(new_n434), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n312), .A2(new_n296), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n421), .A2(G1698), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n592), .B(new_n593), .C1(new_n297), .C2(new_n298), .ZN(new_n594));
  NAND2_X1  g0394(.A1(G33), .A2(G116), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n309), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(G250), .B1(new_n497), .B2(G1), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n302), .A2(new_n597), .B1(new_n497), .B2(new_n307), .ZN(new_n598));
  NOR3_X1   g0398(.A1(new_n596), .A2(G179), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n597), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(new_n309), .B1(new_n456), .B2(G45), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n594), .A2(new_n595), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(new_n309), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n599), .B1(new_n401), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n591), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n588), .A2(new_n270), .B1(new_n268), .B2(new_n434), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n596), .A2(new_n598), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G190), .ZN(new_n608));
  INV_X1    g0408(.A(new_n558), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G87), .ZN(new_n610));
  OAI21_X1  g0410(.A(G200), .B1(new_n596), .B2(new_n598), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n606), .A2(new_n608), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n560), .A2(new_n578), .A3(new_n605), .A4(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(G257), .B(G1698), .C1(new_n297), .C2(new_n298), .ZN(new_n614));
  OAI211_X1 g0414(.A(G250), .B(new_n296), .C1(new_n297), .C2(new_n298), .ZN(new_n615));
  INV_X1    g0415(.A(G294), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n614), .B(new_n615), .C1(new_n278), .C2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(KEYINPUT84), .A3(new_n302), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n501), .A2(G264), .A3(new_n309), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n619), .A2(new_n506), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT84), .B1(new_n617), .B2(new_n302), .ZN(new_n622));
  OAI21_X1  g0422(.A(G169), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n617), .A2(new_n302), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n620), .A2(new_n624), .A3(G179), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n210), .B(G87), .C1(new_n297), .C2(new_n298), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT22), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT22), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n317), .A2(new_n629), .A3(new_n210), .A4(G87), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT24), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n595), .A2(G20), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT23), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n210), .B2(G107), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n547), .A2(KEYINPUT23), .A3(G20), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n631), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n632), .B1(new_n631), .B2(new_n637), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n270), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n259), .A2(new_n547), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(KEYINPUT25), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n609), .B2(G107), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n626), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n621), .A2(G190), .A3(new_n622), .ZN(new_n646));
  AOI21_X1  g0446(.A(G200), .B1(new_n620), .B2(new_n624), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n640), .B(new_n643), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NOR4_X1   g0449(.A1(new_n486), .A2(new_n526), .A3(new_n613), .A4(new_n649), .ZN(G372));
  OR2_X1    g0450(.A1(new_n323), .A2(new_n325), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n442), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n333), .A2(new_n331), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n315), .A2(new_n321), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n332), .B1(new_n654), .B2(G169), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n286), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n397), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n404), .A2(new_n417), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n659), .A2(new_n482), .B1(new_n465), .B2(new_n467), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n610), .A2(new_n589), .A3(new_n590), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n608), .A2(new_n611), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n661), .A2(new_n662), .B1(new_n591), .B2(new_n604), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n648), .A2(new_n663), .A3(new_n560), .A4(new_n578), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n516), .A2(new_n524), .A3(new_n525), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n623), .A2(new_n625), .B1(new_n640), .B2(new_n643), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n605), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n540), .A2(new_n541), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n577), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT26), .B1(new_n670), .B2(new_n663), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n605), .A2(new_n612), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n672), .A2(new_n560), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n660), .B1(new_n486), .B2(new_n676), .ZN(G369));
  NAND2_X1  g0477(.A1(new_n256), .A2(new_n210), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n520), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n526), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n665), .A2(new_n684), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n683), .B1(new_n640), .B2(new_n643), .ZN(new_n690));
  OAI22_X1  g0490(.A1(new_n649), .A2(new_n690), .B1(new_n645), .B2(new_n683), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n665), .A2(new_n683), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n645), .A2(new_n648), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n693), .A2(new_n694), .B1(new_n666), .B2(new_n683), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(G399));
  OAI21_X1  g0496(.A(new_n683), .B1(new_n668), .B2(new_n675), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(KEYINPUT29), .Z(new_n698));
  INV_X1    g0498(.A(new_n613), .ZN(new_n699));
  INV_X1    g0499(.A(new_n526), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n694), .A2(new_n699), .A3(new_n700), .A4(new_n683), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT86), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n502), .A2(new_n506), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n302), .B2(new_n511), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n399), .B1(new_n596), .B2(new_n598), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n513), .A2(KEYINPUT86), .A3(new_n399), .A4(new_n603), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n567), .A2(new_n570), .B1(new_n620), .B2(new_n624), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  INV_X1    g0510(.A(new_n619), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n711), .A2(new_n596), .A3(new_n598), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n567), .A3(new_n570), .A4(new_n624), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n704), .A2(G179), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n607), .A2(new_n624), .A3(new_n619), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n523), .A2(KEYINPUT30), .A3(new_n539), .A4(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n709), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n683), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT31), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n719), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n701), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n698), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n209), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n213), .A2(G41), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n552), .A2(new_n224), .A3(new_n487), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n729), .A2(G1), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n218), .B2(new_n729), .ZN(new_n733));
  XOR2_X1   g0533(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n734));
  XNOR2_X1  g0534(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n727), .A2(new_n735), .ZN(G364));
  XOR2_X1   g0536(.A(new_n688), .B(KEYINPUT87), .Z(new_n737));
  NOR2_X1   g0537(.A1(new_n212), .A2(G20), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G45), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT88), .Z(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(G1), .A3(new_n729), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n737), .B(new_n741), .C1(G330), .C2(new_n687), .ZN(new_n742));
  INV_X1    g0542(.A(new_n741), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n214), .A2(new_n317), .ZN(new_n744));
  INV_X1    g0544(.A(G355), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n744), .A2(new_n745), .B1(G116), .B2(new_n214), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n251), .A2(new_n497), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n214), .A2(new_n344), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n219), .B2(new_n457), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n746), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n220), .B1(G20), .B2(new_n401), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n743), .B1(new_n750), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G179), .A2(G200), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n210), .B1(new_n758), .B2(G190), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n210), .A2(new_n385), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(new_n399), .A3(G200), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n344), .B1(new_n759), .B2(new_n616), .C1(new_n761), .C2(new_n510), .ZN(new_n762));
  NAND3_X1  g0562(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n385), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n762), .B1(G326), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n210), .A2(G190), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(new_n399), .A3(G200), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT90), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G283), .ZN(new_n769));
  XNOR2_X1  g0569(.A(KEYINPUT33), .B(G317), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT91), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n763), .A2(G190), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(KEYINPUT91), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n399), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n760), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n766), .ZN(new_n778));
  INV_X1    g0578(.A(G311), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n766), .A2(new_n758), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n780), .B1(G329), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n765), .A2(new_n769), .A3(new_n774), .A4(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n759), .A2(new_n226), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n782), .A2(G159), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(KEYINPUT32), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n785), .B(new_n787), .C1(G68), .C2(new_n772), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n768), .A2(G107), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n317), .B1(new_n761), .B2(new_n224), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(KEYINPUT32), .B2(new_n786), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n776), .ZN(new_n793));
  INV_X1    g0593(.A(new_n778), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G58), .A2(new_n793), .B1(new_n794), .B2(G77), .ZN(new_n795));
  INV_X1    g0595(.A(new_n764), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n205), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT89), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n784), .B1(new_n792), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n757), .B1(new_n799), .B2(new_n754), .ZN(new_n800));
  INV_X1    g0600(.A(new_n753), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n687), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n742), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(G396));
  INV_X1    g0604(.A(KEYINPUT93), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n719), .B(new_n805), .C1(new_n437), .C2(new_n440), .ZN(new_n806));
  INV_X1    g0606(.A(new_n429), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n427), .ZN(new_n808));
  INV_X1    g0608(.A(new_n441), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n805), .B(new_n471), .C1(new_n430), .C2(new_n441), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n719), .B1(new_n437), .B2(new_n440), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n697), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n813), .B(new_n683), .C1(new_n668), .C2(new_n675), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n743), .B1(new_n817), .B2(new_n725), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n725), .B2(new_n817), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n754), .A2(new_n751), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT92), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n743), .B1(new_n821), .B2(G77), .ZN(new_n822));
  INV_X1    g0622(.A(new_n761), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n317), .B(new_n785), .C1(G107), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n768), .A2(G87), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n772), .A2(G283), .B1(new_n764), .B2(G303), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n778), .A2(new_n487), .B1(new_n781), .B2(new_n779), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G294), .B2(new_n793), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n824), .A2(new_n825), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n768), .A2(G68), .ZN(new_n830));
  INV_X1    g0630(.A(G132), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n317), .B1(new_n781), .B2(new_n831), .C1(new_n761), .C2(new_n205), .ZN(new_n832));
  INV_X1    g0632(.A(new_n759), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(G58), .B2(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G143), .A2(new_n793), .B1(new_n794), .B2(G159), .ZN(new_n835));
  INV_X1    g0635(.A(G137), .ZN(new_n836));
  INV_X1    g0636(.A(new_n772), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n835), .B1(new_n796), .B2(new_n836), .C1(new_n444), .C2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT34), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n830), .B(new_n834), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n829), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n822), .B1(new_n842), .B2(new_n754), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n813), .B2(new_n752), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n819), .A2(new_n844), .ZN(G384));
  OR2_X1    g0645(.A1(new_n554), .A2(KEYINPUT35), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n554), .A2(KEYINPUT35), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n846), .A2(G116), .A3(new_n221), .A4(new_n847), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT36), .Z(new_n849));
  NAND4_X1  g0649(.A1(new_n219), .A2(G77), .A3(new_n351), .A4(new_n352), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n205), .A2(G68), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n209), .B(G13), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n660), .B1(new_n698), .B2(new_n486), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT95), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT96), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT39), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n413), .A2(new_n415), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n413), .A2(new_n682), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(new_n393), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n858), .A2(new_n859), .A3(new_n862), .A4(new_n393), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT94), .ZN(new_n865));
  INV_X1    g0665(.A(new_n859), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n395), .A2(new_n396), .A3(new_n404), .A4(new_n417), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n864), .A2(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n861), .A2(KEYINPUT94), .A3(new_n863), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT38), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n407), .A2(new_n408), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n343), .B1(new_n871), .B2(new_n367), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n363), .A2(new_n373), .A3(new_n359), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n361), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n342), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n393), .B1(new_n875), .B2(new_n403), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n875), .A2(new_n681), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT37), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n863), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n375), .A2(new_n403), .A3(KEYINPUT18), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n416), .B1(new_n413), .B2(new_n415), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT79), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n404), .A2(new_n417), .A3(new_n405), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n397), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n877), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n879), .B(KEYINPUT38), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n857), .B1(new_n870), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n334), .A2(new_n286), .A3(new_n683), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(KEYINPUT39), .A3(new_n886), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n888), .A2(new_n890), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n886), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n286), .A2(new_n719), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n656), .A2(new_n651), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n286), .B(new_n719), .C1(new_n334), .C2(new_n326), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n442), .A2(new_n683), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n900), .B1(new_n816), .B2(new_n901), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n896), .A2(new_n902), .B1(new_n658), .B2(new_n681), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n895), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n856), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n898), .A2(new_n899), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(new_n724), .A3(new_n813), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n420), .A2(new_n877), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n910), .B2(new_n879), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n909), .B1(new_n911), .B2(new_n887), .ZN(new_n912));
  XOR2_X1   g0712(.A(KEYINPUT97), .B(KEYINPUT40), .Z(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AND4_X1   g0715(.A1(KEYINPUT40), .A2(new_n907), .A3(new_n724), .A4(new_n813), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n870), .B2(new_n887), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n484), .A2(new_n485), .A3(new_n724), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(G330), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n906), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n209), .B2(new_n738), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n906), .A2(new_n923), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n853), .B1(new_n925), .B2(new_n926), .ZN(G367));
  NAND2_X1  g0727(.A1(new_n740), .A2(G1), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT99), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n560), .B(new_n578), .C1(new_n577), .C2(new_n683), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n670), .A2(new_n719), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n695), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT44), .ZN(new_n935));
  INV_X1    g0735(.A(new_n692), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n695), .A2(new_n933), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT45), .ZN(new_n938));
  OR3_X1    g0738(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n936), .B1(new_n935), .B2(new_n938), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n693), .A2(new_n694), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n691), .B2(new_n693), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n688), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n737), .B2(new_n944), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(new_n725), .A3(new_n698), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n726), .B1(new_n942), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n728), .B(KEYINPUT41), .Z(new_n950));
  OAI21_X1  g0750(.A(new_n930), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n933), .ZN(new_n952));
  OR3_X1    g0752(.A1(new_n943), .A2(new_n952), .A3(KEYINPUT42), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n933), .A2(new_n693), .A3(new_n694), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n560), .B1(new_n931), .B2(new_n645), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n954), .A2(KEYINPUT42), .B1(new_n683), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT98), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n661), .A2(new_n683), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(new_n591), .A3(new_n604), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n672), .B2(new_n960), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT43), .Z(new_n963));
  OR2_X1    g0763(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n959), .B1(KEYINPUT43), .B2(new_n962), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n936), .A2(new_n933), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n962), .A2(new_n801), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n755), .B1(new_n214), .B2(new_n434), .C1(new_n247), .C2(new_n748), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n743), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G50), .A2(new_n794), .B1(new_n782), .B2(G137), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n275), .B2(new_n767), .C1(new_n444), .C2(new_n776), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n317), .B1(new_n761), .B2(new_n201), .C1(new_n355), .C2(new_n837), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n759), .A2(new_n202), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n764), .A2(G143), .ZN(new_n976));
  NOR4_X1   g0776(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n761), .A2(new_n487), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT46), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G303), .A2(new_n793), .B1(new_n782), .B2(G317), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n527), .B2(new_n778), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n796), .A2(new_n779), .B1(new_n759), .B2(new_n547), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n344), .B1(new_n767), .B2(new_n226), .C1(new_n616), .C2(new_n837), .ZN(new_n983));
  NOR4_X1   g0783(.A1(new_n979), .A2(new_n981), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n977), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT47), .Z(new_n986));
  AOI21_X1  g0786(.A(new_n971), .B1(new_n986), .B2(new_n754), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n951), .A2(new_n968), .B1(new_n969), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(G387));
  OR2_X1    g0789(.A1(new_n691), .A2(new_n801), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n744), .A2(new_n731), .B1(G107), .B2(new_n214), .ZN(new_n991));
  AOI211_X1 g0791(.A(G45), .B(new_n730), .C1(G68), .C2(G77), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(KEYINPUT100), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(KEYINPUT100), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT50), .B1(new_n338), .B2(G50), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n338), .A2(KEYINPUT50), .A3(G50), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n748), .B1(new_n244), .B2(new_n305), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n991), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n743), .B1(new_n1000), .B2(new_n756), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n833), .A2(new_n435), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n205), .B2(new_n776), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT102), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n317), .B1(new_n778), .B2(new_n202), .C1(new_n796), .C2(new_n355), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n338), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1005), .B1(new_n1006), .B2(new_n772), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n823), .A2(G77), .B1(new_n782), .B2(G150), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT101), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1009), .A2(new_n1008), .B1(new_n768), .B2(G97), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1004), .A2(new_n1007), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(G317), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n776), .A2(new_n1013), .B1(new_n778), .B2(new_n510), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1014), .A2(KEYINPUT103), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(KEYINPUT103), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n772), .A2(G311), .B1(new_n764), .B2(G322), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT48), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n761), .A2(new_n616), .B1(new_n759), .B2(new_n527), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1020), .A2(KEYINPUT49), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n317), .B1(new_n782), .B2(G326), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(new_n487), .C2(new_n767), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT49), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1012), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1001), .B1(new_n1027), .B2(new_n754), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n946), .A2(new_n929), .B1(new_n990), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n947), .A2(new_n728), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n946), .B1(new_n725), .B2(new_n698), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(G393));
  OAI21_X1  g0832(.A(new_n728), .B1(new_n941), .B2(new_n947), .ZN(new_n1033));
  OAI21_X1  g0833(.A(KEYINPUT106), .B1(new_n942), .B2(new_n948), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT106), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n941), .A2(new_n947), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1033), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n952), .A2(new_n753), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n755), .B1(new_n226), .B2(new_n214), .C1(new_n254), .C2(new_n748), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n743), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n793), .A2(G159), .B1(G150), .B2(new_n764), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT51), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n344), .B1(new_n794), .B2(new_n1006), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n823), .A2(G68), .B1(new_n782), .B2(G143), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n759), .A2(new_n275), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n772), .B2(G50), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n825), .A2(new_n1044), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n317), .B1(new_n794), .B2(G294), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n823), .A2(G283), .B1(new_n782), .B2(G322), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n833), .A2(G116), .B1(G303), .B2(new_n772), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n789), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n796), .A2(new_n1013), .B1(new_n776), .B2(new_n779), .ZN(new_n1053));
  XOR2_X1   g0853(.A(KEYINPUT104), .B(KEYINPUT52), .Z(new_n1054));
  XNOR2_X1  g0854(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1043), .A2(new_n1048), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT105), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1041), .B1(new_n1057), .B2(new_n754), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n942), .A2(new_n929), .B1(new_n1039), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1038), .A2(new_n1059), .ZN(G390));
  NAND2_X1  g0860(.A1(new_n816), .A2(new_n901), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n890), .B1(new_n1061), .B2(new_n907), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n864), .A2(new_n865), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n867), .A2(new_n866), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n869), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n892), .ZN(new_n1067));
  AOI21_X1  g0867(.A(KEYINPUT39), .B1(new_n1067), .B2(new_n886), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n893), .A2(KEYINPUT39), .A3(new_n886), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1063), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n722), .A2(new_n723), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n649), .A2(new_n613), .A3(new_n526), .A4(new_n719), .ZN(new_n1072));
  OAI211_X1 g0872(.A(G330), .B(new_n813), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1073), .A2(new_n900), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1067), .A2(new_n886), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n1062), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1070), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(KEYINPUT107), .B1(new_n1073), .B2(new_n900), .ZN(new_n1079));
  INV_X1    g0879(.A(G330), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n719), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT31), .B1(new_n718), .B2(new_n719), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1080), .B1(new_n1083), .B2(new_n701), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT107), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1084), .A2(new_n1085), .A3(new_n813), .A4(new_n907), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1079), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1062), .B1(new_n888), .B2(new_n894), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1076), .A2(new_n1062), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1078), .A2(new_n1091), .A3(new_n929), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n751), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n821), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n741), .B1(new_n1094), .B2(new_n338), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n317), .B(new_n1046), .C1(G87), .C2(new_n823), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n772), .A2(G107), .B1(new_n764), .B2(G283), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n776), .A2(new_n487), .B1(new_n781), .B2(new_n616), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G97), .B2(new_n794), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1096), .A2(new_n830), .A3(new_n1097), .A4(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n761), .A2(new_n444), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  XOR2_X1   g0902(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n1103));
  AOI22_X1  g0903(.A1(new_n1102), .A2(new_n1103), .B1(new_n772), .B2(G137), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1103), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1101), .A2(new_n1105), .B1(new_n764), .B2(G128), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(KEYINPUT54), .B(G143), .ZN(new_n1107));
  INV_X1    g0907(.A(G125), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n778), .A2(new_n1107), .B1(new_n781), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G132), .B2(new_n793), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n317), .B1(new_n767), .B2(new_n205), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G159), .B2(new_n833), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1104), .A2(new_n1106), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1100), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1114), .A2(KEYINPUT112), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(KEYINPUT112), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n754), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1093), .B(new_n1095), .C1(new_n1115), .C2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1092), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT110), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n484), .A2(new_n485), .A3(new_n1084), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n660), .B(new_n1121), .C1(new_n698), .C2(new_n486), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1073), .A2(new_n900), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1087), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n1061), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1084), .A2(KEYINPUT108), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n813), .B1(new_n1084), .B2(KEYINPUT108), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n900), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1061), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(new_n1129), .A3(new_n1075), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1122), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(new_n1078), .A3(new_n1091), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT109), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n1133), .A3(new_n728), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1078), .A2(new_n1091), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1122), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1133), .B1(new_n1132), .B2(new_n728), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1120), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1132), .A2(new_n728), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT109), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1144), .A2(KEYINPUT110), .A3(new_n1139), .A4(new_n1134), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1119), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(G378));
  NAND2_X1  g0947(.A1(new_n450), .A2(new_n682), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT116), .Z(new_n1149));
  INV_X1    g0949(.A(KEYINPUT115), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n482), .A2(new_n1150), .A3(new_n464), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1150), .B1(new_n482), .B2(new_n464), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1149), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n482), .A2(new_n464), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT115), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1149), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n1158), .A3(new_n1151), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1154), .A2(new_n1155), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1155), .B1(new_n1154), .B2(new_n1159), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n751), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n837), .A2(new_n831), .B1(new_n759), .B2(new_n444), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n793), .A2(G128), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n836), .B2(new_n778), .C1(new_n761), .C2(new_n1107), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(G125), .C2(new_n764), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n278), .B(new_n308), .C1(new_n767), .C2(new_n355), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G124), .B2(new_n782), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n344), .A2(new_n308), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n761), .A2(new_n275), .B1(new_n778), .B2(new_n434), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(G283), .C2(new_n782), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n796), .A2(new_n487), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n975), .B(new_n1177), .C1(G97), .C2(new_n772), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n767), .A2(new_n201), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT113), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n776), .A2(new_n547), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT114), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1176), .A2(new_n1178), .A3(new_n1180), .A4(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT58), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1174), .B(new_n205), .C1(G33), .C2(G41), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1173), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n754), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1094), .A2(new_n205), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1163), .A2(new_n743), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n908), .B1(new_n893), .B2(new_n886), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n917), .B(G330), .C1(new_n1193), .C2(new_n913), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n1162), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1162), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n915), .A2(new_n1196), .A3(G330), .A4(new_n917), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n905), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n904), .A2(new_n1195), .A3(new_n1197), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1192), .B1(new_n1201), .B2(new_n929), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1122), .B(KEYINPUT117), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1200), .A2(new_n1199), .B1(new_n1132), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n728), .B1(new_n1204), .B2(KEYINPUT57), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1132), .A2(new_n1203), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1201), .A2(KEYINPUT57), .A3(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1202), .B1(new_n1205), .B2(new_n1207), .ZN(G375));
  NAND2_X1  g1008(.A1(new_n900), .A2(new_n751), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n743), .B1(new_n821), .B2(G68), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n823), .A2(G159), .B1(new_n782), .B2(G128), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT119), .Z(new_n1212));
  OAI22_X1  g1012(.A1(new_n837), .A2(new_n1107), .B1(new_n205), .B2(new_n759), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G132), .B2(new_n764), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n317), .B1(new_n778), .B2(new_n444), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G137), .B2(new_n793), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1212), .A2(new_n1180), .A3(new_n1214), .A4(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n317), .B1(new_n768), .B2(G77), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT118), .Z(new_n1219));
  AOI22_X1  g1019(.A1(G107), .A2(new_n794), .B1(new_n782), .B2(G303), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n226), .B2(new_n761), .C1(new_n527), .C2(new_n776), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1002), .B1(new_n796), .B2(new_n616), .C1(new_n487), .C2(new_n837), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1217), .B1(new_n1219), .B2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1210), .B1(new_n1224), .B2(new_n754), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1136), .A2(new_n929), .B1(new_n1209), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n950), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1138), .A2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1226), .B1(new_n1228), .B2(new_n1229), .ZN(G381));
  OR2_X1    g1030(.A1(G393), .A2(G396), .ZN(new_n1231));
  OR3_X1    g1031(.A1(G390), .A2(G384), .A3(new_n1231), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1232), .A2(G387), .A3(G381), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(G375), .B(KEYINPUT120), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1119), .B1(new_n1235), .B2(new_n1144), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1236), .ZN(G407));
  INV_X1    g1037(.A(G213), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1238), .A2(G343), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1234), .A2(new_n1236), .A3(new_n1239), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1240), .B(KEYINPUT121), .Z(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(G213), .A3(G407), .ZN(G409));
  NAND3_X1  g1042(.A1(new_n1229), .A2(KEYINPUT60), .A3(new_n1138), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n728), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1229), .B1(KEYINPUT60), .B2(new_n1138), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(G384), .B1(new_n1246), .B2(new_n1226), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G384), .B(new_n1226), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1239), .A2(G2897), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1250), .A2(G2897), .A3(new_n1239), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT122), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n904), .A2(new_n1195), .A3(new_n1197), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1195), .A2(new_n1197), .B1(new_n895), .B2(new_n903), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1256), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1199), .A2(KEYINPUT122), .A3(new_n1200), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1260), .A3(new_n929), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1201), .A2(new_n1206), .A3(new_n1227), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n1191), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1236), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1146), .B2(G375), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1239), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT61), .B1(new_n1255), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT62), .B1(new_n1267), .B2(new_n1251), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1265), .A2(KEYINPUT123), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT123), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1272), .B(new_n1264), .C1(new_n1146), .C2(G375), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1271), .A2(new_n1266), .A3(new_n1273), .A4(new_n1250), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(KEYINPUT62), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1231), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1038), .A2(new_n1277), .A3(new_n1059), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1059), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1231), .B(new_n1276), .C1(new_n1037), .C2(new_n1279), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1278), .A2(new_n988), .A3(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n988), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n1270), .A2(new_n1275), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1271), .A2(new_n1266), .A3(new_n1273), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT124), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT124), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1271), .A2(new_n1286), .A3(new_n1266), .A4(new_n1273), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1255), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT125), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1265), .A2(new_n1250), .A3(KEYINPUT63), .A4(new_n1266), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1281), .A2(new_n1282), .A3(KEYINPUT61), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1293), .B2(new_n1274), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1288), .A2(new_n1289), .A3(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1289), .B1(new_n1288), .B2(new_n1294), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1283), .B1(new_n1295), .B2(new_n1296), .ZN(G405));
  NOR2_X1   g1097(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1298));
  AND2_X1   g1098(.A1(G375), .A2(new_n1236), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1146), .A2(G375), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT126), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1250), .A2(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1301), .B(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT127), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1298), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1304), .B(new_n1305), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1306), .B1(new_n1307), .B2(new_n1298), .ZN(G402));
endmodule


