//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n202));
  OR2_X1    g001(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n205));
  NAND4_X1  g004(.A1(new_n203), .A2(KEYINPUT23), .A3(new_n204), .A4(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(new_n204), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n206), .A2(KEYINPUT65), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  MUX2_X1   g013(.A(KEYINPUT24), .B(new_n213), .S(new_n214), .Z(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT65), .B1(new_n206), .B2(new_n211), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n202), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n202), .B1(new_n219), .B2(KEYINPUT23), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n215), .A2(new_n211), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT26), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n219), .B1(new_n223), .B2(new_n207), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n225), .B(new_n226), .C1(KEYINPUT26), .C2(new_n210), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT27), .B(G183gat), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT28), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(KEYINPUT28), .A3(new_n229), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n232), .A2(new_n233), .B1(G183gat), .B2(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n227), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n222), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g036(.A(G113gat), .B(G120gat), .ZN(new_n238));
  INV_X1    g037(.A(G127gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(G134gat), .ZN(new_n240));
  INV_X1    g039(.A(G134gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(G127gat), .ZN(new_n242));
  OAI22_X1  g041(.A1(new_n238), .A2(KEYINPUT1), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G120gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G113gat), .ZN(new_n245));
  INV_X1    g044(.A(G113gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G120gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G127gat), .B(G134gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n243), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G227gat), .A2(G233gat), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n218), .A2(new_n221), .B1(new_n227), .B2(new_n234), .ZN(new_n255));
  INV_X1    g054(.A(new_n252), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT67), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n255), .A2(new_n256), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n253), .B(new_n254), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT34), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n261), .B1(new_n259), .B2(new_n260), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT68), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT32), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n253), .B1(new_n257), .B2(new_n258), .ZN(new_n266));
  INV_X1    g065(.A(new_n254), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT33), .B1(new_n266), .B2(new_n267), .ZN(new_n269));
  XOR2_X1   g068(.A(G15gat), .B(G43gat), .Z(new_n270));
  XNOR2_X1  g069(.A(G71gat), .B(G99gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n268), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  AOI221_X4 g073(.A(new_n265), .B1(KEYINPUT33), .B2(new_n272), .C1(new_n266), .C2(new_n267), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n264), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n263), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n268), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n267), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT33), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n281), .A2(new_n284), .A3(new_n272), .ZN(new_n285));
  INV_X1    g084(.A(new_n275), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n276), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n288), .A2(KEYINPUT36), .ZN(new_n289));
  OAI22_X1  g088(.A1(new_n274), .A2(new_n275), .B1(new_n263), .B2(new_n262), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n285), .A2(new_n286), .A3(new_n277), .A4(new_n279), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT36), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G8gat), .B(G36gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT71), .ZN(new_n295));
  XOR2_X1   g094(.A(G64gat), .B(G92gat), .Z(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT72), .ZN(new_n298));
  AND2_X1   g097(.A1(G226gat), .A2(G233gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n236), .A2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(KEYINPUT70), .B(KEYINPUT29), .Z(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n255), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n300), .B1(new_n303), .B2(new_n299), .ZN(new_n304));
  XNOR2_X1  g103(.A(G197gat), .B(G204gat), .ZN(new_n305));
  INV_X1    g104(.A(G211gat), .ZN(new_n306));
  INV_X1    g105(.A(G218gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n305), .B1(KEYINPUT22), .B2(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(G211gat), .B(G218gat), .Z(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n304), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n255), .A2(KEYINPUT29), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n300), .B(new_n311), .C1(new_n315), .C2(new_n299), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n298), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n313), .A2(KEYINPUT30), .A3(new_n316), .A4(new_n297), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT73), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n313), .A2(new_n316), .A3(new_n297), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(KEYINPUT30), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n318), .A2(new_n319), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT6), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT78), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n243), .A2(new_n251), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n330), .B1(new_n243), .B2(new_n251), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G155gat), .B(G162gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT2), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(G155gat), .B2(G162gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(G141gat), .B(G148gat), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(KEYINPUT74), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n339));
  INV_X1    g138(.A(G148gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(G141gat), .ZN(new_n341));
  INV_X1    g140(.A(G141gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(G148gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n339), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n334), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT2), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT76), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n346), .A2(KEYINPUT76), .A3(KEYINPUT2), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n334), .A3(new_n350), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n342), .A2(KEYINPUT75), .A3(G148gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n340), .A2(G141gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n340), .B2(G141gat), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n352), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT3), .B1(new_n345), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n342), .A2(G148gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(new_n353), .A3(KEYINPUT74), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n360), .A3(new_n347), .ZN(new_n361));
  INV_X1    g160(.A(new_n334), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n355), .A2(new_n353), .ZN(new_n364));
  INV_X1    g163(.A(new_n352), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n366), .A2(new_n334), .A3(new_n350), .A4(new_n349), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n363), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n333), .A2(new_n358), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G225gat), .A2(G233gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n256), .A2(new_n363), .A3(new_n367), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n345), .A2(new_n357), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(KEYINPUT4), .A3(new_n256), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n370), .A2(new_n371), .A3(new_n374), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n252), .A2(KEYINPUT77), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n243), .A2(new_n251), .A3(new_n330), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n372), .B1(new_n380), .B2(new_n375), .ZN(new_n381));
  INV_X1    g180(.A(new_n371), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT5), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT5), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n377), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT0), .ZN(new_n390));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  AOI21_X1  g191(.A(new_n329), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n377), .A2(new_n386), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n386), .B1(new_n377), .B2(new_n383), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n329), .B(new_n392), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n328), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT79), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n400), .B(new_n328), .C1(new_n393), .C2(new_n397), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n388), .A2(new_n392), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n328), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n327), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n311), .A2(new_n301), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n375), .B1(new_n409), .B2(new_n368), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n311), .B1(new_n369), .B2(new_n301), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT29), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT3), .B1(new_n311), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n415), .B2(new_n375), .ZN(new_n416));
  OAI22_X1  g215(.A1(new_n412), .A2(new_n413), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(G22gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(G78gat), .B(G106gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT31), .B(G50gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  MUX2_X1   g221(.A(G22gat), .B(new_n419), .S(new_n422), .Z(new_n423));
  XNOR2_X1  g222(.A(new_n417), .B(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n293), .B1(new_n408), .B2(new_n424), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n425), .A2(KEYINPUT81), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT37), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n313), .A2(new_n427), .A3(new_n316), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT85), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n313), .A2(KEYINPUT85), .A3(new_n427), .A4(new_n316), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n297), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT37), .B1(new_n314), .B2(new_n317), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT38), .ZN(new_n436));
  INV_X1    g235(.A(new_n298), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n300), .B(new_n312), .C1(new_n315), .C2(new_n299), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n427), .B1(new_n304), .B2(new_n311), .ZN(new_n439));
  AOI211_X1 g238(.A(KEYINPUT38), .B(new_n437), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n322), .B1(new_n432), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n398), .A2(new_n403), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n407), .ZN(new_n444));
  OR2_X1    g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n322), .A2(KEYINPUT30), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n446), .A2(new_n318), .A3(new_n319), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT39), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n381), .A2(new_n382), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT83), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n370), .A2(new_n374), .A3(new_n376), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n382), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n451), .B(new_n453), .C1(new_n450), .C2(new_n449), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n392), .B1(new_n453), .B2(KEYINPUT39), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT82), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(KEYINPUT82), .B(new_n392), .C1(new_n453), .C2(KEYINPUT39), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n454), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT40), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n403), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n459), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT84), .B1(new_n462), .B2(KEYINPUT40), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT84), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n459), .A2(new_n464), .A3(new_n460), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n447), .B(new_n461), .C1(new_n463), .C2(new_n465), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n466), .A2(new_n424), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n425), .A2(KEYINPUT81), .B1(new_n445), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n326), .A2(new_n325), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n469), .A2(new_n323), .A3(new_n320), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n276), .A2(new_n287), .A3(new_n424), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n403), .B1(new_n399), .B2(new_n401), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(new_n406), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT86), .B1(new_n473), .B2(KEYINPUT35), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n473), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n290), .A2(new_n291), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(new_n447), .ZN(new_n480));
  INV_X1    g279(.A(new_n424), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(KEYINPUT35), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n444), .A3(new_n482), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n426), .A2(new_n468), .B1(new_n477), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT16), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n485), .A2(G1gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(G15gat), .B(G22gat), .ZN(new_n487));
  MUX2_X1   g286(.A(G1gat), .B(new_n486), .S(new_n487), .Z(new_n488));
  INV_X1    g287(.A(G8gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(G57gat), .A2(G64gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(G57gat), .A2(G64gat), .ZN(new_n492));
  AND2_X1   g291(.A1(G71gat), .A2(G78gat), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n491), .B(new_n492), .C1(new_n493), .C2(KEYINPUT9), .ZN(new_n494));
  XNOR2_X1  g293(.A(G71gat), .B(G78gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n490), .B1(KEYINPUT21), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n496), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT94), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G231gat), .A2(G233gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G127gat), .B(G155gat), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n505), .B(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n505), .B(new_n506), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n509), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n498), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n511), .A2(new_n513), .A3(new_n498), .ZN(new_n516));
  XOR2_X1   g315(.A(G183gat), .B(G211gat), .Z(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n516), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n517), .B1(new_n520), .B2(new_n514), .ZN(new_n521));
  XNOR2_X1  g320(.A(G190gat), .B(G218gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G43gat), .B(G50gat), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n524), .A2(KEYINPUT15), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n525), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(G29gat), .A2(G36gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT14), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n526), .B(new_n529), .C1(KEYINPUT15), .C2(new_n524), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n529), .A2(KEYINPUT87), .ZN(new_n531));
  NAND2_X1  g330(.A1(G29gat), .A2(G36gat), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(new_n529), .B2(KEYINPUT87), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n525), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g335(.A1(G85gat), .A2(G92gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(G99gat), .A2(G106gat), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n536), .A2(new_n537), .B1(new_n538), .B2(KEYINPUT8), .ZN(new_n539));
  NAND3_X1  g338(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT96), .B(G92gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(G85gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G99gat), .B(G106gat), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n544), .B(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT41), .ZN(new_n548));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549));
  OAI22_X1  g348(.A1(new_n535), .A2(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT97), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n530), .A2(new_n534), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(new_n535), .B2(KEYINPUT17), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n553), .A2(KEYINPUT88), .A3(new_n554), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n547), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n523), .B1(new_n552), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n561), .A2(KEYINPUT98), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n552), .A2(new_n560), .A3(new_n523), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n561), .B2(KEYINPUT98), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT95), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n548), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n568), .ZN(new_n570));
  OAI211_X1 g369(.A(KEYINPUT95), .B(new_n570), .C1(new_n562), .C2(new_n564), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n519), .A2(new_n521), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT89), .ZN(new_n573));
  INV_X1    g372(.A(new_n490), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n559), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT88), .B1(new_n553), .B2(new_n554), .ZN(new_n576));
  AOI211_X1 g375(.A(new_n556), .B(KEYINPUT17), .C1(new_n530), .C2(new_n534), .ZN(new_n577));
  OAI22_X1  g376(.A1(new_n576), .A2(new_n577), .B1(new_n554), .B2(new_n553), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT89), .B1(new_n578), .B2(new_n490), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n574), .A2(new_n535), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n575), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT92), .ZN(new_n583));
  NAND2_X1  g382(.A1(G229gat), .A2(G233gat), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT18), .A4(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n575), .A2(new_n579), .A3(new_n584), .A4(new_n581), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT18), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT92), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n553), .B(new_n490), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n584), .B(KEYINPUT13), .Z(new_n590));
  AOI22_X1  g389(.A1(new_n585), .A2(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT90), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n582), .A2(new_n592), .A3(new_n584), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n586), .A2(KEYINPUT90), .ZN(new_n594));
  XOR2_X1   g393(.A(KEYINPUT91), .B(KEYINPUT18), .Z(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G113gat), .B(G141gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT11), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(new_n209), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G197gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n600), .B(KEYINPUT12), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n591), .A2(new_n596), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n602), .B1(new_n591), .B2(new_n596), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G230gat), .ZN(new_n607));
  INV_X1    g406(.A(G233gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT99), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n546), .B1(new_n544), .B2(new_n610), .ZN(new_n611));
  OAI211_X1 g410(.A(KEYINPUT99), .B(new_n545), .C1(new_n541), .C2(new_n543), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n611), .A2(new_n496), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n547), .A2(new_n499), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n547), .A2(new_n619), .A3(new_n499), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT101), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n609), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n618), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n609), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n630), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n624), .A2(new_n626), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n572), .A2(new_n606), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n484), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n405), .A2(new_n407), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G1gat), .ZN(G1324gat));
  INV_X1    g440(.A(new_n447), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n484), .A2(new_n642), .A3(new_n636), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT42), .B1(new_n643), .B2(new_n489), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT16), .B(G8gat), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  MUX2_X1   g445(.A(KEYINPUT42), .B(new_n644), .S(new_n646), .Z(G1325gat));
  INV_X1    g446(.A(G15gat), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n637), .A2(new_n648), .A3(new_n478), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n484), .A2(new_n293), .A3(new_n636), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n649), .B1(new_n650), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT102), .ZN(G1326gat));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n481), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT43), .B(G22gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  NAND2_X1  g454(.A1(new_n569), .A2(new_n571), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n484), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(G29gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n519), .A2(new_n521), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n605), .A2(new_n659), .A3(new_n634), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n657), .A2(new_n658), .A3(new_n639), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT45), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n473), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n483), .B1(new_n663), .B2(new_n474), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI211_X1 g465(.A(KEYINPUT104), .B(new_n483), .C1(new_n663), .C2(new_n474), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n424), .B(new_n466), .C1(new_n442), .C2(new_n444), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n668), .B(new_n293), .C1(new_n408), .C2(new_n424), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  INV_X1    g470(.A(new_n656), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n670), .A2(KEYINPUT105), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT44), .B1(new_n484), .B2(new_n656), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n669), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n664), .B2(new_n665), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n656), .B1(new_n677), .B2(new_n667), .ZN(new_n678));
  AOI21_X1  g477(.A(KEYINPUT105), .B1(new_n678), .B2(new_n671), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n660), .B(KEYINPUT103), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n639), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n662), .B1(new_n683), .B2(new_n658), .ZN(G1328gat));
  NAND2_X1  g483(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  OAI21_X1  g484(.A(G36gat), .B1(new_n685), .B2(new_n642), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n642), .A2(G36gat), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n657), .A2(new_n660), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT46), .Z(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(G1329gat));
  INV_X1    g489(.A(new_n293), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n680), .A2(G43gat), .A3(new_n691), .A4(new_n681), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n657), .A2(new_n478), .A3(new_n660), .ZN(new_n693));
  INV_X1    g492(.A(G43gat), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n696));
  AND3_X1   g495(.A1(new_n692), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n692), .B2(new_n695), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(G1330gat));
  NAND3_X1  g498(.A1(new_n657), .A2(new_n481), .A3(new_n660), .ZN(new_n700));
  INV_X1    g499(.A(G50gat), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n481), .A2(G50gat), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n685), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT48), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n702), .B(new_n706), .C1(new_n685), .C2(new_n703), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(G1331gat));
  NAND3_X1  g507(.A1(new_n572), .A2(new_n605), .A3(new_n634), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT107), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n670), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n639), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g514(.A(new_n711), .B(KEYINPUT108), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT109), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n642), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT110), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n717), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n722), .B(new_n723), .Z(G1333gat));
  INV_X1    g523(.A(G71gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n478), .B(KEYINPUT111), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n716), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n717), .A2(new_n719), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n691), .A2(G71gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT50), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n733), .B(new_n728), .C1(new_n729), .C2(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1334gat));
  NAND3_X1  g534(.A1(new_n717), .A2(new_n719), .A3(new_n481), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G78gat), .ZN(G1335gat));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n606), .A2(new_n659), .A3(new_n635), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n680), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n740), .B2(new_n638), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n680), .A2(KEYINPUT112), .A3(new_n639), .A4(new_n739), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n741), .A2(G85gat), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n638), .A2(G85gat), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n606), .A2(new_n659), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n670), .A2(new_n672), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT51), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n678), .A2(new_n748), .A3(new_n745), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n750), .A2(KEYINPUT113), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(KEYINPUT113), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n634), .B(new_n744), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n743), .A2(new_n753), .ZN(G1336gat));
  OAI211_X1 g553(.A(new_n447), .B(new_n739), .C1(new_n675), .C2(new_n679), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n542), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n635), .A2(G92gat), .A3(new_n642), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n756), .B(new_n757), .C1(new_n750), .C2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n761), .A3(new_n748), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n678), .B(new_n745), .C1(KEYINPUT115), .C2(KEYINPUT51), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n758), .B(KEYINPUT114), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT116), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n764), .A2(new_n768), .A3(new_n765), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n767), .A2(new_n756), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n760), .B1(new_n770), .B2(new_n757), .ZN(G1337gat));
  OAI21_X1  g570(.A(G99gat), .B1(new_n740), .B2(new_n293), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n479), .A2(G99gat), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n634), .B(new_n773), .C1(new_n751), .C2(new_n752), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(G1338gat));
  INV_X1    g574(.A(KEYINPUT118), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n481), .B(new_n739), .C1(new_n675), .C2(new_n679), .ZN(new_n778));
  XOR2_X1   g577(.A(KEYINPUT117), .B(G106gat), .Z(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n635), .A2(G106gat), .A3(new_n424), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n777), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n747), .A2(new_n749), .A3(new_n781), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n777), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n778), .B2(new_n779), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n776), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n785), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n780), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n778), .A2(new_n779), .B1(new_n764), .B2(new_n781), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n789), .B(KEYINPUT118), .C1(new_n777), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(G1339gat));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n620), .A2(new_n622), .A3(new_n609), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n624), .A2(KEYINPUT54), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n632), .B1(new_n623), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n795), .A2(KEYINPUT55), .A3(new_n797), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n633), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n603), .B2(new_n604), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n591), .A2(new_n596), .A3(new_n602), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n582), .A2(new_n584), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n589), .A2(new_n590), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n600), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n634), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n672), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n805), .A2(new_n808), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n811), .A2(new_n672), .A3(new_n803), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n793), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n591), .A2(new_n596), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n601), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n802), .B1(new_n815), .B2(new_n805), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n805), .A2(new_n634), .A3(new_n808), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n656), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n811), .A2(new_n672), .A3(new_n803), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(KEYINPUT119), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n659), .B1(new_n813), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n572), .A2(new_n605), .A3(new_n635), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n824), .A2(new_n639), .A3(new_n424), .A4(new_n480), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n825), .A2(new_n246), .A3(new_n605), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n639), .B1(new_n821), .B2(new_n823), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n827), .A2(new_n481), .A3(new_n288), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n642), .A3(new_n606), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n826), .B1(new_n829), .B2(new_n246), .ZN(G1340gat));
  NOR3_X1   g629(.A1(new_n825), .A2(new_n244), .A3(new_n635), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n642), .A3(new_n634), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(new_n244), .ZN(G1341gat));
  INV_X1    g632(.A(new_n659), .ZN(new_n834));
  OAI21_X1  g633(.A(G127gat), .B1(new_n825), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n828), .A2(new_n642), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n659), .A2(new_n239), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(G1342gat));
  OAI21_X1  g637(.A(G134gat), .B1(new_n825), .B2(new_n656), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n656), .A2(new_n447), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT120), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(G134gat), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n828), .A2(KEYINPUT56), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT56), .B1(new_n828), .B2(new_n842), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n839), .B1(new_n843), .B2(new_n844), .ZN(G1343gat));
  NAND2_X1  g644(.A1(new_n827), .A2(KEYINPUT121), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n847), .B(new_n639), .C1(new_n821), .C2(new_n823), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n691), .A2(new_n424), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n846), .A2(new_n642), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n342), .B1(new_n850), .B2(new_n605), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n824), .A2(new_n852), .A3(new_n481), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n691), .A2(new_n638), .A3(new_n447), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n818), .A2(new_n819), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n823), .B1(new_n855), .B2(new_n834), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT57), .B1(new_n856), .B2(new_n424), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n853), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n606), .A2(G141gat), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n851), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n851), .B(KEYINPUT58), .C1(new_n858), .C2(new_n859), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1344gat));
  NOR2_X1   g663(.A1(new_n858), .A2(new_n635), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n865), .A2(KEYINPUT59), .A3(new_n340), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867));
  OAI211_X1 g666(.A(KEYINPUT57), .B(new_n481), .C1(new_n821), .C2(new_n823), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n834), .B1(new_n810), .B2(new_n812), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n424), .B1(new_n870), .B2(new_n822), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n869), .B1(new_n871), .B2(KEYINPUT57), .ZN(new_n872));
  OAI211_X1 g671(.A(KEYINPUT122), .B(new_n852), .C1(new_n856), .C2(new_n424), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n868), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n634), .A3(new_n854), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n867), .B1(new_n875), .B2(G148gat), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n634), .A2(new_n340), .ZN(new_n877));
  OAI22_X1  g676(.A1(new_n866), .A2(new_n876), .B1(new_n850), .B2(new_n877), .ZN(G1345gat));
  INV_X1    g677(.A(G155gat), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n858), .A2(new_n879), .A3(new_n834), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n850), .A2(new_n834), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(KEYINPUT123), .ZN(new_n882));
  AOI21_X1  g681(.A(G155gat), .B1(new_n881), .B2(KEYINPUT123), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(G1346gat));
  OAI21_X1  g683(.A(G162gat), .B1(new_n858), .B2(new_n656), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n841), .A2(G162gat), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n846), .A2(new_n848), .A3(new_n849), .A4(new_n886), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n887), .A2(KEYINPUT124), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(KEYINPUT124), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n885), .A2(new_n888), .A3(new_n889), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n639), .A2(new_n642), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n824), .A2(new_n424), .A3(new_n726), .A4(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(G169gat), .B1(new_n892), .B2(new_n605), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n824), .A2(new_n471), .A3(new_n891), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n606), .A2(new_n203), .A3(new_n205), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(G1348gat));
  OAI21_X1  g695(.A(G176gat), .B1(new_n892), .B2(new_n635), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n634), .A2(new_n204), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n894), .B2(new_n898), .ZN(G1349gat));
  OAI21_X1  g698(.A(G183gat), .B1(new_n892), .B2(new_n834), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n659), .A2(new_n228), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n894), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT60), .ZN(G1350gat));
  OR2_X1    g702(.A1(new_n892), .A2(new_n656), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n905), .A3(G190gat), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n905), .B1(new_n904), .B2(G190gat), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n672), .A2(new_n229), .ZN(new_n909));
  OAI22_X1  g708(.A1(new_n907), .A2(new_n908), .B1(new_n894), .B2(new_n909), .ZN(G1351gat));
  NAND3_X1  g709(.A1(new_n824), .A2(new_n849), .A3(new_n891), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(KEYINPUT125), .B(G197gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n606), .A3(new_n913), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n691), .A2(new_n639), .A3(new_n642), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n874), .A2(new_n606), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n914), .B1(new_n916), .B2(new_n913), .ZN(G1352gat));
  NOR3_X1   g716(.A1(new_n911), .A2(G204gat), .A3(new_n635), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT62), .ZN(new_n919));
  INV_X1    g718(.A(G204gat), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n874), .A2(new_n634), .A3(new_n915), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(G1353gat));
  NAND3_X1  g721(.A1(new_n874), .A2(new_n659), .A3(new_n915), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n923), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n923), .A2(G211gat), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT63), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n926), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n912), .A2(new_n306), .A3(new_n659), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1354gat));
  NAND3_X1  g732(.A1(new_n912), .A2(new_n307), .A3(new_n672), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n874), .A2(new_n672), .A3(new_n915), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n935), .B2(new_n307), .ZN(G1355gat));
endmodule


