

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U545 ( .A1(n572), .A2(n517), .ZN(n791) );
  AND2_X1 U546 ( .A1(n530), .A2(G2104), .ZN(n868) );
  NAND2_X1 U547 ( .A1(n603), .A2(n602), .ZN(n966) );
  NOR2_X2 U548 ( .A1(n600), .A2(n599), .ZN(n601) );
  AND2_X2 U549 ( .A1(G160), .A2(G40), .ZN(n699) );
  AND2_X1 U550 ( .A1(n544), .A2(n543), .ZN(G164) );
  BUF_X1 U551 ( .A(n683), .Z(n684) );
  NOR2_X1 U552 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  BUF_X2 U553 ( .A(n869), .Z(n511) );
  XOR2_X1 U554 ( .A(KEYINPUT17), .B(n527), .Z(n869) );
  INV_X1 U555 ( .A(KEYINPUT29), .ZN(n633) );
  AND2_X1 U556 ( .A1(n636), .A2(G1996), .ZN(n591) );
  AND2_X1 U557 ( .A1(n641), .A2(G8), .ZN(n643) );
  XNOR2_X1 U558 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U559 ( .A(n649), .B(KEYINPUT102), .ZN(n650) );
  AND2_X1 U560 ( .A1(G2105), .A2(G2104), .ZN(n872) );
  NAND2_X1 U561 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U562 ( .A(n634), .B(n633), .ZN(n640) );
  INV_X2 U563 ( .A(n654), .ZN(n636) );
  XOR2_X1 U564 ( .A(KEYINPUT87), .B(n541), .Z(n512) );
  INV_X1 U565 ( .A(KEYINPUT30), .ZN(n642) );
  NOR2_X1 U566 ( .A1(G168), .A2(n644), .ZN(n645) );
  INV_X1 U567 ( .A(KEYINPUT31), .ZN(n649) );
  NAND2_X1 U568 ( .A1(G8), .A2(n654), .ZN(n715) );
  XNOR2_X1 U569 ( .A(KEYINPUT71), .B(KEYINPUT13), .ZN(n597) );
  XNOR2_X1 U570 ( .A(n598), .B(n597), .ZN(n599) );
  NOR2_X1 U571 ( .A1(G651), .A2(n572), .ZN(n787) );
  XOR2_X1 U572 ( .A(KEYINPUT1), .B(n518), .Z(n786) );
  INV_X1 U573 ( .A(KEYINPUT88), .ZN(n539) );
  XNOR2_X1 U574 ( .A(n540), .B(n539), .ZN(n544) );
  NOR2_X1 U575 ( .A1(G651), .A2(G543), .ZN(n790) );
  NAND2_X1 U576 ( .A1(n790), .A2(G89), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(KEYINPUT4), .ZN(n515) );
  XOR2_X1 U578 ( .A(KEYINPUT0), .B(G543), .Z(n572) );
  INV_X1 U579 ( .A(G651), .ZN(n517) );
  NAND2_X1 U580 ( .A1(G76), .A2(n791), .ZN(n514) );
  NAND2_X1 U581 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(KEYINPUT5), .B(n516), .ZN(n524) );
  NOR2_X1 U583 ( .A1(G543), .A2(n517), .ZN(n518) );
  NAND2_X1 U584 ( .A1(G63), .A2(n786), .ZN(n520) );
  NAND2_X1 U585 ( .A1(G51), .A2(n787), .ZN(n519) );
  NAND2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n522) );
  XOR2_X1 U587 ( .A(KEYINPUT74), .B(KEYINPUT6), .Z(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(n523) );
  NAND2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U590 ( .A(KEYINPUT7), .B(n525), .ZN(G168) );
  INV_X1 U591 ( .A(G2105), .ZN(n530) );
  NOR2_X1 U592 ( .A1(n530), .A2(G2104), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n526), .B(KEYINPUT66), .ZN(n683) );
  NAND2_X1 U594 ( .A1(n683), .A2(G125), .ZN(n535) );
  NAND2_X1 U595 ( .A1(G137), .A2(n511), .ZN(n529) );
  NAND2_X1 U596 ( .A1(G113), .A2(n872), .ZN(n528) );
  NAND2_X1 U597 ( .A1(n529), .A2(n528), .ZN(n533) );
  NAND2_X1 U598 ( .A1(G101), .A2(n868), .ZN(n531) );
  XNOR2_X1 U599 ( .A(KEYINPUT23), .B(n531), .ZN(n532) );
  NOR2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X2 U601 ( .A(n536), .B(KEYINPUT65), .ZN(G160) );
  NAND2_X1 U602 ( .A1(G102), .A2(n868), .ZN(n538) );
  NAND2_X1 U603 ( .A1(G138), .A2(n511), .ZN(n537) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n540) );
  NAND2_X1 U605 ( .A1(G126), .A2(n683), .ZN(n542) );
  NAND2_X1 U606 ( .A1(G114), .A2(n872), .ZN(n541) );
  AND2_X1 U607 ( .A1(n542), .A2(n512), .ZN(n543) );
  NAND2_X1 U608 ( .A1(G65), .A2(n786), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n545), .B(KEYINPUT68), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G91), .A2(n790), .ZN(n547) );
  NAND2_X1 U611 ( .A1(G53), .A2(n787), .ZN(n546) );
  NAND2_X1 U612 ( .A1(n547), .A2(n546), .ZN(n550) );
  NAND2_X1 U613 ( .A1(G78), .A2(n791), .ZN(n548) );
  XNOR2_X1 U614 ( .A(KEYINPUT67), .B(n548), .ZN(n549) );
  NOR2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U617 ( .A(KEYINPUT69), .B(n553), .Z(G299) );
  NAND2_X1 U618 ( .A1(G64), .A2(n786), .ZN(n555) );
  NAND2_X1 U619 ( .A1(G52), .A2(n787), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n560) );
  NAND2_X1 U621 ( .A1(G90), .A2(n790), .ZN(n557) );
  NAND2_X1 U622 ( .A1(G77), .A2(n791), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(G171) );
  XOR2_X1 U626 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U627 ( .A1(G88), .A2(n790), .ZN(n562) );
  NAND2_X1 U628 ( .A1(G75), .A2(n791), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G62), .A2(n786), .ZN(n563) );
  XOR2_X1 U631 ( .A(KEYINPUT81), .B(n563), .Z(n565) );
  NAND2_X1 U632 ( .A1(n787), .A2(G50), .ZN(n564) );
  NAND2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U634 ( .A1(n567), .A2(n566), .ZN(G166) );
  XNOR2_X1 U635 ( .A(KEYINPUT89), .B(G166), .ZN(G303) );
  NAND2_X1 U636 ( .A1(G49), .A2(n787), .ZN(n569) );
  NAND2_X1 U637 ( .A1(G74), .A2(G651), .ZN(n568) );
  NAND2_X1 U638 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U639 ( .A(KEYINPUT78), .B(n570), .ZN(n571) );
  NOR2_X1 U640 ( .A1(n786), .A2(n571), .ZN(n574) );
  NAND2_X1 U641 ( .A1(n572), .A2(G87), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(G288) );
  NAND2_X1 U643 ( .A1(G73), .A2(n791), .ZN(n575) );
  XOR2_X1 U644 ( .A(KEYINPUT79), .B(n575), .Z(n576) );
  XNOR2_X1 U645 ( .A(n576), .B(KEYINPUT2), .ZN(n578) );
  NAND2_X1 U646 ( .A1(G61), .A2(n786), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U648 ( .A1(G86), .A2(n790), .ZN(n580) );
  NAND2_X1 U649 ( .A1(G48), .A2(n787), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U652 ( .A(KEYINPUT80), .B(n583), .Z(G305) );
  NAND2_X1 U653 ( .A1(G85), .A2(n790), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G72), .A2(n791), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U656 ( .A1(G60), .A2(n786), .ZN(n587) );
  NAND2_X1 U657 ( .A1(G47), .A2(n787), .ZN(n586) );
  NAND2_X1 U658 ( .A1(n587), .A2(n586), .ZN(n588) );
  OR2_X1 U659 ( .A1(n589), .A2(n588), .ZN(G290) );
  NOR2_X1 U660 ( .A1(G164), .A2(G1384), .ZN(n701) );
  NAND2_X2 U661 ( .A1(n699), .A2(n701), .ZN(n654) );
  XOR2_X1 U662 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n590) );
  XNOR2_X1 U663 ( .A(n591), .B(n590), .ZN(n606) );
  AND2_X1 U664 ( .A1(n654), .A2(G1341), .ZN(n604) );
  XOR2_X1 U665 ( .A(KEYINPUT14), .B(KEYINPUT70), .Z(n593) );
  NAND2_X1 U666 ( .A1(G56), .A2(n786), .ZN(n592) );
  XNOR2_X1 U667 ( .A(n593), .B(n592), .ZN(n600) );
  NAND2_X1 U668 ( .A1(n790), .A2(G81), .ZN(n594) );
  XNOR2_X1 U669 ( .A(n594), .B(KEYINPUT12), .ZN(n596) );
  NAND2_X1 U670 ( .A1(G68), .A2(n791), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n598) );
  XNOR2_X1 U672 ( .A(n601), .B(KEYINPUT72), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G43), .A2(n787), .ZN(n602) );
  NOR2_X1 U674 ( .A1(n604), .A2(n966), .ZN(n605) );
  AND2_X1 U675 ( .A1(n606), .A2(n605), .ZN(n619) );
  NAND2_X1 U676 ( .A1(G66), .A2(n786), .ZN(n608) );
  NAND2_X1 U677 ( .A1(G92), .A2(n790), .ZN(n607) );
  NAND2_X1 U678 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U679 ( .A1(G79), .A2(n791), .ZN(n610) );
  NAND2_X1 U680 ( .A1(G54), .A2(n787), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U683 ( .A(KEYINPUT15), .B(n613), .Z(n969) );
  NAND2_X1 U684 ( .A1(n619), .A2(n969), .ZN(n617) );
  NOR2_X1 U685 ( .A1(n636), .A2(G1348), .ZN(n615) );
  NOR2_X1 U686 ( .A1(G2067), .A2(n654), .ZN(n614) );
  NOR2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n618), .B(KEYINPUT100), .ZN(n621) );
  OR2_X1 U690 ( .A1(n619), .A2(n969), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n621), .A2(n620), .ZN(n626) );
  INV_X1 U692 ( .A(G299), .ZN(n628) );
  NAND2_X1 U693 ( .A1(n636), .A2(G2072), .ZN(n622) );
  XNOR2_X1 U694 ( .A(n622), .B(KEYINPUT27), .ZN(n624) );
  INV_X1 U695 ( .A(G1956), .ZN(n981) );
  NOR2_X1 U696 ( .A1(n981), .A2(n636), .ZN(n623) );
  NOR2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U698 ( .A1(n628), .A2(n627), .ZN(n625) );
  NAND2_X1 U699 ( .A1(n626), .A2(n625), .ZN(n632) );
  NOR2_X1 U700 ( .A1(n628), .A2(n627), .ZN(n630) );
  XNOR2_X1 U701 ( .A(KEYINPUT99), .B(KEYINPUT28), .ZN(n629) );
  XNOR2_X1 U702 ( .A(n630), .B(n629), .ZN(n631) );
  NAND2_X1 U703 ( .A1(n632), .A2(n631), .ZN(n634) );
  NOR2_X1 U704 ( .A1(n636), .A2(G1961), .ZN(n635) );
  XOR2_X1 U705 ( .A(KEYINPUT98), .B(n635), .Z(n638) );
  XNOR2_X1 U706 ( .A(G2078), .B(KEYINPUT25), .ZN(n939) );
  NAND2_X1 U707 ( .A1(n636), .A2(n939), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n638), .A2(n637), .ZN(n646) );
  NAND2_X1 U709 ( .A1(n646), .A2(G171), .ZN(n639) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n653) );
  NOR2_X1 U711 ( .A1(G1966), .A2(n715), .ZN(n666) );
  NOR2_X1 U712 ( .A1(G2084), .A2(n654), .ZN(n667) );
  NOR2_X1 U713 ( .A1(n666), .A2(n667), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U715 ( .A(KEYINPUT101), .B(n645), .ZN(n648) );
  OR2_X1 U716 ( .A1(G171), .A2(n646), .ZN(n647) );
  AND2_X1 U717 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U718 ( .A1(n653), .A2(n652), .ZN(n664) );
  NAND2_X1 U719 ( .A1(n664), .A2(G286), .ZN(n661) );
  NOR2_X1 U720 ( .A1(G2090), .A2(n654), .ZN(n655) );
  XOR2_X1 U721 ( .A(KEYINPUT105), .B(n655), .Z(n657) );
  NOR2_X1 U722 ( .A1(G1971), .A2(n715), .ZN(n656) );
  NOR2_X1 U723 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U724 ( .A(n658), .B(KEYINPUT106), .ZN(n659) );
  NAND2_X1 U725 ( .A1(n659), .A2(G303), .ZN(n660) );
  NAND2_X1 U726 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U727 ( .A1(n662), .A2(G8), .ZN(n663) );
  XNOR2_X1 U728 ( .A(KEYINPUT32), .B(n663), .ZN(n672) );
  XNOR2_X1 U729 ( .A(n664), .B(KEYINPUT103), .ZN(n665) );
  NOR2_X1 U730 ( .A1(n666), .A2(n665), .ZN(n669) );
  NAND2_X1 U731 ( .A1(G8), .A2(n667), .ZN(n668) );
  NAND2_X1 U732 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U733 ( .A(n670), .B(KEYINPUT104), .ZN(n671) );
  NAND2_X1 U734 ( .A1(n672), .A2(n671), .ZN(n711) );
  NOR2_X1 U735 ( .A1(G1976), .A2(G288), .ZN(n955) );
  NOR2_X1 U736 ( .A1(G1971), .A2(G303), .ZN(n962) );
  NOR2_X1 U737 ( .A1(n955), .A2(n962), .ZN(n673) );
  NAND2_X1 U738 ( .A1(n711), .A2(n673), .ZN(n675) );
  NAND2_X1 U739 ( .A1(G288), .A2(G1976), .ZN(n674) );
  XOR2_X1 U740 ( .A(KEYINPUT107), .B(n674), .Z(n956) );
  NAND2_X1 U741 ( .A1(n675), .A2(n956), .ZN(n676) );
  NOR2_X1 U742 ( .A1(n715), .A2(n676), .ZN(n677) );
  NOR2_X1 U743 ( .A1(KEYINPUT33), .A2(n677), .ZN(n680) );
  NAND2_X1 U744 ( .A1(n955), .A2(KEYINPUT33), .ZN(n678) );
  NOR2_X1 U745 ( .A1(n678), .A2(n715), .ZN(n679) );
  NOR2_X1 U746 ( .A1(n680), .A2(n679), .ZN(n708) );
  XOR2_X1 U747 ( .A(G305), .B(G1981), .Z(n952) );
  NAND2_X1 U748 ( .A1(G95), .A2(n868), .ZN(n682) );
  NAND2_X1 U749 ( .A1(G107), .A2(n872), .ZN(n681) );
  NAND2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n688) );
  NAND2_X1 U751 ( .A1(G131), .A2(n511), .ZN(n686) );
  NAND2_X1 U752 ( .A1(G119), .A2(n684), .ZN(n685) );
  NAND2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  OR2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n885) );
  NAND2_X1 U755 ( .A1(G1991), .A2(n885), .ZN(n698) );
  NAND2_X1 U756 ( .A1(G105), .A2(n868), .ZN(n689) );
  XNOR2_X1 U757 ( .A(n689), .B(KEYINPUT38), .ZN(n696) );
  NAND2_X1 U758 ( .A1(G141), .A2(n511), .ZN(n691) );
  NAND2_X1 U759 ( .A1(G129), .A2(n684), .ZN(n690) );
  NAND2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n694) );
  NAND2_X1 U761 ( .A1(n872), .A2(G117), .ZN(n692) );
  XOR2_X1 U762 ( .A(KEYINPUT94), .B(n692), .Z(n693) );
  NOR2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n866) );
  NAND2_X1 U765 ( .A1(G1996), .A2(n866), .ZN(n697) );
  NAND2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n904) );
  INV_X1 U767 ( .A(n699), .ZN(n700) );
  NOR2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n747) );
  XOR2_X1 U769 ( .A(n747), .B(KEYINPUT95), .Z(n702) );
  NAND2_X1 U770 ( .A1(n904), .A2(n702), .ZN(n703) );
  XOR2_X1 U771 ( .A(KEYINPUT96), .B(n703), .Z(n739) );
  XNOR2_X1 U772 ( .A(n739), .B(KEYINPUT97), .ZN(n705) );
  XNOR2_X1 U773 ( .A(G1986), .B(G290), .ZN(n975) );
  NAND2_X1 U774 ( .A1(n975), .A2(n747), .ZN(n704) );
  NAND2_X1 U775 ( .A1(n705), .A2(n704), .ZN(n719) );
  INV_X1 U776 ( .A(n719), .ZN(n706) );
  AND2_X1 U777 ( .A1(n952), .A2(n706), .ZN(n707) );
  NAND2_X1 U778 ( .A1(n708), .A2(n707), .ZN(n721) );
  NOR2_X1 U779 ( .A1(G2090), .A2(G303), .ZN(n709) );
  NAND2_X1 U780 ( .A1(G8), .A2(n709), .ZN(n710) );
  NAND2_X1 U781 ( .A1(n711), .A2(n710), .ZN(n712) );
  AND2_X1 U782 ( .A1(n712), .A2(n715), .ZN(n717) );
  NOR2_X1 U783 ( .A1(G305), .A2(G1981), .ZN(n713) );
  XOR2_X1 U784 ( .A(n713), .B(KEYINPUT24), .Z(n714) );
  NOR2_X1 U785 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n718) );
  OR2_X1 U787 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n735) );
  XNOR2_X1 U789 ( .A(G2067), .B(KEYINPUT37), .ZN(n722) );
  XNOR2_X1 U790 ( .A(n722), .B(KEYINPUT90), .ZN(n744) );
  NAND2_X1 U791 ( .A1(G104), .A2(n868), .ZN(n724) );
  NAND2_X1 U792 ( .A1(G140), .A2(n511), .ZN(n723) );
  NAND2_X1 U793 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U794 ( .A(n725), .B(KEYINPUT34), .ZN(n726) );
  XNOR2_X1 U795 ( .A(n726), .B(KEYINPUT91), .ZN(n732) );
  XNOR2_X1 U796 ( .A(KEYINPUT35), .B(KEYINPUT92), .ZN(n730) );
  NAND2_X1 U797 ( .A1(G116), .A2(n872), .ZN(n728) );
  NAND2_X1 U798 ( .A1(G128), .A2(n684), .ZN(n727) );
  NAND2_X1 U799 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U800 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U801 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U802 ( .A(KEYINPUT36), .B(n733), .Z(n880) );
  NOR2_X1 U803 ( .A1(n744), .A2(n880), .ZN(n906) );
  NAND2_X1 U804 ( .A1(n906), .A2(n747), .ZN(n734) );
  XOR2_X1 U805 ( .A(KEYINPUT93), .B(n734), .Z(n742) );
  NAND2_X1 U806 ( .A1(n735), .A2(n742), .ZN(n736) );
  XNOR2_X1 U807 ( .A(n736), .B(KEYINPUT108), .ZN(n749) );
  NOR2_X1 U808 ( .A1(G1996), .A2(n866), .ZN(n914) );
  NOR2_X1 U809 ( .A1(G1986), .A2(G290), .ZN(n737) );
  NOR2_X1 U810 ( .A1(G1991), .A2(n885), .ZN(n905) );
  NOR2_X1 U811 ( .A1(n737), .A2(n905), .ZN(n738) );
  NOR2_X1 U812 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U813 ( .A1(n914), .A2(n740), .ZN(n741) );
  XNOR2_X1 U814 ( .A(n741), .B(KEYINPUT39), .ZN(n743) );
  NAND2_X1 U815 ( .A1(n743), .A2(n742), .ZN(n745) );
  NAND2_X1 U816 ( .A1(n744), .A2(n880), .ZN(n920) );
  NAND2_X1 U817 ( .A1(n745), .A2(n920), .ZN(n746) );
  NAND2_X1 U818 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U819 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U820 ( .A(n750), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U821 ( .A(G2435), .B(G2454), .Z(n752) );
  XNOR2_X1 U822 ( .A(G2430), .B(G2438), .ZN(n751) );
  XNOR2_X1 U823 ( .A(n752), .B(n751), .ZN(n759) );
  XOR2_X1 U824 ( .A(G2446), .B(KEYINPUT109), .Z(n754) );
  XNOR2_X1 U825 ( .A(G2451), .B(G2443), .ZN(n753) );
  XNOR2_X1 U826 ( .A(n754), .B(n753), .ZN(n755) );
  XOR2_X1 U827 ( .A(n755), .B(G2427), .Z(n757) );
  XNOR2_X1 U828 ( .A(G1341), .B(G1348), .ZN(n756) );
  XNOR2_X1 U829 ( .A(n757), .B(n756), .ZN(n758) );
  XNOR2_X1 U830 ( .A(n759), .B(n758), .ZN(n760) );
  AND2_X1 U831 ( .A1(n760), .A2(G14), .ZN(G401) );
  AND2_X1 U832 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U833 ( .A(G57), .ZN(G237) );
  NAND2_X1 U834 ( .A1(G7), .A2(G661), .ZN(n761) );
  XNOR2_X1 U835 ( .A(n761), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U836 ( .A(G223), .ZN(n824) );
  NAND2_X1 U837 ( .A1(n824), .A2(G567), .ZN(n762) );
  XOR2_X1 U838 ( .A(KEYINPUT11), .B(n762), .Z(G234) );
  INV_X1 U839 ( .A(G860), .ZN(n768) );
  OR2_X1 U840 ( .A1(n966), .A2(n768), .ZN(G153) );
  XNOR2_X1 U841 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U842 ( .A1(G868), .A2(G301), .ZN(n764) );
  OR2_X1 U843 ( .A1(n969), .A2(G868), .ZN(n763) );
  NAND2_X1 U844 ( .A1(n764), .A2(n763), .ZN(G284) );
  XNOR2_X1 U845 ( .A(KEYINPUT75), .B(G868), .ZN(n765) );
  NOR2_X1 U846 ( .A1(G286), .A2(n765), .ZN(n767) );
  NOR2_X1 U847 ( .A1(G868), .A2(G299), .ZN(n766) );
  NOR2_X1 U848 ( .A1(n767), .A2(n766), .ZN(G297) );
  NAND2_X1 U849 ( .A1(n768), .A2(G559), .ZN(n769) );
  NAND2_X1 U850 ( .A1(n769), .A2(n969), .ZN(n770) );
  XNOR2_X1 U851 ( .A(n770), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U852 ( .A1(G868), .A2(n966), .ZN(n773) );
  NAND2_X1 U853 ( .A1(n969), .A2(G868), .ZN(n771) );
  NOR2_X1 U854 ( .A1(G559), .A2(n771), .ZN(n772) );
  NOR2_X1 U855 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U856 ( .A(KEYINPUT76), .B(n774), .ZN(G282) );
  NAND2_X1 U857 ( .A1(G99), .A2(n868), .ZN(n776) );
  NAND2_X1 U858 ( .A1(G111), .A2(n872), .ZN(n775) );
  NAND2_X1 U859 ( .A1(n776), .A2(n775), .ZN(n782) );
  NAND2_X1 U860 ( .A1(G123), .A2(n684), .ZN(n777) );
  XNOR2_X1 U861 ( .A(n777), .B(KEYINPUT18), .ZN(n779) );
  NAND2_X1 U862 ( .A1(G135), .A2(n511), .ZN(n778) );
  NAND2_X1 U863 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U864 ( .A(KEYINPUT77), .B(n780), .Z(n781) );
  NOR2_X1 U865 ( .A1(n782), .A2(n781), .ZN(n923) );
  XNOR2_X1 U866 ( .A(n923), .B(G2096), .ZN(n784) );
  INV_X1 U867 ( .A(G2100), .ZN(n783) );
  NAND2_X1 U868 ( .A1(n784), .A2(n783), .ZN(G156) );
  NAND2_X1 U869 ( .A1(G559), .A2(n969), .ZN(n785) );
  XNOR2_X1 U870 ( .A(n785), .B(n966), .ZN(n804) );
  NOR2_X1 U871 ( .A1(n804), .A2(G860), .ZN(n796) );
  NAND2_X1 U872 ( .A1(G67), .A2(n786), .ZN(n789) );
  NAND2_X1 U873 ( .A1(G55), .A2(n787), .ZN(n788) );
  NAND2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n795) );
  NAND2_X1 U875 ( .A1(G93), .A2(n790), .ZN(n793) );
  NAND2_X1 U876 ( .A1(G80), .A2(n791), .ZN(n792) );
  NAND2_X1 U877 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U878 ( .A1(n795), .A2(n794), .ZN(n799) );
  XNOR2_X1 U879 ( .A(n796), .B(n799), .ZN(G145) );
  NOR2_X1 U880 ( .A1(G868), .A2(n799), .ZN(n797) );
  XOR2_X1 U881 ( .A(n797), .B(KEYINPUT82), .Z(n807) );
  XNOR2_X1 U882 ( .A(KEYINPUT19), .B(G290), .ZN(n798) );
  XNOR2_X1 U883 ( .A(n798), .B(G288), .ZN(n800) );
  XOR2_X1 U884 ( .A(n800), .B(n799), .Z(n802) );
  XNOR2_X1 U885 ( .A(G166), .B(G305), .ZN(n801) );
  XNOR2_X1 U886 ( .A(n802), .B(n801), .ZN(n803) );
  XNOR2_X1 U887 ( .A(n803), .B(G299), .ZN(n894) );
  XNOR2_X1 U888 ( .A(n894), .B(n804), .ZN(n805) );
  NAND2_X1 U889 ( .A1(G868), .A2(n805), .ZN(n806) );
  NAND2_X1 U890 ( .A1(n807), .A2(n806), .ZN(G295) );
  NAND2_X1 U891 ( .A1(G2084), .A2(G2078), .ZN(n808) );
  XNOR2_X1 U892 ( .A(n808), .B(KEYINPUT20), .ZN(n809) );
  XNOR2_X1 U893 ( .A(KEYINPUT83), .B(n809), .ZN(n810) );
  NAND2_X1 U894 ( .A1(n810), .A2(G2090), .ZN(n811) );
  XNOR2_X1 U895 ( .A(KEYINPUT21), .B(n811), .ZN(n812) );
  NAND2_X1 U896 ( .A1(n812), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U897 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U898 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n814) );
  NAND2_X1 U899 ( .A1(G132), .A2(G82), .ZN(n813) );
  XNOR2_X1 U900 ( .A(n814), .B(n813), .ZN(n815) );
  XNOR2_X1 U901 ( .A(n815), .B(KEYINPUT84), .ZN(n816) );
  NOR2_X1 U902 ( .A1(G218), .A2(n816), .ZN(n817) );
  XNOR2_X1 U903 ( .A(KEYINPUT86), .B(n817), .ZN(n818) );
  NAND2_X1 U904 ( .A1(n818), .A2(G96), .ZN(n829) );
  NAND2_X1 U905 ( .A1(n829), .A2(G2106), .ZN(n822) );
  NAND2_X1 U906 ( .A1(G120), .A2(G108), .ZN(n819) );
  NOR2_X1 U907 ( .A1(G237), .A2(n819), .ZN(n820) );
  NAND2_X1 U908 ( .A1(G69), .A2(n820), .ZN(n830) );
  NAND2_X1 U909 ( .A1(n830), .A2(G567), .ZN(n821) );
  NAND2_X1 U910 ( .A1(n822), .A2(n821), .ZN(n831) );
  NAND2_X1 U911 ( .A1(G483), .A2(G661), .ZN(n823) );
  NOR2_X1 U912 ( .A1(n831), .A2(n823), .ZN(n826) );
  NAND2_X1 U913 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n824), .ZN(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U916 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G1), .A2(G3), .ZN(n827) );
  NAND2_X1 U918 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U919 ( .A(n828), .B(KEYINPUT110), .ZN(G188) );
  XNOR2_X1 U920 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U922 ( .A(G132), .ZN(G219) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  INV_X1 U925 ( .A(G82), .ZN(G220) );
  NOR2_X1 U926 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  INV_X1 U928 ( .A(n831), .ZN(G319) );
  XNOR2_X1 U929 ( .A(G1996), .B(G2474), .ZN(n841) );
  XOR2_X1 U930 ( .A(G1981), .B(G1956), .Z(n833) );
  XNOR2_X1 U931 ( .A(G1986), .B(G1991), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U933 ( .A(G1976), .B(G1966), .Z(n835) );
  XNOR2_X1 U934 ( .A(G1971), .B(G1961), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U936 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U937 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(G229) );
  XOR2_X1 U940 ( .A(KEYINPUT111), .B(G2084), .Z(n843) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2090), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U943 ( .A(n844), .B(G2100), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2072), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U946 ( .A(G2096), .B(KEYINPUT43), .Z(n848) );
  XNOR2_X1 U947 ( .A(G2678), .B(KEYINPUT42), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U949 ( .A(n850), .B(n849), .Z(G227) );
  NAND2_X1 U950 ( .A1(G100), .A2(n868), .ZN(n852) );
  NAND2_X1 U951 ( .A1(G112), .A2(n872), .ZN(n851) );
  NAND2_X1 U952 ( .A1(n852), .A2(n851), .ZN(n857) );
  NAND2_X1 U953 ( .A1(n684), .A2(G124), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U955 ( .A1(n511), .A2(G136), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U957 ( .A1(n857), .A2(n856), .ZN(G162) );
  NAND2_X1 U958 ( .A1(G106), .A2(n868), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G142), .A2(n511), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n860), .B(KEYINPUT45), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G118), .A2(n872), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G130), .A2(n684), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U965 ( .A(KEYINPUT113), .B(n863), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n882) );
  NAND2_X1 U968 ( .A1(G103), .A2(n868), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G139), .A2(n511), .ZN(n870) );
  NAND2_X1 U970 ( .A1(n871), .A2(n870), .ZN(n878) );
  NAND2_X1 U971 ( .A1(G115), .A2(n872), .ZN(n874) );
  NAND2_X1 U972 ( .A1(G127), .A2(n684), .ZN(n873) );
  NAND2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U974 ( .A(KEYINPUT114), .B(n875), .Z(n876) );
  XNOR2_X1 U975 ( .A(KEYINPUT47), .B(n876), .ZN(n877) );
  NOR2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n909) );
  XOR2_X1 U977 ( .A(G160), .B(n909), .Z(n879) );
  XNOR2_X1 U978 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n884) );
  XNOR2_X1 U980 ( .A(G162), .B(n923), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n890) );
  XNOR2_X1 U982 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n887) );
  XNOR2_X1 U983 ( .A(n885), .B(KEYINPUT46), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U985 ( .A(G164), .B(n888), .Z(n889) );
  XNOR2_X1 U986 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U987 ( .A1(G37), .A2(n891), .ZN(G395) );
  XNOR2_X1 U988 ( .A(n966), .B(KEYINPUT116), .ZN(n893) );
  XNOR2_X1 U989 ( .A(G171), .B(n969), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n896) );
  XOR2_X1 U991 ( .A(G286), .B(n894), .Z(n895) );
  XNOR2_X1 U992 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U993 ( .A1(G37), .A2(n897), .ZN(G397) );
  NOR2_X1 U994 ( .A1(G229), .A2(G227), .ZN(n898) );
  XNOR2_X1 U995 ( .A(KEYINPUT49), .B(n898), .ZN(n899) );
  NOR2_X1 U996 ( .A1(G401), .A2(n899), .ZN(n900) );
  AND2_X1 U997 ( .A1(G319), .A2(n900), .ZN(n902) );
  NOR2_X1 U998 ( .A1(G395), .A2(G397), .ZN(n901) );
  NAND2_X1 U999 ( .A1(n902), .A2(n901), .ZN(G225) );
  INV_X1 U1000 ( .A(G225), .ZN(G308) );
  INV_X1 U1001 ( .A(G69), .ZN(G235) );
  INV_X1 U1002 ( .A(KEYINPUT55), .ZN(n927) );
  XNOR2_X1 U1003 ( .A(KEYINPUT52), .B(KEYINPUT118), .ZN(n925) );
  XOR2_X1 U1004 ( .A(G160), .B(G2084), .Z(n903) );
  NOR2_X1 U1005 ( .A1(n904), .A2(n903), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(n919) );
  XOR2_X1 U1008 ( .A(G2072), .B(n909), .Z(n911) );
  XOR2_X1 U1009 ( .A(G164), .B(G2078), .Z(n910) );
  NOR2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(KEYINPUT50), .B(n912), .ZN(n917) );
  XOR2_X1 U1012 ( .A(G2090), .B(G162), .Z(n913) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1014 ( .A(KEYINPUT51), .B(n915), .Z(n916) );
  NAND2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n921) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1019 ( .A(n925), .B(n924), .ZN(n926) );
  NAND2_X1 U1020 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1021 ( .A1(n928), .A2(G29), .ZN(n951) );
  XOR2_X1 U1022 ( .A(G2090), .B(G35), .Z(n931) );
  XOR2_X1 U1023 ( .A(G34), .B(KEYINPUT54), .Z(n929) );
  XNOR2_X1 U1024 ( .A(G2084), .B(n929), .ZN(n930) );
  NAND2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n944) );
  XNOR2_X1 U1026 ( .A(G1996), .B(G32), .ZN(n933) );
  XNOR2_X1 U1027 ( .A(G33), .B(G2072), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n938) );
  XOR2_X1 U1029 ( .A(G1991), .B(G25), .Z(n934) );
  NAND2_X1 U1030 ( .A1(n934), .A2(G28), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(G26), .B(G2067), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n941) );
  XOR2_X1 U1034 ( .A(G27), .B(n939), .Z(n940) );
  NOR2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(n942), .B(KEYINPUT53), .ZN(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(KEYINPUT55), .B(n945), .ZN(n946) );
  XNOR2_X1 U1039 ( .A(n946), .B(KEYINPUT119), .ZN(n947) );
  OR2_X1 U1040 ( .A1(G29), .A2(n947), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n948), .A2(G11), .ZN(n949) );
  XOR2_X1 U1042 ( .A(KEYINPUT120), .B(n949), .Z(n950) );
  NAND2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n1009) );
  XNOR2_X1 U1044 ( .A(G16), .B(KEYINPUT56), .ZN(n979) );
  XNOR2_X1 U1045 ( .A(G168), .B(G1966), .ZN(n953) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(n954), .B(KEYINPUT57), .ZN(n965) );
  INV_X1 U1048 ( .A(n955), .ZN(n957) );
  NAND2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(n958), .B(KEYINPUT121), .ZN(n960) );
  NAND2_X1 U1051 ( .A1(G1971), .A2(G303), .ZN(n959) );
  NAND2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1053 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(n963), .B(KEYINPUT122), .ZN(n964) );
  NAND2_X1 U1055 ( .A1(n965), .A2(n964), .ZN(n968) );
  XNOR2_X1 U1056 ( .A(G1341), .B(n966), .ZN(n967) );
  NOR2_X1 U1057 ( .A1(n968), .A2(n967), .ZN(n977) );
  XNOR2_X1 U1058 ( .A(n969), .B(G1348), .ZN(n973) );
  XOR2_X1 U1059 ( .A(G171), .B(G1961), .Z(n971) );
  XNOR2_X1 U1060 ( .A(G299), .B(G1956), .ZN(n970) );
  NOR2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1062 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1063 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1064 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1065 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1066 ( .A(n980), .B(KEYINPUT123), .ZN(n1006) );
  XNOR2_X1 U1067 ( .A(G20), .B(n981), .ZN(n985) );
  XNOR2_X1 U1068 ( .A(G1341), .B(G19), .ZN(n983) );
  XNOR2_X1 U1069 ( .A(G1981), .B(G6), .ZN(n982) );
  NOR2_X1 U1070 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1071 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1072 ( .A(KEYINPUT59), .B(G1348), .Z(n986) );
  XNOR2_X1 U1073 ( .A(G4), .B(n986), .ZN(n987) );
  NOR2_X1 U1074 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1075 ( .A(KEYINPUT60), .B(n989), .Z(n991) );
  XNOR2_X1 U1076 ( .A(G1961), .B(G5), .ZN(n990) );
  NOR2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n1002) );
  XOR2_X1 U1078 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n998) );
  XNOR2_X1 U1079 ( .A(G1971), .B(G22), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(G23), .B(G1976), .ZN(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n996) );
  XOR2_X1 U1082 ( .A(G1986), .B(KEYINPUT124), .Z(n994) );
  XNOR2_X1 U1083 ( .A(G24), .B(n994), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(n998), .B(n997), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(G21), .B(G1966), .ZN(n999) );
  NOR2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(KEYINPUT61), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1090 ( .A1(n1004), .A2(G16), .ZN(n1005) );
  NOR2_X1 U1091 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1092 ( .A(n1007), .B(KEYINPUT126), .Z(n1008) );
  NOR2_X1 U1093 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1094 ( .A(KEYINPUT62), .B(n1010), .Z(n1011) );
  XNOR2_X1 U1095 ( .A(KEYINPUT127), .B(n1011), .ZN(G311) );
  INV_X1 U1096 ( .A(G311), .ZN(G150) );
endmodule

