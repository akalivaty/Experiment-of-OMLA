//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1265, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(new_n203), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G97), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n202), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n210), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n213), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT64), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n221), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n234), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT74), .ZN(new_n247));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  INV_X1    g0048(.A(G45), .ZN(new_n249));
  AOI21_X1  g0049(.A(G1), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n252), .A3(G274), .ZN(new_n253));
  INV_X1    g0053(.A(G226), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n253), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT65), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n253), .B(KEYINPUT65), .C1(new_n254), .C2(new_n256), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G223), .A3(G1698), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G77), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT66), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n265), .A2(new_n272), .A3(G222), .A4(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n265), .A2(G222), .A3(new_n273), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT66), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n271), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n259), .B(new_n260), .C1(new_n277), .C2(new_n252), .ZN(new_n278));
  INV_X1    g0078(.A(G190), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n247), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n276), .A2(new_n274), .ZN(new_n281));
  INV_X1    g0081(.A(new_n271), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n252), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n259), .A2(new_n260), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(KEYINPUT74), .A3(G190), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT9), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n201), .B1(new_n207), .B2(G20), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT69), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT68), .ZN(new_n291));
  INV_X1    g0091(.A(G13), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n292), .A2(new_n208), .A3(G1), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n217), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n291), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n293), .A2(new_n295), .A3(new_n291), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n290), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n292), .A2(G1), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G20), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n299), .B1(G50), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n295), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT8), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G58), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n262), .A2(G20), .ZN(new_n308));
  NOR2_X1   g0108(.A1(G20), .A2(G33), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n307), .A2(new_n308), .B1(G150), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT67), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n310), .A2(new_n311), .B1(G20), .B2(new_n204), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT8), .B(G58), .ZN(new_n313));
  INV_X1    g0113(.A(new_n308), .ZN(new_n314));
  INV_X1    g0114(.A(G150), .ZN(new_n315));
  INV_X1    g0115(.A(new_n309), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n313), .A2(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT67), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n303), .B1(new_n312), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n288), .B1(new_n302), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n298), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n296), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(new_n290), .B1(new_n201), .B2(new_n293), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n204), .A2(G20), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n317), .B2(KEYINPUT67), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n310), .A2(new_n311), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n295), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n323), .A2(KEYINPUT9), .A3(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT73), .B(G200), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n283), .B2(new_n284), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n320), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n287), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT10), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT10), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n287), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n293), .A2(new_n203), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT12), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n309), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n340));
  INV_X1    g0140(.A(G77), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n314), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT11), .A3(new_n295), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n293), .A2(new_n295), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n207), .A2(G20), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(G68), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n339), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT11), .B1(new_n342), .B2(new_n295), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G169), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(KEYINPUT76), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n221), .A2(G1698), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(G226), .B2(G1698), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n354), .B1(new_n356), .B2(new_n269), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n252), .A2(G238), .A3(new_n255), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n253), .A2(new_n360), .A3(KEYINPUT75), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT75), .B1(new_n253), .B2(new_n360), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT13), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n365), .B(new_n359), .C1(new_n361), .C2(new_n362), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n353), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT14), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n364), .A2(G179), .A3(new_n366), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n367), .B2(new_n368), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n350), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n364), .A2(G190), .A3(new_n366), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n349), .ZN(new_n375));
  INV_X1    g0175(.A(G200), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n364), .B2(new_n366), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n307), .A2(new_n309), .B1(G20), .B2(G77), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT71), .ZN(new_n381));
  XNOR2_X1  g0181(.A(KEYINPUT15), .B(G87), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n380), .A2(new_n381), .B1(new_n314), .B2(new_n382), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n313), .A2(new_n316), .B1(new_n208), .B2(new_n341), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(KEYINPUT71), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n295), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT72), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n386), .B(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n265), .A2(G238), .A3(G1698), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n265), .A2(G232), .A3(new_n273), .ZN(new_n390));
  INV_X1    g0190(.A(G107), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n389), .B(new_n390), .C1(new_n391), .C2(new_n265), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n358), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n252), .A2(G244), .A3(new_n255), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n253), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT70), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n396), .B1(new_n393), .B2(new_n395), .ZN(new_n398));
  OAI21_X1  g0198(.A(G190), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n393), .A2(new_n395), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT70), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n330), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n341), .B1(new_n207), .B2(G20), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n344), .A2(new_n404), .B1(new_n341), .B2(new_n293), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n388), .A2(new_n399), .A3(new_n403), .A4(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n382), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n384), .A2(KEYINPUT71), .B1(new_n308), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(KEYINPUT71), .B2(new_n384), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT72), .B1(new_n409), .B2(new_n295), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n386), .A2(new_n387), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n405), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G179), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n397), .B2(new_n398), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n401), .A2(new_n351), .A3(new_n402), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n285), .A2(new_n413), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n278), .A2(new_n351), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n323), .A2(new_n327), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n406), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n337), .A2(new_n373), .A3(new_n379), .A4(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n307), .A2(new_n345), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n322), .A2(new_n423), .B1(new_n293), .B2(new_n313), .ZN(new_n424));
  XNOR2_X1  g0224(.A(G58), .B(G68), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n425), .A2(G20), .B1(G159), .B2(new_n309), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT7), .ZN(new_n427));
  NOR4_X1   g0227(.A1(new_n267), .A2(new_n268), .A3(new_n427), .A4(G20), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT77), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n267), .B2(new_n268), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n263), .A2(KEYINPUT77), .A3(new_n264), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n431), .A3(new_n208), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n428), .B1(new_n432), .B2(new_n427), .ZN(new_n433));
  OAI211_X1 g0233(.A(KEYINPUT16), .B(new_n426), .C1(new_n433), .C2(new_n203), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n295), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n427), .B1(new_n265), .B2(G20), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT78), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n269), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n269), .A2(KEYINPUT78), .A3(KEYINPUT7), .A4(new_n208), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(G68), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT16), .B1(new_n441), .B2(new_n426), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n424), .B1(new_n435), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n254), .A2(G1698), .ZN(new_n444));
  OAI221_X1 g0244(.A(new_n444), .B1(G223), .B2(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G87), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n252), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n253), .B1(new_n221), .B2(new_n256), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G179), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n351), .B2(new_n449), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n443), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT18), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n443), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n449), .A2(new_n376), .ZN(new_n456));
  AND2_X1   g0256(.A1(KEYINPUT79), .A2(G190), .ZN(new_n457));
  NOR2_X1   g0257(.A1(KEYINPUT79), .A2(G190), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n447), .A2(new_n448), .A3(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n461), .B(new_n424), .C1(new_n435), .C2(new_n442), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT17), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n441), .A2(new_n426), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n295), .B(new_n434), .C1(new_n465), .C2(KEYINPUT16), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n466), .A2(KEYINPUT17), .A3(new_n424), .A4(new_n461), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n453), .A2(new_n455), .A3(new_n464), .A4(new_n467), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n468), .A2(KEYINPUT80), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(KEYINPUT80), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n422), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT84), .ZN(new_n472));
  OAI211_X1 g0272(.A(G244), .B(new_n273), .C1(new_n267), .C2(new_n268), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT4), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT83), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT83), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n473), .A2(new_n477), .A3(new_n474), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n265), .A2(KEYINPUT4), .A3(G244), .A4(new_n273), .ZN(new_n479));
  OAI211_X1 g0279(.A(G250), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n476), .A2(new_n478), .A3(new_n479), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n358), .ZN(new_n484));
  AND2_X1   g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  NOR2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n249), .A2(G1), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n487), .A2(G274), .A3(new_n252), .A4(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n485), .B2(new_n486), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n252), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n491), .B2(new_n223), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n472), .B1(new_n484), .B2(new_n493), .ZN(new_n494));
  AOI211_X1 g0294(.A(KEYINPUT84), .B(new_n492), .C1(new_n483), .C2(new_n358), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n351), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n439), .A2(G107), .A3(new_n440), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n309), .A2(G77), .ZN(new_n498));
  XNOR2_X1  g0298(.A(new_n498), .B(KEYINPUT81), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n391), .A2(KEYINPUT6), .A3(G97), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n222), .A2(new_n391), .ZN(new_n501));
  NOR2_X1   g0301(.A1(G97), .A2(G107), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n500), .B1(new_n503), .B2(KEYINPUT6), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n499), .B1(G20), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n303), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n303), .B(new_n301), .C1(G1), .C2(new_n262), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT82), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n301), .B2(G97), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n293), .A2(KEYINPUT82), .A3(new_n222), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n509), .A2(G97), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n492), .B1(new_n483), .B2(new_n358), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n507), .A2(new_n513), .B1(new_n514), .B2(new_n413), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n496), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n481), .B(new_n480), .C1(new_n473), .C2(new_n474), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n477), .B1(new_n473), .B2(new_n474), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n252), .B1(new_n519), .B2(new_n478), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT84), .B1(new_n520), .B2(new_n492), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n484), .A2(new_n472), .A3(new_n493), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(G190), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n513), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n506), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n514), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G200), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n523), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n252), .A2(G274), .A3(new_n488), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n207), .A2(G45), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n252), .A2(G250), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(G238), .B(new_n273), .C1(new_n267), .C2(new_n268), .ZN(new_n533));
  OAI211_X1 g0333(.A(G244), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G116), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n532), .B1(new_n536), .B2(new_n358), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(G169), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n413), .B2(new_n537), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n407), .A2(new_n301), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n265), .A2(new_n208), .A3(G68), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT85), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT85), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n265), .A2(new_n543), .A3(new_n208), .A4(G68), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n308), .A2(new_n545), .A3(G97), .ZN(new_n546));
  INV_X1    g0346(.A(G87), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n502), .A2(new_n547), .B1(new_n354), .B2(new_n208), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n548), .B2(new_n545), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n542), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n540), .B1(new_n550), .B2(new_n295), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n508), .B2(new_n382), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n537), .A2(new_n329), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n536), .A2(new_n358), .ZN(new_n554));
  INV_X1    g0354(.A(new_n532), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n554), .A2(G190), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n508), .A2(new_n547), .ZN(new_n558));
  AOI211_X1 g0358(.A(new_n540), .B(new_n558), .C1(new_n550), .C2(new_n295), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n539), .A2(new_n552), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n516), .A2(new_n528), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT23), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n208), .B2(G107), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n391), .A2(KEYINPUT23), .A3(G20), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT87), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n535), .B2(G20), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n208), .A2(KEYINPUT87), .A3(G33), .A4(G116), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n208), .B(G87), .C1(new_n267), .C2(new_n268), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n570), .A2(KEYINPUT22), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n570), .A2(KEYINPUT22), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT24), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT24), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n569), .B(new_n575), .C1(new_n571), .C2(new_n572), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n295), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT25), .B1(new_n293), .B2(new_n391), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n293), .A2(KEYINPUT25), .A3(new_n391), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n509), .A2(G107), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  OR2_X1    g0383(.A1(G250), .A2(G1698), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n223), .A2(G1698), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n584), .B(new_n585), .C1(new_n267), .C2(new_n268), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT88), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G294), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n587), .B1(new_n586), .B2(new_n588), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n589), .A2(new_n590), .A3(new_n252), .ZN(new_n591));
  INV_X1    g0391(.A(G264), .ZN(new_n592));
  OAI21_X1  g0392(.A(KEYINPUT89), .B1(new_n491), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT89), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n490), .A2(new_n594), .A3(G264), .A4(new_n252), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT90), .B1(new_n591), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n586), .A2(new_n588), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT88), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n358), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT90), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(new_n593), .A4(new_n595), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n597), .A2(new_n489), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n376), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n601), .A2(new_n489), .A3(new_n593), .A4(new_n595), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(G190), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n583), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT21), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n481), .B(new_n208), .C1(G33), .C2(new_n222), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n611), .B(new_n295), .C1(new_n208), .C2(G116), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n612), .B(KEYINPUT20), .ZN(new_n613));
  INV_X1    g0413(.A(G116), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n293), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n508), .B2(new_n614), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(G303), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n252), .B1(new_n269), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(G257), .A2(G1698), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n273), .A2(G264), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n265), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n490), .A2(G270), .A3(new_n252), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n489), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G169), .ZN(new_n626));
  OAI211_X1 g0426(.A(KEYINPUT86), .B(new_n610), .C1(new_n617), .C2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n623), .A2(G179), .A3(new_n489), .A4(new_n624), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n617), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n625), .A2(G200), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n617), .B(new_n630), .C1(new_n625), .C2(new_n459), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n625), .A2(G169), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n610), .A2(KEYINPUT86), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n632), .B(new_n633), .C1(new_n613), .C2(new_n616), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n627), .A2(new_n629), .A3(new_n631), .A4(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n597), .A2(new_n603), .A3(G179), .A4(new_n489), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n606), .A2(G169), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n636), .A2(new_n637), .B1(new_n578), .B2(new_n582), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n609), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n471), .A2(new_n561), .A3(new_n639), .ZN(G372));
  INV_X1    g0440(.A(new_n420), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT91), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n287), .A2(new_n332), .A3(new_n335), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n335), .B1(new_n287), .B2(new_n332), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n334), .A2(KEYINPUT91), .A3(new_n336), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n453), .A2(new_n455), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n373), .A2(new_n416), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n379), .A2(new_n464), .A3(new_n467), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n641), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n471), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n539), .A2(new_n552), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n516), .A2(new_n528), .A3(new_n560), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n627), .A2(new_n629), .A3(new_n634), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n607), .B1(new_n604), .B2(new_n376), .ZN(new_n657));
  OAI22_X1  g0457(.A1(new_n638), .A2(new_n656), .B1(new_n657), .B2(new_n583), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n654), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n478), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n660), .A2(new_n517), .A3(new_n518), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n413), .B(new_n493), .C1(new_n661), .C2(new_n252), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n506), .B2(new_n524), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n521), .A2(new_n522), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n351), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT26), .B1(new_n665), .B2(new_n560), .ZN(new_n666));
  AND4_X1   g0466(.A1(KEYINPUT26), .A2(new_n560), .A3(new_n496), .A4(new_n515), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n659), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n652), .B1(new_n653), .B2(new_n670), .ZN(G369));
  NOR2_X1   g0471(.A1(new_n609), .A2(new_n638), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n300), .A2(new_n208), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(G213), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n583), .A2(new_n678), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n672), .A2(new_n679), .B1(new_n638), .B2(new_n678), .ZN(new_n680));
  INV_X1    g0480(.A(new_n678), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n617), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n656), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n635), .B2(new_n682), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n656), .A2(new_n681), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n672), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n638), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n689), .B2(new_n678), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n686), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n211), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n502), .A2(new_n547), .A3(new_n614), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n694), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n697), .A2(KEYINPUT92), .B1(new_n215), .B2(new_n694), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(KEYINPUT92), .B2(new_n697), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n669), .B2(new_n681), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n701), .B(new_n681), .C1(new_n659), .C2(new_n668), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n554), .A2(new_n555), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n628), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n597), .A2(new_n603), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n706), .B1(new_n664), .B2(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n597), .A2(new_n708), .A3(new_n603), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(KEYINPUT30), .A3(new_n521), .A4(new_n522), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n707), .A2(new_n413), .A3(new_n625), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT93), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n604), .B(new_n526), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n710), .A2(new_n712), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n678), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n639), .A2(new_n561), .A3(new_n681), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n705), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n700), .B1(new_n727), .B2(G1), .ZN(G364));
  NOR2_X1   g0528(.A1(new_n292), .A2(G20), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n207), .B1(new_n729), .B2(G45), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n693), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n217), .B1(G20), .B2(new_n351), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n692), .A2(new_n269), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G355), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(G116), .B2(new_n211), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n430), .A2(new_n431), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n692), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(new_n249), .B2(new_n216), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n242), .A2(new_n249), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n741), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G179), .A2(G200), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(G20), .A3(new_n279), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n265), .B1(new_n750), .B2(G329), .ZN(new_n751));
  INV_X1    g0551(.A(G322), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n208), .A2(new_n413), .A3(G200), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(new_n458), .B2(new_n457), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n751), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n208), .A2(new_n413), .A3(new_n376), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n459), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(G190), .ZN(new_n759));
  AND2_X1   g0559(.A1(KEYINPUT33), .A2(G317), .ZN(new_n760));
  NOR2_X1   g0560(.A1(KEYINPUT33), .A2(G317), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G326), .A2(new_n758), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G294), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n208), .B1(new_n748), .B2(G190), .ZN(new_n765));
  INV_X1    g0565(.A(G311), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n753), .A2(new_n279), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n763), .B1(new_n764), .B2(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NOR4_X1   g0568(.A1(new_n329), .A2(new_n208), .A3(G179), .A4(new_n279), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n755), .B(new_n768), .C1(G303), .C2(new_n769), .ZN(new_n770));
  NOR4_X1   g0570(.A1(new_n329), .A2(new_n208), .A3(G179), .A4(G190), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT96), .Z(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G283), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(G107), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n767), .A2(KEYINPUT95), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n767), .A2(KEYINPUT95), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n765), .B(KEYINPUT97), .Z(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n778), .A2(new_n341), .B1(new_n780), .B2(new_n222), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n750), .A2(G159), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n759), .A2(G68), .B1(new_n782), .B2(KEYINPUT32), .ZN(new_n783));
  INV_X1    g0583(.A(new_n758), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n783), .B1(new_n201), .B2(new_n784), .C1(new_n202), .C2(new_n754), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n769), .A2(G87), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n786), .B(new_n265), .C1(KEYINPUT32), .C2(new_n782), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n781), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n770), .A2(new_n773), .B1(new_n774), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n736), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n732), .B1(new_n738), .B2(new_n747), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT98), .ZN(new_n792));
  INV_X1    g0592(.A(new_n735), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n684), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n684), .A2(G330), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT94), .Z(new_n796));
  INV_X1    g0596(.A(new_n732), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n796), .A2(new_n685), .A3(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  NOR2_X1   g0600(.A1(new_n736), .A2(new_n733), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n732), .B1(G77), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n269), .B1(new_n749), .B2(new_n766), .ZN(new_n804));
  INV_X1    g0604(.A(new_n759), .ZN(new_n805));
  INV_X1    g0605(.A(G283), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n805), .A2(new_n806), .B1(new_n764), .B2(new_n754), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n804), .B(new_n807), .C1(G303), .C2(new_n758), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n772), .A2(G87), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n769), .A2(G107), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n777), .A2(G116), .B1(new_n779), .B2(G97), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G137), .A2(new_n758), .B1(new_n759), .B2(G150), .ZN(new_n813));
  INV_X1    g0613(.A(G143), .ZN(new_n814));
  INV_X1    g0614(.A(G159), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n813), .B1(new_n814), .B2(new_n754), .C1(new_n778), .C2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n772), .A2(G68), .ZN(new_n819));
  INV_X1    g0619(.A(G132), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n742), .B1(new_n202), .B2(new_n765), .C1(new_n820), .C2(new_n749), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G50), .B2(new_n769), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n818), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n816), .A2(new_n817), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n812), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n803), .B1(new_n825), .B2(new_n736), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n416), .A2(new_n678), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n412), .A2(new_n678), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n406), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n827), .B1(new_n416), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n826), .B1(new_n830), .B2(new_n734), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n669), .A2(new_n681), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n829), .A2(new_n416), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n416), .A2(new_n678), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n681), .B(new_n830), .C1(new_n659), .C2(new_n668), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n836), .A2(KEYINPUT99), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT99), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n832), .A2(new_n839), .A3(new_n835), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n838), .A2(new_n725), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n797), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n725), .B1(new_n838), .B2(new_n840), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n831), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT100), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT100), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n846), .B(new_n831), .C1(new_n842), .C2(new_n843), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(new_n847), .ZN(G384));
  OR2_X1    g0648(.A1(new_n504), .A2(KEYINPUT35), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n504), .A2(KEYINPUT35), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n849), .A2(G116), .A3(new_n218), .A4(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT36), .Z(new_n852));
  OAI211_X1 g0652(.A(new_n216), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n201), .A2(G68), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n207), .B(G13), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n426), .B1(new_n433), .B2(new_n203), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT16), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n424), .B1(new_n859), .B2(new_n435), .ZN(new_n860));
  INV_X1    g0660(.A(new_n676), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n462), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n860), .A2(new_n451), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT37), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n443), .A2(KEYINPUT101), .A3(new_n861), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT101), .B1(new_n443), .B2(new_n861), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n452), .B(new_n462), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n865), .B1(new_n868), .B2(KEYINPUT37), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n468), .A2(new_n861), .A3(new_n860), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n866), .A2(new_n867), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n468), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT104), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n468), .A2(KEYINPUT104), .A3(new_n872), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n443), .A2(new_n861), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT101), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n443), .A2(KEYINPUT101), .A3(new_n861), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT103), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n452), .A2(new_n462), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n882), .A2(new_n883), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n877), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n452), .A2(new_n462), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n880), .B2(new_n881), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n883), .B1(new_n889), .B2(new_n884), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n875), .B(new_n876), .C1(new_n887), .C2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n871), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT39), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n870), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT102), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT102), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n869), .A2(new_n898), .A3(KEYINPUT38), .A4(new_n870), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n869), .A2(new_n870), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n892), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n897), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT39), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n895), .A2(new_n903), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n367), .A2(new_n368), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(new_n369), .A3(new_n371), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(new_n350), .A3(new_n681), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n373), .B(new_n379), .C1(new_n349), .C2(new_n681), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n350), .B(new_n678), .C1(new_n906), .C2(new_n378), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n837), .A2(new_n834), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n902), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n648), .A2(new_n861), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n909), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n471), .B1(new_n702), .B2(new_n704), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n652), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(KEYINPUT105), .A2(KEYINPUT31), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n718), .A2(new_n678), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n718), .B2(new_n678), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n722), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n835), .B1(new_n910), .B2(new_n911), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT40), .B1(new_n893), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(KEYINPUT40), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n902), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n471), .A3(new_n923), .ZN(new_n930));
  INV_X1    g0730(.A(new_n925), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n468), .A2(KEYINPUT104), .A3(new_n872), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT104), .B1(new_n468), .B2(new_n872), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT103), .B1(new_n868), .B2(KEYINPUT37), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(new_n877), .A3(new_n886), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT38), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n931), .B1(new_n937), .B2(new_n871), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n938), .A2(KEYINPUT40), .B1(new_n902), .B2(new_n927), .ZN(new_n939));
  INV_X1    g0739(.A(new_n923), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n939), .B1(new_n653), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n930), .A2(new_n941), .A3(G330), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n919), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n207), .B2(new_n729), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n919), .A2(new_n942), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n856), .B1(new_n944), .B2(new_n945), .ZN(G367));
  NAND2_X1  g0746(.A1(new_n234), .A2(new_n743), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n947), .B(new_n737), .C1(new_n211), .C2(new_n382), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n732), .B1(new_n949), .B2(KEYINPUT109), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(KEYINPUT109), .B2(new_n949), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n654), .A2(new_n559), .A3(new_n681), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n560), .B1(new_n559), .B2(new_n681), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n742), .ZN(new_n955));
  INV_X1    g0755(.A(G317), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n955), .B1(new_n956), .B2(new_n749), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n805), .A2(new_n764), .B1(new_n391), .B2(new_n765), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n957), .B(new_n958), .C1(G97), .C2(new_n771), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n769), .A2(KEYINPUT46), .A3(G116), .ZN(new_n960));
  INV_X1    g0760(.A(new_n754), .ZN(new_n961));
  AOI22_X1  g0761(.A1(G311), .A2(new_n758), .B1(new_n961), .B2(G303), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(KEYINPUT110), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(G283), .B2(new_n777), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT46), .B1(new_n769), .B2(G116), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(new_n962), .B2(KEYINPUT110), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n959), .A2(new_n960), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n777), .A2(G50), .B1(G159), .B2(new_n759), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(KEYINPUT111), .ZN(new_n970));
  INV_X1    g0770(.A(G137), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n265), .B1(new_n971), .B2(new_n749), .C1(new_n784), .C2(new_n814), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(G150), .B2(new_n961), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n779), .A2(G68), .ZN(new_n974));
  AOI22_X1  g0774(.A1(G58), .A2(new_n769), .B1(new_n771), .B2(G77), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n970), .A2(new_n973), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n969), .A2(KEYINPUT111), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n967), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT47), .Z(new_n979));
  OAI221_X1 g0779(.A(new_n951), .B1(new_n793), .B2(new_n954), .C1(new_n979), .C2(new_n790), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n516), .B(new_n528), .C1(new_n525), .C2(new_n681), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n665), .A2(new_n678), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT106), .Z(new_n984));
  OAI21_X1  g0784(.A(new_n516), .B1(new_n984), .B2(new_n689), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n681), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n983), .A2(new_n688), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT42), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n986), .A2(new_n988), .B1(KEYINPUT43), .B2(new_n954), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n989), .A2(new_n991), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n686), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n984), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n994), .B(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n690), .A2(new_n983), .ZN(new_n999));
  XOR2_X1   g0799(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n690), .A2(new_n983), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT44), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(new_n686), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n687), .ZN(new_n1007));
  AOI21_X1  g0807(.A(KEYINPUT108), .B1(new_n680), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n672), .B2(new_n687), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n688), .A2(KEYINPUT108), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n685), .ZN(new_n1012));
  OAI211_X1 g0812(.A(G330), .B(new_n684), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n727), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n727), .B1(new_n1006), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n693), .B(KEYINPUT41), .Z(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n731), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n980), .B1(new_n998), .B2(new_n1019), .ZN(G387));
  OR3_X1    g0820(.A1(new_n1014), .A2(new_n727), .A3(KEYINPUT114), .ZN(new_n1021));
  OAI21_X1  g0821(.A(KEYINPUT114), .B1(new_n1014), .B2(new_n727), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1021), .A2(new_n693), .A3(new_n1015), .A4(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n739), .A2(new_n695), .B1(new_n391), .B2(new_n692), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n238), .A2(new_n249), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n307), .A2(new_n201), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n696), .B(new_n249), .C1(new_n203), .C2(new_n341), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n743), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1024), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n797), .B1(new_n1031), .B2(new_n737), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT113), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n784), .B2(new_n815), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n758), .A2(KEYINPUT113), .A3(G159), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n955), .B1(G150), .B2(new_n750), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n769), .A2(G77), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n767), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n961), .A2(G50), .B1(new_n1039), .B2(G68), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n313), .B2(new_n805), .C1(new_n780), .C2(new_n382), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1038), .B(new_n1041), .C1(G97), .C2(new_n772), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n771), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1043), .A2(new_n614), .ZN(new_n1044));
  INV_X1    g0844(.A(G326), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n955), .B1(new_n1045), .B2(new_n749), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G311), .A2(new_n759), .B1(new_n961), .B2(G317), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n752), .B2(new_n784), .C1(new_n778), .C2(new_n618), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n769), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n1052), .A2(new_n764), .B1(new_n806), .B2(new_n765), .ZN(new_n1053));
  OR3_X1    g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1044), .B(new_n1046), .C1(new_n1055), .C2(KEYINPUT49), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(KEYINPUT49), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1042), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1032), .B1(new_n1058), .B2(new_n790), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n680), .B2(new_n735), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n1014), .B2(new_n731), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1023), .A2(new_n1061), .ZN(G393));
  INV_X1    g0862(.A(new_n1015), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n694), .B1(new_n1005), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n1005), .B2(new_n1063), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1005), .A2(new_n731), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n984), .A2(new_n735), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n269), .B1(new_n749), .B2(new_n752), .C1(new_n614), .C2(new_n765), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n805), .A2(new_n618), .B1(new_n767), .B2(new_n764), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(G283), .C2(new_n769), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n784), .A2(new_n956), .B1(new_n766), .B2(new_n754), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT52), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1070), .A2(new_n774), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n955), .B1(G143), .B2(new_n750), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n809), .B(new_n1074), .C1(new_n203), .C2(new_n1052), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT115), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n777), .A2(new_n307), .B1(G50), .B2(new_n759), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(KEYINPUT116), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(KEYINPUT116), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n784), .A2(new_n315), .B1(new_n815), .B2(new_n754), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT51), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1081), .A2(new_n1082), .B1(G77), .B2(new_n779), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1079), .A2(new_n1080), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1073), .B1(new_n1076), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n736), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n737), .B1(new_n222), .B2(new_n211), .C1(new_n744), .C2(new_n245), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1067), .A2(new_n732), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1065), .A2(new_n1066), .A3(new_n1089), .ZN(G390));
  INV_X1    g0890(.A(KEYINPUT123), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n895), .A2(new_n903), .A3(new_n733), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n732), .B1(new_n307), .B2(new_n802), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT122), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n269), .B1(new_n749), .B2(new_n764), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n391), .A2(new_n805), .B1(new_n784), .B2(new_n806), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(G116), .C2(new_n961), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n777), .A2(G97), .B1(new_n779), .B2(G77), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1097), .A2(new_n786), .A3(new_n819), .A4(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n754), .A2(new_n820), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n269), .B1(new_n750), .B2(G125), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n805), .B2(new_n971), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1100), .B(new_n1102), .C1(G128), .C2(new_n758), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(KEYINPUT54), .B(G143), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n777), .A2(new_n1105), .B1(new_n779), .B2(G159), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1103), .B(new_n1106), .C1(new_n201), .C2(new_n1043), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n769), .A2(G150), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT53), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1099), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1094), .B1(new_n1110), .B2(new_n736), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1092), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n913), .A2(new_n912), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n907), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n895), .A2(new_n903), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n724), .A2(new_n924), .A3(G330), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT118), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n724), .A2(new_n924), .A3(KEYINPUT118), .A4(G330), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n913), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT117), .ZN(new_n1122));
  AOI21_X1  g0922(.A(KEYINPUT117), .B1(new_n910), .B2(new_n911), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n907), .B1(new_n937), .B2(new_n871), .C1(new_n1121), .C2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1115), .A2(new_n1120), .A3(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1115), .A2(new_n1125), .ZN(new_n1127));
  INV_X1    g0927(.A(G330), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n940), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n924), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1126), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1091), .B(new_n1112), .C1(new_n1131), .C2(new_n730), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1115), .A2(new_n1120), .A3(new_n1125), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1130), .B1(new_n1115), .B2(new_n1125), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n1133), .A2(new_n1134), .A3(new_n730), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1112), .ZN(new_n1136));
  OAI21_X1  g0936(.A(KEYINPUT123), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n910), .B(new_n911), .C1(new_n725), .C2(new_n835), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1121), .B1(new_n1130), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n923), .A2(G330), .A3(new_n830), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1124), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT120), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1140), .A2(new_n1124), .A3(KEYINPUT120), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1120), .A2(new_n1143), .A3(new_n1121), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT121), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1140), .A2(new_n1124), .A3(KEYINPUT120), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT120), .B1(new_n1140), .B2(new_n1124), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n913), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1150), .A2(KEYINPUT121), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1139), .B1(new_n1147), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1129), .A2(new_n471), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n917), .A2(new_n652), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT119), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT119), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n917), .A2(new_n1154), .A3(new_n1157), .A4(new_n652), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1153), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n693), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1139), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1164));
  AOI21_X1  g0964(.A(KEYINPUT121), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1159), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(new_n1131), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1132), .B(new_n1137), .C1(new_n1162), .C2(new_n1169), .ZN(G378));
  INV_X1    g0970(.A(KEYINPUT57), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n914), .A2(new_n915), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n908), .B2(new_n904), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n645), .A2(new_n646), .A3(new_n420), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n419), .A2(new_n861), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n645), .A2(new_n646), .A3(new_n420), .A4(new_n1175), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1179), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n939), .B2(new_n1128), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1182), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT40), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n887), .A2(new_n890), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n875), .A2(new_n876), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n892), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n896), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1185), .B1(new_n1189), .B2(new_n931), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n928), .ZN(new_n1191));
  OAI211_X1 g0991(.A(G330), .B(new_n1184), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1173), .A2(new_n1183), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1173), .B1(new_n1183), .B2(new_n1192), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1159), .B1(new_n1161), .B2(new_n1166), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1171), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1183), .A2(new_n1192), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT125), .B1(new_n1198), .B2(new_n916), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1184), .B1(new_n929), .B2(G330), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1128), .B(new_n1182), .C1(new_n926), .C2(new_n928), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n916), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1173), .A2(new_n1183), .A3(new_n1192), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1199), .B1(new_n1204), .B2(KEYINPUT125), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1167), .B1(new_n1131), .B2(new_n1153), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT57), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1197), .B(new_n693), .C1(new_n1205), .C2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1182), .A2(new_n733), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n955), .A2(new_n248), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1037), .B1(new_n806), .B2(new_n749), .C1(new_n805), .C2(new_n222), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(G58), .C2(new_n771), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n758), .A2(G116), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n961), .A2(G107), .B1(new_n1039), .B2(new_n407), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1212), .A2(new_n974), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  AOI21_X1  g1016(.A(G50), .B1(new_n262), .B2(new_n248), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1215), .A2(new_n1216), .B1(new_n1210), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1216), .B2(new_n1215), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G132), .A2(new_n759), .B1(new_n961), .B2(G128), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n758), .A2(G125), .B1(new_n1039), .B2(G137), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n315), .B2(new_n780), .C1(new_n1052), .C2(new_n1104), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n771), .A2(G159), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G33), .B(G41), .C1(new_n750), .C2(G124), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n736), .B1(new_n1219), .B2(new_n1229), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT124), .Z(new_n1231));
  AOI21_X1  g1031(.A(new_n797), .B1(new_n201), .B2(new_n801), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1209), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1204), .B2(new_n731), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1208), .A2(new_n1235), .ZN(G375));
  NAND2_X1  g1036(.A1(new_n1153), .A2(new_n1159), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1168), .A2(new_n1018), .A3(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n758), .A2(G132), .B1(new_n1039), .B2(G150), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n971), .B2(new_n754), .C1(new_n805), .C2(new_n1104), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n955), .B1(G128), .B2(new_n750), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n1043), .B2(new_n202), .C1(new_n815), .C2(new_n1052), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1240), .B(new_n1242), .C1(G50), .C2(new_n779), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n778), .A2(new_n391), .B1(new_n780), .B2(new_n382), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1052), .A2(new_n222), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n269), .B1(new_n618), .B2(new_n749), .C1(new_n784), .C2(new_n764), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n805), .A2(new_n614), .B1(new_n806), .B2(new_n754), .ZN(new_n1247));
  NOR4_X1   g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n772), .A2(G77), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1243), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n732), .B1(G68), .B2(new_n802), .C1(new_n1250), .C2(new_n790), .ZN(new_n1251));
  XOR2_X1   g1051(.A(new_n1251), .B(KEYINPUT126), .Z(new_n1252));
  NAND2_X1  g1052(.A1(new_n1124), .A2(new_n733), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1153), .B2(new_n730), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1238), .A2(new_n1257), .ZN(G381));
  NAND3_X1  g1058(.A1(new_n1023), .A2(new_n799), .A3(new_n1061), .ZN(new_n1259));
  OR2_X1    g1059(.A1(G390), .A2(new_n1259), .ZN(new_n1260));
  NOR4_X1   g1060(.A1(new_n1260), .A2(G387), .A3(G384), .A4(G381), .ZN(new_n1261));
  INV_X1    g1061(.A(G378), .ZN(new_n1262));
  INV_X1    g1062(.A(G375), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(G407));
  NAND2_X1  g1064(.A1(new_n677), .A2(G213), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n1262), .A3(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G407), .A2(G213), .A3(new_n1267), .ZN(G409));
  NAND2_X1  g1068(.A1(new_n1266), .A2(G2897), .ZN(new_n1269));
  INV_X1    g1069(.A(G384), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1147), .A2(new_n1152), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1271), .A2(KEYINPUT60), .A3(new_n1159), .A4(new_n1163), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1272), .A2(new_n693), .ZN(new_n1273));
  OAI21_X1  g1073(.A(KEYINPUT60), .B1(new_n1153), .B2(new_n1159), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1237), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1270), .B1(new_n1276), .B2(new_n1257), .ZN(new_n1277));
  AOI211_X1 g1077(.A(G384), .B(new_n1256), .C1(new_n1273), .C2(new_n1275), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1269), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1272), .A2(new_n693), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1237), .B2(new_n1274), .ZN(new_n1281));
  OAI21_X1  g1081(.A(G384), .B1(new_n1281), .B2(new_n1256), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1276), .A2(new_n1270), .A3(new_n1257), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1269), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1279), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1197), .A2(new_n693), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G378), .B(new_n1235), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1290));
  OR2_X1    g1090(.A1(new_n1162), .A2(new_n1169), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1137), .A2(new_n1132), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1205), .A2(new_n730), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1206), .A2(new_n1204), .A3(new_n1018), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1233), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1291), .B(new_n1292), .C1(new_n1293), .C2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1290), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1265), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1287), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT63), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1300), .B1(new_n1298), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(G390), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G387), .A2(new_n1303), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n980), .B(G390), .C1(new_n998), .C2(new_n1019), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G393), .A2(G396), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT127), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(new_n1308), .A3(new_n1259), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1308), .B1(new_n1307), .B2(new_n1259), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1306), .B(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1266), .B1(new_n1290), .B2(new_n1296), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1301), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(KEYINPUT63), .A3(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1299), .A2(new_n1302), .A3(new_n1313), .A4(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1314), .A2(new_n1318), .A3(new_n1315), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT61), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1320), .B1(new_n1314), .B2(new_n1286), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1318), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1319), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1317), .B1(new_n1323), .B2(new_n1313), .ZN(G405));
  NAND2_X1  g1124(.A1(G375), .A2(new_n1262), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1290), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1315), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1325), .A2(new_n1301), .A3(new_n1290), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1330));
  XNOR2_X1  g1130(.A(new_n1306), .B(new_n1330), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1329), .B(new_n1331), .ZN(G402));
endmodule


