//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n599, new_n600, new_n601, new_n603,
    new_n604, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT71), .B(KEYINPUT22), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n210), .A2(KEYINPUT65), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(KEYINPUT65), .ZN(new_n212));
  NOR2_X1   g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  AND2_X1   g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(KEYINPUT24), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  OR2_X1    g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n221), .A2(new_n222), .B1(new_n220), .B2(new_n219), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n217), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT25), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT27), .B(G183gat), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT28), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n219), .A2(KEYINPUT26), .ZN(new_n233));
  INV_X1    g032(.A(new_n218), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n219), .B1(new_n234), .B2(KEYINPUT26), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n214), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  AOI211_X1 g035(.A(KEYINPUT25), .B(new_n221), .C1(new_n220), .C2(new_n219), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n215), .B1(KEYINPUT24), .B2(new_n214), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n232), .A2(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n227), .A2(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(G226gat), .A2(G233gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT29), .B1(new_n227), .B2(new_n239), .ZN(new_n244));
  OAI22_X1  g043(.A1(new_n243), .A2(KEYINPUT72), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT72), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n209), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n244), .A2(new_n241), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n249), .A2(new_n243), .A3(new_n209), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G8gat), .B(G36gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(G64gat), .B(G92gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n252), .A2(KEYINPUT73), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT73), .B1(new_n252), .B2(new_n255), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT30), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n249), .B1(new_n246), .B2(new_n242), .ZN(new_n259));
  INV_X1    g058(.A(new_n247), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n250), .B1(new_n261), .B2(new_n209), .ZN(new_n262));
  INV_X1    g061(.A(new_n255), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n258), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AND4_X1   g063(.A1(new_n258), .A2(new_n248), .A3(new_n251), .A4(new_n263), .ZN(new_n265));
  OAI22_X1  g064(.A1(new_n256), .A2(new_n257), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(new_n209), .B2(KEYINPUT29), .ZN(new_n269));
  NAND2_X1  g068(.A1(G155gat), .A2(G162gat), .ZN(new_n270));
  INV_X1    g069(.A(G155gat), .ZN(new_n271));
  INV_X1    g070(.A(G162gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G141gat), .B(G148gat), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n270), .B(new_n273), .C1(new_n274), .C2(KEYINPUT2), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n270), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT75), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT75), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n273), .A2(new_n278), .A3(new_n270), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n270), .A2(KEYINPUT2), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G148gat), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n282), .A2(G141gat), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT74), .B(G141gat), .Z(new_n284));
  AOI21_X1  g083(.A(new_n283), .B1(new_n284), .B2(G148gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n275), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n268), .B(new_n275), .C1(new_n281), .C2(new_n285), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n209), .B1(new_n289), .B2(KEYINPUT29), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G228gat), .ZN(new_n292));
  INV_X1    g091(.A(G233gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G22gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n287), .A2(new_n294), .A3(new_n290), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n299), .A2(KEYINPUT83), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(KEYINPUT83), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n296), .A2(new_n298), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G22gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G78gat), .B(G106gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(G50gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n297), .A2(KEYINPUT84), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n308), .B1(new_n302), .B2(new_n310), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G15gat), .B(G43gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(KEYINPUT69), .ZN(new_n316));
  XOR2_X1   g115(.A(G71gat), .B(G99gat), .Z(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G127gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G134gat), .ZN(new_n320));
  INV_X1    g119(.A(G134gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G127gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT67), .ZN(new_n323));
  OR3_X1    g122(.A1(new_n321), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(G113gat), .B(G120gat), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n323), .B(new_n324), .C1(KEYINPUT1), .C2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT68), .ZN(new_n327));
  INV_X1    g126(.A(G113gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n328), .A3(G120gat), .ZN(new_n329));
  INV_X1    g128(.A(G120gat), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT68), .B1(new_n330), .B2(G113gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(G113gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n320), .A2(new_n322), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n326), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n240), .B(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G227gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(new_n293), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT33), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n318), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(KEYINPUT32), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n341), .B(KEYINPUT32), .C1(new_n342), .C2(new_n318), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n240), .B(new_n337), .Z(new_n348));
  INV_X1    g147(.A(KEYINPUT34), .ZN(new_n349));
  INV_X1    g148(.A(new_n340), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n349), .B1(new_n348), .B2(new_n350), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n352), .A2(new_n353), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n356), .A2(new_n346), .A3(new_n345), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n314), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT0), .ZN(new_n361));
  XNOR2_X1  g160(.A(G57gat), .B(G85gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  AND3_X1   g162(.A1(new_n326), .A2(new_n336), .A3(KEYINPUT76), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT76), .B1(new_n326), .B2(new_n336), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n286), .A2(KEYINPUT3), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n288), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n286), .A2(new_n337), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n286), .A2(KEYINPUT4), .A3(new_n337), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n376));
  OR3_X1    g175(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n337), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n326), .A2(new_n336), .A3(KEYINPUT76), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n286), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT78), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT78), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n380), .A2(new_n384), .A3(new_n286), .A4(new_n381), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n369), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n376), .B1(new_n386), .B2(new_n374), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT80), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT80), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n389), .B(new_n376), .C1(new_n386), .C2(new_n374), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n368), .A2(new_n374), .ZN(new_n392));
  INV_X1    g191(.A(new_n369), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT4), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT77), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n372), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n371), .A2(KEYINPUT77), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n392), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n378), .B1(new_n391), .B2(new_n399), .ZN(new_n400));
  AOI211_X1 g199(.A(KEYINPUT81), .B(new_n398), .C1(new_n388), .C2(new_n390), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n363), .B(new_n377), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n384), .B1(new_n366), .B2(new_n286), .ZN(new_n405));
  INV_X1    g204(.A(new_n385), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n393), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n375), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n389), .B1(new_n408), .B2(new_n376), .ZN(new_n409));
  INV_X1    g208(.A(new_n390), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n399), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT81), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n391), .A2(new_n378), .A3(new_n399), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n363), .B1(new_n414), .B2(new_n377), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n404), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n377), .B1(new_n400), .B2(new_n401), .ZN(new_n417));
  INV_X1    g216(.A(new_n363), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(KEYINPUT6), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n267), .B(new_n359), .C1(new_n416), .C2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT35), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n417), .A2(new_n418), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(new_n403), .A3(new_n402), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n419), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT35), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n267), .A4(new_n359), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  AOI211_X1 g228(.A(new_n266), .B(new_n358), .C1(new_n425), .C2(new_n419), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT86), .B1(new_n430), .B2(new_n427), .ZN(new_n431));
  INV_X1    g230(.A(new_n314), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n373), .A2(new_n375), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT39), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n375), .B2(new_n407), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n418), .B1(new_n433), .B2(new_n434), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n438), .B(KEYINPUT40), .Z(new_n439));
  NOR2_X1   g238(.A1(new_n267), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n432), .B1(new_n440), .B2(new_n424), .ZN(new_n441));
  INV_X1    g240(.A(new_n209), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n261), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT37), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n249), .A2(new_n243), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(new_n209), .ZN(new_n446));
  AOI211_X1 g245(.A(KEYINPUT38), .B(new_n263), .C1(new_n443), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n262), .A2(new_n444), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n447), .A2(new_n448), .B1(new_n262), .B2(new_n263), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n425), .A2(new_n419), .A3(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n450), .A2(KEYINPUT85), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT85), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n425), .A2(new_n452), .A3(new_n419), .A4(new_n449), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n448), .A2(new_n255), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n262), .A2(new_n444), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT38), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n441), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n314), .B1(new_n426), .B2(new_n267), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n355), .A2(new_n357), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT70), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n461), .A2(KEYINPUT70), .A3(KEYINPUT36), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n429), .A2(new_n431), .B1(new_n458), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT88), .B(G1gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT89), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT16), .ZN(new_n471));
  XNOR2_X1  g270(.A(G15gat), .B(G22gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n470), .B1(new_n469), .B2(KEYINPUT16), .ZN(new_n474));
  OAI22_X1  g273(.A1(new_n473), .A2(new_n474), .B1(G1gat), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT90), .B1(new_n472), .B2(G1gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(G8gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n475), .B(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n478), .B(KEYINPUT91), .Z(new_n479));
  XNOR2_X1  g278(.A(G43gat), .B(G50gat), .ZN(new_n480));
  OR3_X1    g279(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n481), .A2(new_n482), .B1(G29gat), .B2(G36gat), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n480), .B1(new_n483), .B2(KEYINPUT15), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(KEYINPUT15), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n484), .B(new_n485), .Z(new_n486));
  INV_X1    g285(.A(KEYINPUT17), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n479), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n478), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n489), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G229gat), .A2(G233gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT18), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n491), .A2(KEYINPUT18), .A3(new_n492), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n478), .B(new_n486), .Z(new_n497));
  XOR2_X1   g296(.A(new_n492), .B(KEYINPUT13), .Z(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G113gat), .B(G141gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(G169gat), .B(G197gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XOR2_X1   g302(.A(KEYINPUT87), .B(KEYINPUT11), .Z(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n505), .B(KEYINPUT12), .Z(new_n506));
  NAND2_X1  g305(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n506), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n495), .A2(new_n496), .A3(new_n499), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n468), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(G57gat), .A2(G64gat), .ZN(new_n513));
  AND2_X1   g312(.A1(G57gat), .A2(G64gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT9), .ZN(new_n515));
  NAND2_X1  g314(.A1(G71gat), .A2(G78gat), .ZN(new_n516));
  AOI211_X1 g315(.A(new_n513), .B(new_n514), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(G71gat), .A2(G78gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT92), .ZN(new_n519));
  INV_X1    g318(.A(new_n516), .ZN(new_n520));
  OR3_X1    g319(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OR3_X1    g320(.A1(new_n520), .A2(new_n518), .A3(KEYINPUT93), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT93), .B1(new_n520), .B2(new_n518), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n517), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT21), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G127gat), .B(G155gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n521), .A2(new_n524), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n490), .B1(KEYINPUT21), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n533), .B(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G183gat), .B(G211gat), .Z(new_n537));
  OR2_X1    g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G134gat), .B(G162gat), .Z(new_n541));
  AND2_X1   g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(KEYINPUT41), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n541), .B(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G85gat), .A2(G92gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  NAND2_X1  g345(.A1(G99gat), .A2(G106gat), .ZN(new_n547));
  INV_X1    g346(.A(G85gat), .ZN(new_n548));
  INV_X1    g347(.A(G92gat), .ZN(new_n549));
  AOI22_X1  g348(.A1(KEYINPUT8), .A2(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT94), .ZN(new_n551));
  XNOR2_X1  g350(.A(G99gat), .B(G106gat), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n546), .B(new_n550), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n551), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n553), .B(new_n554), .Z(new_n555));
  AOI22_X1  g354(.A1(new_n486), .A2(new_n555), .B1(KEYINPUT41), .B2(new_n542), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(new_n488), .B2(new_n555), .ZN(new_n557));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT95), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n544), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n560), .B2(new_n559), .ZN(new_n562));
  INV_X1    g361(.A(new_n559), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(KEYINPUT95), .A3(new_n544), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n540), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G230gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(new_n293), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n555), .A2(new_n534), .A3(KEYINPUT10), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT96), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n555), .B(new_n525), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT10), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n569), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n572), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n575), .B1(new_n576), .B2(new_n569), .ZN(new_n577));
  XNOR2_X1  g376(.A(G120gat), .B(G148gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT97), .ZN(new_n579));
  XOR2_X1   g378(.A(G176gat), .B(G204gat), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n577), .A2(new_n582), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n567), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n512), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n426), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n266), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT16), .B(G8gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n594), .B(KEYINPUT42), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(G8gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT98), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(G1325gat));
  AOI21_X1  g397(.A(G15gat), .B1(new_n588), .B2(new_n462), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n466), .A2(G15gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n600), .B(KEYINPUT99), .Z(new_n601));
  AOI21_X1  g400(.A(new_n599), .B1(new_n588), .B2(new_n601), .ZN(G1326gat));
  NOR2_X1   g401(.A1(new_n587), .A2(new_n314), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT43), .B(G22gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(G1327gat));
  NAND2_X1  g404(.A1(new_n458), .A2(new_n467), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n431), .A2(new_n423), .A3(new_n428), .ZN(new_n607));
  AOI211_X1 g406(.A(KEYINPUT44), .B(new_n566), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n607), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n565), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT101), .B1(new_n611), .B2(KEYINPUT44), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n566), .B1(new_n606), .B2(new_n607), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT44), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n609), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT102), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n540), .B(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n585), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n510), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n617), .A2(new_n618), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n614), .B1(new_n613), .B2(new_n615), .ZN(new_n625));
  OAI211_X1 g424(.A(KEYINPUT101), .B(KEYINPUT44), .C1(new_n468), .C2(new_n566), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n608), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(KEYINPUT102), .B1(new_n627), .B2(new_n622), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(G29gat), .B1(new_n629), .B2(new_n426), .ZN(new_n630));
  INV_X1    g429(.A(new_n540), .ZN(new_n631));
  AND4_X1   g430(.A1(new_n512), .A2(new_n631), .A3(new_n565), .A4(new_n621), .ZN(new_n632));
  INV_X1    g431(.A(G29gat), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n632), .A2(new_n633), .A3(new_n589), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT45), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n630), .A2(new_n635), .ZN(G1328gat));
  INV_X1    g435(.A(G36gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n632), .A2(new_n637), .A3(new_n266), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT103), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT46), .ZN(new_n640));
  OAI21_X1  g439(.A(G36gat), .B1(new_n629), .B2(new_n267), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(G1329gat));
  INV_X1    g441(.A(KEYINPUT47), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n624), .A2(new_n628), .A3(new_n466), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n645), .A3(G43gat), .ZN(new_n646));
  INV_X1    g445(.A(G43gat), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n632), .A2(new_n647), .A3(new_n462), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n645), .B1(new_n644), .B2(G43gat), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n643), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n617), .A2(new_n623), .ZN(new_n652));
  INV_X1    g451(.A(new_n466), .ZN(new_n653));
  OAI21_X1  g452(.A(G43gat), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n654), .A2(KEYINPUT47), .A3(new_n648), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n655), .ZN(G1330gat));
  OAI21_X1  g455(.A(KEYINPUT105), .B1(new_n652), .B2(new_n314), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n617), .A2(new_n658), .A3(new_n432), .A4(new_n623), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(G50gat), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n314), .A2(G50gat), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n632), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT48), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n660), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n661), .B1(new_n660), .B2(new_n665), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n624), .A2(new_n628), .A3(new_n432), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n663), .B1(new_n668), .B2(G50gat), .ZN(new_n669));
  OAI22_X1  g468(.A1(new_n666), .A2(new_n667), .B1(KEYINPUT48), .B2(new_n669), .ZN(G1331gat));
  NOR2_X1   g469(.A1(new_n567), .A2(new_n510), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n610), .A2(new_n585), .A3(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n672), .A2(KEYINPUT107), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(KEYINPUT107), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n589), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n266), .ZN(new_n679));
  NOR2_X1   g478(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n680));
  AND2_X1   g479(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n680), .B2(new_n679), .ZN(G1333gat));
  NAND3_X1  g482(.A1(new_n676), .A2(G71gat), .A3(new_n466), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n675), .A2(new_n461), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n684), .B1(G71gat), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g486(.A1(new_n676), .A2(new_n432), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g488(.A1(new_n540), .A2(new_n510), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n613), .B(new_n690), .C1(new_n691), .C2(KEYINPUT51), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n691), .A2(KEYINPUT51), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n694), .A2(new_n585), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(G85gat), .B1(new_n696), .B2(new_n589), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n690), .A2(new_n585), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n627), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n426), .A2(new_n548), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n697), .B1(new_n699), .B2(new_n700), .ZN(G1336gat));
  NAND3_X1  g500(.A1(new_n696), .A2(new_n549), .A3(new_n266), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n617), .A2(new_n585), .A3(new_n690), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n267), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n549), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT52), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n704), .A2(KEYINPUT109), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(KEYINPUT109), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n549), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT52), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n702), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n706), .B1(new_n709), .B2(new_n711), .ZN(G1337gat));
  AOI21_X1  g511(.A(G99gat), .B1(new_n696), .B2(new_n462), .ZN(new_n713));
  INV_X1    g512(.A(G99gat), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n703), .A2(new_n714), .A3(new_n653), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n713), .A2(new_n715), .ZN(G1338gat));
  INV_X1    g515(.A(G106gat), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n699), .B2(new_n432), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n314), .A2(G106gat), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n694), .A2(new_n585), .A3(new_n695), .A4(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT53), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT110), .B1(new_n699), .B2(new_n432), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n724));
  NOR4_X1   g523(.A1(new_n627), .A2(new_n724), .A3(new_n314), .A4(new_n698), .ZN(new_n725));
  OAI21_X1  g524(.A(G106gat), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n721), .A2(KEYINPUT53), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n727), .B1(new_n726), .B2(new_n728), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n722), .B1(new_n729), .B2(new_n730), .ZN(G1339gat));
  NOR2_X1   g530(.A1(new_n491), .A2(new_n492), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n497), .A2(new_n498), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n505), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n565), .A2(new_n509), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT54), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n575), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n571), .A2(new_n574), .A3(new_n569), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g539(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n741));
  AOI21_X1  g540(.A(new_n582), .B1(new_n575), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n736), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n740), .A2(KEYINPUT55), .A3(new_n742), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n584), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n743), .A2(new_n736), .A3(new_n744), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n746), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n735), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n565), .A2(new_n509), .A3(new_n734), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n746), .A2(new_n749), .A3(new_n750), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT114), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n510), .A2(new_n746), .A3(new_n749), .A4(new_n750), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n585), .A2(new_n509), .A3(new_n734), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n565), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n620), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n671), .A2(new_n621), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n426), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n267), .A3(new_n359), .ZN(new_n764));
  OAI21_X1  g563(.A(G113gat), .B1(new_n764), .B2(new_n511), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n510), .A2(new_n328), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT115), .Z(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n764), .B2(new_n767), .ZN(G1340gat));
  NOR2_X1   g567(.A1(new_n764), .A2(new_n621), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(new_n330), .ZN(G1341gat));
  OAI21_X1  g569(.A(G127gat), .B1(new_n764), .B2(new_n620), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n540), .A2(new_n319), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n764), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT116), .ZN(G1342gat));
  NOR2_X1   g573(.A1(new_n566), .A2(new_n266), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n358), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n763), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n777), .B(new_n778), .Z(G1343gat));
  NOR2_X1   g578(.A1(new_n466), .A2(new_n314), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n763), .A2(KEYINPUT117), .A3(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n785), .A2(new_n266), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n511), .A2(G141gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT58), .ZN(new_n789));
  INV_X1    g588(.A(new_n284), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n466), .A2(new_n426), .A3(new_n266), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n743), .A2(new_n744), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n749), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n759), .B1(new_n511), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n566), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(new_n756), .A3(new_n753), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n631), .ZN(new_n798));
  AOI211_X1 g597(.A(new_n792), .B(new_n314), .C1(new_n798), .C2(new_n762), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n314), .B1(new_n761), .B2(new_n762), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(KEYINPUT57), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n791), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n790), .B1(new_n802), .B2(new_n511), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n789), .A3(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n763), .A2(new_n267), .A3(new_n780), .A4(new_n787), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n806), .B2(new_n789), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n804), .B(KEYINPUT118), .C1(new_n789), .C2(new_n806), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(G1344gat));
  NAND3_X1  g610(.A1(new_n786), .A2(new_n282), .A3(new_n585), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n762), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n671), .A2(KEYINPUT120), .A3(new_n621), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n796), .B1(new_n755), .B2(new_n754), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n815), .A2(new_n816), .B1(new_n817), .B2(new_n631), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n792), .B1(new_n818), .B2(new_n314), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n800), .A2(new_n820), .A3(KEYINPUT57), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n800), .B2(KEYINPUT57), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n585), .A3(new_n791), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n813), .B1(new_n824), .B2(G148gat), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n802), .A2(new_n621), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(KEYINPUT59), .A3(new_n282), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n812), .B1(new_n825), .B2(new_n827), .ZN(G1345gat));
  NAND3_X1  g627(.A1(new_n786), .A2(new_n271), .A3(new_n540), .ZN(new_n829));
  OAI21_X1  g628(.A(G155gat), .B1(new_n802), .B2(new_n620), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(G1346gat));
  OAI21_X1  g630(.A(KEYINPUT121), .B1(new_n802), .B2(new_n566), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(G162gat), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n802), .A2(KEYINPUT121), .A3(new_n566), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n775), .A2(new_n272), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n833), .A2(new_n834), .B1(new_n785), .B2(new_n835), .ZN(G1347gat));
  AOI211_X1 g635(.A(new_n589), .B(new_n267), .C1(new_n761), .C2(new_n762), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n359), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n510), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G169gat), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT122), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(G169gat), .B2(new_n840), .ZN(G1348gat));
  NAND2_X1  g642(.A1(new_n839), .A2(new_n585), .ZN(new_n844));
  INV_X1    g643(.A(G176gat), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n844), .A2(KEYINPUT123), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT123), .B1(new_n844), .B2(new_n845), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n844), .A2(new_n845), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(G1349gat));
  OAI21_X1  g648(.A(G183gat), .B1(new_n838), .B2(new_n620), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n540), .A2(new_n228), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n850), .B1(new_n838), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g651(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n852), .B(new_n853), .ZN(G1350gat));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n565), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(G190gat), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT125), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(G190gat), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT126), .B1(new_n858), .B2(KEYINPUT61), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(KEYINPUT61), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n858), .A2(KEYINPUT126), .A3(KEYINPUT61), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n857), .B1(new_n861), .B2(new_n862), .ZN(G1351gat));
  AND2_X1   g662(.A1(new_n837), .A2(new_n780), .ZN(new_n864));
  AOI21_X1  g663(.A(G197gat), .B1(new_n864), .B2(new_n510), .ZN(new_n865));
  INV_X1    g664(.A(new_n823), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n589), .A2(new_n267), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n653), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n510), .A2(G197gat), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n865), .B1(new_n869), .B2(new_n870), .ZN(G1352gat));
  INV_X1    g670(.A(G204gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n864), .A2(new_n872), .A3(new_n585), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT62), .Z(new_n874));
  NOR3_X1   g673(.A1(new_n866), .A2(new_n621), .A3(new_n868), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(new_n872), .ZN(G1353gat));
  NAND3_X1  g675(.A1(new_n864), .A2(new_n204), .A3(new_n540), .ZN(new_n877));
  INV_X1    g676(.A(new_n868), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n823), .A2(new_n540), .A3(new_n878), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n879), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT63), .B1(new_n879), .B2(G211gat), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT127), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT127), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n884), .B(new_n877), .C1(new_n880), .C2(new_n881), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(G1354gat));
  NAND3_X1  g685(.A1(new_n864), .A2(new_n205), .A3(new_n565), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n866), .A2(new_n566), .A3(new_n868), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(new_n205), .ZN(G1355gat));
endmodule


