

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U322 ( .A(KEYINPUT47), .B(KEYINPUT119), .ZN(n384) );
  XNOR2_X1 U323 ( .A(n460), .B(n459), .ZN(n568) );
  XNOR2_X1 U324 ( .A(n385), .B(n384), .ZN(n392) );
  XNOR2_X1 U325 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U326 ( .A(n493), .B(n492), .ZN(n502) );
  XOR2_X1 U327 ( .A(KEYINPUT79), .B(KEYINPUT20), .Z(n290) );
  XNOR2_X1 U328 ( .A(n441), .B(n440), .ZN(n442) );
  NOR2_X1 U329 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U330 ( .A(n458), .B(KEYINPUT95), .ZN(n459) );
  XNOR2_X1 U331 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U332 ( .A(n446), .B(n290), .ZN(n447) );
  XNOR2_X1 U333 ( .A(n340), .B(n339), .ZN(n386) );
  XNOR2_X1 U334 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U335 ( .A(n394), .B(n393), .ZN(n547) );
  INV_X1 U336 ( .A(KEYINPUT108), .ZN(n496) );
  XNOR2_X1 U337 ( .A(n452), .B(G190GAT), .ZN(n453) );
  XNOR2_X1 U338 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U339 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(G169GAT), .B(G8GAT), .Z(n356) );
  XOR2_X1 U341 ( .A(KEYINPUT94), .B(KEYINPUT92), .Z(n292) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(KEYINPUT93), .ZN(n291) );
  XNOR2_X1 U343 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U344 ( .A(n356), .B(n293), .Z(n295) );
  NAND2_X1 U345 ( .A1(G226GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n300) );
  INV_X1 U347 ( .A(G204GAT), .ZN(n299) );
  XOR2_X1 U348 ( .A(G92GAT), .B(G64GAT), .Z(n297) );
  XNOR2_X1 U349 ( .A(G176GAT), .B(KEYINPUT73), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n334) );
  XOR2_X1 U352 ( .A(n300), .B(n334), .Z(n310) );
  XOR2_X1 U353 ( .A(G183GAT), .B(KEYINPUT17), .Z(n302) );
  XNOR2_X1 U354 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U356 ( .A(n303), .B(KEYINPUT18), .Z(n305) );
  XNOR2_X1 U357 ( .A(KEYINPUT81), .B(G190GAT), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n450) );
  XOR2_X1 U359 ( .A(KEYINPUT21), .B(G218GAT), .Z(n307) );
  XNOR2_X1 U360 ( .A(KEYINPUT84), .B(G211GAT), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U362 ( .A(G197GAT), .B(n308), .Z(n429) );
  XNOR2_X1 U363 ( .A(n450), .B(n429), .ZN(n309) );
  XNOR2_X1 U364 ( .A(n310), .B(n309), .ZN(n519) );
  INV_X1 U365 ( .A(KEYINPUT48), .ZN(n394) );
  XNOR2_X1 U366 ( .A(G183GAT), .B(G127GAT), .ZN(n312) );
  XNOR2_X1 U367 ( .A(G15GAT), .B(G22GAT), .ZN(n355) );
  INV_X1 U368 ( .A(n355), .ZN(n311) );
  XOR2_X1 U369 ( .A(n312), .B(n311), .Z(n325) );
  XOR2_X1 U370 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n314) );
  NAND2_X1 U371 ( .A1(G231GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U373 ( .A(KEYINPUT13), .B(G71GAT), .Z(n327) );
  XOR2_X1 U374 ( .A(n315), .B(n327), .Z(n323) );
  XOR2_X1 U375 ( .A(G57GAT), .B(G78GAT), .Z(n317) );
  XNOR2_X1 U376 ( .A(G155GAT), .B(G211GAT), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U378 ( .A(KEYINPUT12), .B(G64GAT), .Z(n319) );
  XNOR2_X1 U379 ( .A(G8GAT), .B(G1GAT), .ZN(n318) );
  XNOR2_X1 U380 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U381 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U383 ( .A(n325), .B(n324), .Z(n537) );
  INV_X1 U384 ( .A(n537), .ZN(n579) );
  XOR2_X1 U385 ( .A(KEYINPUT117), .B(KEYINPUT46), .Z(n326) );
  XNOR2_X1 U386 ( .A(KEYINPUT116), .B(n326), .ZN(n361) );
  XOR2_X1 U387 ( .A(G99GAT), .B(G85GAT), .Z(n364) );
  XOR2_X1 U388 ( .A(n327), .B(n364), .Z(n329) );
  XOR2_X1 U389 ( .A(G106GAT), .B(G78GAT), .Z(n422) );
  XOR2_X1 U390 ( .A(G120GAT), .B(G57GAT), .Z(n409) );
  XNOR2_X1 U391 ( .A(n422), .B(n409), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U393 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n331) );
  NAND2_X1 U394 ( .A1(G230GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U395 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U396 ( .A(n333), .B(n332), .Z(n340) );
  XNOR2_X1 U397 ( .A(n334), .B(KEYINPUT32), .ZN(n338) );
  XOR2_X1 U398 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n336) );
  XNOR2_X1 U399 ( .A(G148GAT), .B(KEYINPUT74), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n337) );
  INV_X1 U401 ( .A(KEYINPUT64), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n386), .B(n341), .ZN(n342) );
  XOR2_X1 U403 ( .A(n342), .B(KEYINPUT41), .Z(n533) );
  INV_X1 U404 ( .A(n533), .ZN(n560) );
  XNOR2_X1 U405 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n343) );
  XNOR2_X1 U406 ( .A(n343), .B(G36GAT), .ZN(n344) );
  XOR2_X1 U407 ( .A(n344), .B(KEYINPUT68), .Z(n346) );
  XNOR2_X1 U408 ( .A(G50GAT), .B(KEYINPUT8), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n346), .B(n345), .ZN(n376) );
  XOR2_X1 U410 ( .A(G1GAT), .B(G141GAT), .Z(n348) );
  XNOR2_X1 U411 ( .A(G29GAT), .B(G113GAT), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n410) );
  XOR2_X1 U413 ( .A(n410), .B(KEYINPUT29), .Z(n350) );
  NAND2_X1 U414 ( .A1(G229GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U416 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n352) );
  XNOR2_X1 U417 ( .A(G197GAT), .B(KEYINPUT67), .ZN(n351) );
  XNOR2_X1 U418 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U419 ( .A(n354), .B(n353), .Z(n358) );
  XOR2_X1 U420 ( .A(n356), .B(n355), .Z(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n376), .B(n359), .ZN(n571) );
  NAND2_X1 U423 ( .A1(n560), .A2(n571), .ZN(n360) );
  XOR2_X1 U424 ( .A(n361), .B(n360), .Z(n362) );
  NOR2_X1 U425 ( .A1(n579), .A2(n362), .ZN(n363) );
  XNOR2_X1 U426 ( .A(KEYINPUT118), .B(n363), .ZN(n383) );
  XOR2_X1 U427 ( .A(KEYINPUT65), .B(n364), .Z(n366) );
  XNOR2_X1 U428 ( .A(G218GAT), .B(KEYINPUT75), .ZN(n365) );
  XNOR2_X1 U429 ( .A(n366), .B(n365), .ZN(n380) );
  XOR2_X1 U430 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n368) );
  XNOR2_X1 U431 ( .A(G106GAT), .B(G92GAT), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U433 ( .A(KEYINPUT66), .B(G162GAT), .Z(n370) );
  XNOR2_X1 U434 ( .A(G190GAT), .B(G134GAT), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U436 ( .A(n372), .B(n371), .Z(n378) );
  XOR2_X1 U437 ( .A(KEYINPUT77), .B(KEYINPUT9), .Z(n374) );
  XNOR2_X1 U438 ( .A(G29GAT), .B(KEYINPUT76), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U440 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U442 ( .A(n380), .B(n379), .Z(n382) );
  NAND2_X1 U443 ( .A1(G232GAT), .A2(G233GAT), .ZN(n381) );
  XOR2_X1 U444 ( .A(n382), .B(n381), .Z(n555) );
  INV_X1 U445 ( .A(n555), .ZN(n541) );
  NAND2_X1 U446 ( .A1(n383), .A2(n541), .ZN(n385) );
  XOR2_X1 U447 ( .A(n555), .B(KEYINPUT106), .Z(n387) );
  XNOR2_X1 U448 ( .A(n387), .B(KEYINPUT36), .ZN(n583) );
  NOR2_X1 U449 ( .A1(n583), .A2(n537), .ZN(n388) );
  XOR2_X1 U450 ( .A(KEYINPUT45), .B(n388), .Z(n389) );
  NOR2_X1 U451 ( .A1(n386), .A2(n389), .ZN(n390) );
  XOR2_X1 U452 ( .A(KEYINPUT70), .B(n571), .Z(n557) );
  NAND2_X1 U453 ( .A1(n390), .A2(n557), .ZN(n391) );
  NAND2_X1 U454 ( .A1(n392), .A2(n391), .ZN(n393) );
  NOR2_X1 U455 ( .A1(n519), .A2(n547), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n395), .B(KEYINPUT54), .ZN(n567) );
  XOR2_X1 U457 ( .A(KEYINPUT2), .B(G162GAT), .Z(n397) );
  XNOR2_X1 U458 ( .A(G155GAT), .B(G148GAT), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U460 ( .A(KEYINPUT3), .B(n398), .ZN(n430) );
  INV_X1 U461 ( .A(n430), .ZN(n418) );
  XOR2_X1 U462 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n400) );
  XNOR2_X1 U463 ( .A(KEYINPUT89), .B(KEYINPUT85), .ZN(n399) );
  XNOR2_X1 U464 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U465 ( .A(KEYINPUT1), .B(KEYINPUT86), .Z(n402) );
  XNOR2_X1 U466 ( .A(KEYINPUT6), .B(KEYINPUT4), .ZN(n401) );
  XNOR2_X1 U467 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U468 ( .A(n404), .B(n403), .Z(n416) );
  XOR2_X1 U469 ( .A(G127GAT), .B(KEYINPUT0), .Z(n406) );
  XNOR2_X1 U470 ( .A(G134GAT), .B(KEYINPUT78), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n406), .B(n405), .ZN(n446) );
  XOR2_X1 U472 ( .A(n446), .B(KEYINPUT5), .Z(n408) );
  NAND2_X1 U473 ( .A1(G225GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U474 ( .A(n408), .B(n407), .ZN(n414) );
  XOR2_X1 U475 ( .A(n409), .B(KEYINPUT90), .Z(n412) );
  XNOR2_X1 U476 ( .A(n410), .B(G85GAT), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U480 ( .A(n418), .B(n417), .Z(n466) );
  XOR2_X1 U481 ( .A(KEYINPUT91), .B(n466), .Z(n545) );
  XOR2_X1 U482 ( .A(G204GAT), .B(KEYINPUT75), .Z(n420) );
  XNOR2_X1 U483 ( .A(G50GAT), .B(G141GAT), .ZN(n419) );
  XNOR2_X1 U484 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U485 ( .A(n422), .B(n421), .Z(n424) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U488 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n426) );
  XNOR2_X1 U489 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n425) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U491 ( .A(n428), .B(n427), .Z(n432) );
  XOR2_X1 U492 ( .A(n430), .B(n429), .Z(n431) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n468) );
  NOR2_X1 U494 ( .A1(n545), .A2(n468), .ZN(n433) );
  AND2_X1 U495 ( .A1(n567), .A2(n433), .ZN(n435) );
  XNOR2_X1 U496 ( .A(KEYINPUT124), .B(KEYINPUT55), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n435), .B(n434), .ZN(n451) );
  XOR2_X1 U498 ( .A(G71GAT), .B(G120GAT), .Z(n437) );
  XNOR2_X1 U499 ( .A(G169GAT), .B(G113GAT), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n445) );
  XOR2_X1 U501 ( .A(G176GAT), .B(KEYINPUT80), .Z(n439) );
  XNOR2_X1 U502 ( .A(G15GAT), .B(KEYINPUT83), .ZN(n438) );
  XNOR2_X1 U503 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U504 ( .A(G43GAT), .B(G99GAT), .Z(n441) );
  NAND2_X1 U505 ( .A1(G227GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n457) );
  NOR2_X2 U508 ( .A1(n451), .A2(n457), .ZN(n564) );
  NAND2_X1 U509 ( .A1(n564), .A2(n555), .ZN(n454) );
  XOR2_X1 U510 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n452) );
  NOR2_X1 U511 ( .A1(n557), .A2(n386), .ZN(n491) );
  NOR2_X1 U512 ( .A1(n519), .A2(n457), .ZN(n455) );
  NOR2_X1 U513 ( .A1(n468), .A2(n455), .ZN(n456) );
  XOR2_X1 U514 ( .A(KEYINPUT25), .B(n456), .Z(n463) );
  XOR2_X1 U515 ( .A(n519), .B(KEYINPUT27), .Z(n469) );
  INV_X1 U516 ( .A(n469), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n468), .A2(n457), .ZN(n460) );
  XOR2_X1 U518 ( .A(KEYINPUT96), .B(KEYINPUT26), .Z(n458) );
  NOR2_X1 U519 ( .A1(n461), .A2(n568), .ZN(n544) );
  XOR2_X1 U520 ( .A(n544), .B(KEYINPUT97), .Z(n462) );
  NOR2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT98), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n467), .B(KEYINPUT99), .ZN(n472) );
  INV_X1 U524 ( .A(n545), .ZN(n566) );
  XOR2_X1 U525 ( .A(n468), .B(KEYINPUT28), .Z(n525) );
  NAND2_X1 U526 ( .A1(n469), .A2(n525), .ZN(n470) );
  NOR2_X1 U527 ( .A1(n566), .A2(n470), .ZN(n529) );
  NAND2_X1 U528 ( .A1(n529), .A2(n457), .ZN(n471) );
  NAND2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n488) );
  NAND2_X1 U530 ( .A1(n541), .A2(n579), .ZN(n473) );
  XOR2_X1 U531 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  AND2_X1 U532 ( .A1(n488), .A2(n474), .ZN(n506) );
  NAND2_X1 U533 ( .A1(n491), .A2(n506), .ZN(n475) );
  XNOR2_X1 U534 ( .A(KEYINPUT100), .B(n475), .ZN(n486) );
  NOR2_X1 U535 ( .A1(n486), .A2(n566), .ZN(n480) );
  XOR2_X1 U536 ( .A(KEYINPUT34), .B(KEYINPUT103), .Z(n477) );
  XNOR2_X1 U537 ( .A(G1GAT), .B(KEYINPUT102), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U539 ( .A(KEYINPUT101), .B(n478), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(G1324GAT) );
  NOR2_X1 U541 ( .A1(n519), .A2(n486), .ZN(n481) );
  XOR2_X1 U542 ( .A(G8GAT), .B(n481), .Z(G1325GAT) );
  NOR2_X1 U543 ( .A1(n457), .A2(n486), .ZN(n485) );
  XOR2_X1 U544 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n483) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT105), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n525), .A2(n486), .ZN(n487) );
  XOR2_X1 U549 ( .A(G22GAT), .B(n487), .Z(G1327GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT38), .B(KEYINPUT107), .Z(n493) );
  NOR2_X1 U551 ( .A1(n579), .A2(n583), .ZN(n489) );
  NAND2_X1 U552 ( .A1(n489), .A2(n488), .ZN(n490) );
  XNOR2_X1 U553 ( .A(KEYINPUT37), .B(n490), .ZN(n517) );
  NAND2_X1 U554 ( .A1(n491), .A2(n517), .ZN(n492) );
  NOR2_X1 U555 ( .A1(n502), .A2(n566), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U558 ( .A1(n519), .A2(n502), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(n498), .ZN(G1329GAT) );
  NOR2_X1 U560 ( .A1(n502), .A2(n457), .ZN(n500) );
  XNOR2_X1 U561 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NOR2_X1 U564 ( .A1(n525), .A2(n502), .ZN(n503) );
  XOR2_X1 U565 ( .A(KEYINPUT110), .B(n503), .Z(n504) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n504), .ZN(G1331GAT) );
  NOR2_X1 U567 ( .A1(n533), .A2(n571), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n505), .B(KEYINPUT112), .ZN(n516) );
  NAND2_X1 U569 ( .A1(n516), .A2(n506), .ZN(n507) );
  XOR2_X1 U570 ( .A(KEYINPUT113), .B(n507), .Z(n513) );
  NOR2_X1 U571 ( .A1(n566), .A2(n513), .ZN(n509) );
  XNOR2_X1 U572 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n519), .A2(n513), .ZN(n511) );
  XOR2_X1 U576 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U577 ( .A1(n457), .A2(n513), .ZN(n512) );
  XOR2_X1 U578 ( .A(G71GAT), .B(n512), .Z(G1334GAT) );
  NOR2_X1 U579 ( .A1(n525), .A2(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  NAND2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n524) );
  NOR2_X1 U583 ( .A1(n566), .A2(n524), .ZN(n518) );
  XOR2_X1 U584 ( .A(G85GAT), .B(n518), .Z(G1336GAT) );
  NOR2_X1 U585 ( .A1(n519), .A2(n524), .ZN(n520) );
  XOR2_X1 U586 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  NOR2_X1 U587 ( .A1(n457), .A2(n524), .ZN(n521) );
  XOR2_X1 U588 ( .A(G99GAT), .B(n521), .Z(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT114), .Z(n523) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(KEYINPUT115), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(n527) );
  NOR2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U593 ( .A(n527), .B(n526), .Z(G1339GAT) );
  NOR2_X1 U594 ( .A1(n457), .A2(n547), .ZN(n528) );
  NAND2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(KEYINPUT120), .B(n530), .ZN(n540) );
  NOR2_X1 U597 ( .A1(n540), .A2(n557), .ZN(n532) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(KEYINPUT121), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(G1340GAT) );
  NOR2_X1 U600 ( .A1(n540), .A2(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(KEYINPUT122), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(n536), .ZN(G1341GAT) );
  NOR2_X1 U604 ( .A1(n540), .A2(n537), .ZN(n538) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(n538), .Z(n539) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n543) );
  NOR2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n571), .A2(n554), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n548), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  NAND2_X1 U615 ( .A1(n554), .A2(n560), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n552) );
  XOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT123), .Z(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n554), .A2(n579), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 U623 ( .A(n557), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n564), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n564), .A2(n560), .ZN(n562) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G176GAT), .ZN(G1349GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n579), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n574) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n569) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  INV_X1 U635 ( .A(n570), .ZN(n582) );
  INV_X1 U636 ( .A(n582), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n572), .A2(n386), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  XOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT127), .Z(n581) );
  NAND2_X1 U645 ( .A1(n572), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

