//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G134), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT11), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(KEYINPUT11), .A3(G134), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G137), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(new_n196), .A3(new_n197), .A4(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n196), .B1(G134), .B2(G137), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n190), .A2(new_n192), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G137), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n200), .A2(KEYINPUT67), .A3(new_n203), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n208), .B(G146), .C1(new_n209), .C2(KEYINPUT1), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n211), .A3(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n211), .A2(G143), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n208), .A2(G146), .ZN(new_n220));
  AND4_X1   g034(.A1(new_n215), .A2(new_n217), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n214), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n206), .A2(new_n207), .A3(new_n222), .ZN(new_n223));
  OR2_X1    g037(.A1(KEYINPUT2), .A2(G113), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT2), .A2(G113), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  INV_X1    g041(.A(G119), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(G116), .A2(G119), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n230), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(new_n224), .A3(new_n225), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n219), .A2(new_n220), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT0), .A2(G128), .ZN(new_n237));
  NAND2_X1  g051(.A1(KEYINPUT0), .A2(G128), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n236), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n216), .A2(new_n238), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n200), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n197), .A2(new_n199), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n196), .B1(new_n245), .B2(new_n195), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n242), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n223), .A2(new_n235), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT28), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n222), .A2(new_n200), .A3(new_n203), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n247), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n234), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT28), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n250), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G237), .ZN(new_n257));
  INV_X1    g071(.A(G953), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(G210), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT27), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT26), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT27), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n259), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT26), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n261), .A2(new_n265), .A3(G101), .ZN(new_n266));
  AOI21_X1  g080(.A(G101), .B1(new_n261), .B2(new_n265), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n256), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n248), .A2(KEYINPUT69), .A3(new_n268), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT69), .B1(new_n248), .B2(new_n268), .ZN(new_n273));
  OR2_X1    g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT31), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT65), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n216), .A2(new_n215), .A3(new_n217), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n213), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(new_n204), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n282));
  OAI21_X1  g096(.A(G131), .B1(new_n282), .B2(new_n244), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n283), .A2(new_n200), .B1(new_n240), .B2(new_n241), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n276), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT66), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n223), .A2(KEYINPUT30), .A3(new_n247), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT66), .B(new_n276), .C1(new_n281), .C2(new_n284), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n287), .A2(new_n234), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n290), .A2(KEYINPUT68), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(KEYINPUT68), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n274), .B(new_n275), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT71), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n272), .A2(new_n273), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT66), .B1(new_n252), .B2(new_n276), .ZN(new_n296));
  AOI211_X1 g110(.A(new_n286), .B(KEYINPUT30), .C1(new_n251), .C2(new_n247), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT68), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n298), .A2(new_n299), .A3(new_n234), .A4(new_n288), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n290), .A2(KEYINPUT68), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n295), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(new_n275), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n271), .B1(new_n294), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n302), .B2(new_n275), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n274), .B1(new_n291), .B2(new_n292), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n188), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n300), .A2(new_n301), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n248), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n269), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n256), .A2(new_n269), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n223), .A2(new_n247), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n234), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n250), .A2(new_n255), .A3(new_n319), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n320), .A2(new_n315), .A3(new_n269), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(G902), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n311), .A2(KEYINPUT32), .B1(new_n323), .B2(G472), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n294), .A2(new_n304), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n310), .A2(new_n325), .A3(new_n270), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n187), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT32), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G478), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n331), .A2(KEYINPUT15), .ZN(new_n332));
  INV_X1    g146(.A(G107), .ZN(new_n333));
  XNOR2_X1  g147(.A(G116), .B(G122), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT92), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n334), .A2(KEYINPUT92), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n333), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n337), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n335), .A3(G107), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n208), .A2(G128), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n209), .A2(G143), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT95), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT95), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n190), .A3(new_n192), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n343), .A2(KEYINPUT13), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n342), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT93), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n209), .A2(G143), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n352), .B1(new_n353), .B2(KEYINPUT13), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n189), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT94), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n350), .A2(new_n352), .A3(new_n342), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n356), .B1(new_n355), .B2(new_n357), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n341), .B(new_n349), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n345), .A2(new_n202), .A3(new_n347), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n349), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n227), .A2(KEYINPUT14), .A3(G122), .ZN(new_n363));
  XOR2_X1   g177(.A(G116), .B(G122), .Z(new_n364));
  OAI211_X1 g178(.A(G107), .B(new_n363), .C1(new_n364), .C2(KEYINPUT14), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n365), .A2(KEYINPUT96), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(KEYINPUT96), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n362), .A2(new_n338), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT9), .B(G234), .ZN(new_n370));
  INV_X1    g184(.A(G217), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n370), .A2(new_n371), .A3(G953), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n360), .A2(new_n368), .A3(new_n372), .ZN(new_n375));
  AOI21_X1  g189(.A(G902), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT97), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n332), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G902), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n360), .A2(new_n368), .A3(new_n372), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n372), .B1(new_n360), .B2(new_n368), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT97), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n374), .A2(new_n375), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n377), .A3(new_n379), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n378), .B1(new_n386), .B2(new_n332), .ZN(new_n387));
  INV_X1    g201(.A(G475), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n257), .A2(new_n258), .A3(G214), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n208), .ZN(new_n390));
  NOR2_X1   g204(.A1(G237), .A2(G953), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(G143), .A3(G214), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G131), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT17), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT91), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n196), .B1(new_n390), .B2(new_n392), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT91), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT17), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G125), .B(G140), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT16), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT16), .ZN(new_n403));
  INV_X1    g217(.A(G140), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(G125), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(G146), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(G146), .B1(new_n402), .B2(new_n405), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT90), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n408), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT90), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(new_n406), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n390), .A2(new_n196), .A3(new_n392), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n394), .A2(new_n395), .A3(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n400), .A2(new_n409), .A3(new_n412), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(KEYINPUT18), .A2(G131), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n393), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n390), .A2(KEYINPUT18), .A3(G131), .A4(new_n392), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n404), .A2(G125), .ZN(new_n420));
  INV_X1    g234(.A(G125), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G140), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G146), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n401), .A2(new_n211), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n426), .B1(new_n424), .B2(new_n425), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n419), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n415), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G104), .ZN(new_n431));
  XNOR2_X1  g245(.A(G113), .B(G122), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n432), .A2(new_n433), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n436), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(G104), .A3(new_n434), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n430), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(KEYINPUT89), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT89), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n437), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n415), .A2(new_n429), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n388), .B1(new_n446), .B2(new_n379), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n394), .A2(new_n413), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n401), .A2(KEYINPUT19), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n401), .A2(KEYINPUT19), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n211), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(new_n406), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n429), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n453), .A2(new_n454), .A3(new_n440), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n454), .B1(new_n453), .B2(new_n440), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n445), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(G475), .A2(G902), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT20), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n461), .A3(new_n458), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n447), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G952), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n464), .A2(KEYINPUT98), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(KEYINPUT98), .ZN(new_n466));
  AOI21_X1  g280(.A(G953), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(G234), .A2(G237), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n469), .B(KEYINPUT99), .Z(new_n470));
  AND3_X1   g284(.A1(new_n468), .A2(G902), .A3(G953), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(G898), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n387), .A2(new_n463), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G221), .B1(new_n370), .B2(G902), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n210), .A2(KEYINPUT79), .A3(new_n212), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT79), .B1(new_n210), .B2(new_n212), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n278), .A2(new_n279), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT78), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n484), .B1(new_n431), .B2(G107), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n431), .A2(G107), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n333), .A2(KEYINPUT78), .A3(G104), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G101), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT3), .B1(new_n431), .B2(G107), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT3), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n333), .A3(G104), .ZN(new_n492));
  INV_X1    g306(.A(G101), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n490), .A2(new_n492), .A3(new_n493), .A4(new_n486), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n483), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT10), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n490), .A2(new_n492), .A3(new_n486), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(G101), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n499), .A2(G101), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n242), .B(new_n501), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n283), .A2(new_n200), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT80), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT80), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n283), .A2(new_n507), .A3(new_n200), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n495), .A2(new_n222), .A3(KEYINPUT10), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n498), .A2(new_n504), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n489), .A2(new_n494), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n280), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n496), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT12), .B1(new_n514), .B2(new_n505), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT12), .ZN(new_n516));
  INV_X1    g330(.A(new_n505), .ZN(new_n517));
  AOI211_X1 g331(.A(new_n516), .B(new_n517), .C1(new_n496), .C2(new_n513), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n511), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n258), .A2(G227), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(G140), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT77), .B(G110), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n512), .B1(new_n482), .B2(new_n481), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n510), .B(new_n504), .C1(new_n524), .C2(KEYINPUT10), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n506), .A2(new_n508), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(new_n523), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n505), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n519), .A2(new_n523), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(G469), .B1(new_n530), .B2(G902), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n511), .A2(new_n529), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n523), .ZN(new_n533));
  INV_X1    g347(.A(new_n523), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n511), .B(new_n534), .C1(new_n515), .C2(new_n518), .ZN(new_n535));
  AOI21_X1  g349(.A(G902), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT81), .B(G469), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n478), .B1(new_n531), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT23), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n228), .B2(G128), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n541), .B(new_n542), .C1(G119), .C2(new_n209), .ZN(new_n543));
  XNOR2_X1  g357(.A(G119), .B(G128), .ZN(new_n544));
  XOR2_X1   g358(.A(KEYINPUT24), .B(G110), .Z(new_n545));
  AOI22_X1  g359(.A1(new_n543), .A2(G110), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n407), .B2(new_n408), .ZN(new_n547));
  NAND2_X1  g361(.A1(G221), .A2(G234), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT74), .B1(new_n548), .B2(G953), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT74), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n550), .A2(new_n258), .A3(G221), .A4(G234), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT22), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n552), .B1(new_n549), .B2(new_n551), .ZN(new_n555));
  OR3_X1    g369(.A1(new_n554), .A2(new_n193), .A3(new_n555), .ZN(new_n556));
  OAI22_X1  g370(.A1(new_n543), .A2(G110), .B1(new_n544), .B2(new_n545), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(new_n406), .A3(new_n425), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n193), .B1(new_n554), .B2(new_n555), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n547), .A2(new_n556), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT76), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n547), .A2(new_n558), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n556), .A2(new_n559), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT75), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(KEYINPUT75), .A3(new_n564), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G234), .ZN(new_n571));
  OAI21_X1  g385(.A(G217), .B1(new_n571), .B2(G902), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT72), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(G902), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n573), .B(KEYINPUT73), .Z(new_n578));
  NAND3_X1  g392(.A1(new_n562), .A2(new_n569), .A3(new_n379), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n578), .B1(new_n579), .B2(KEYINPUT25), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT25), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n562), .A2(new_n569), .A3(new_n581), .A4(new_n379), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n577), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n539), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT85), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT84), .ZN(new_n586));
  XNOR2_X1  g400(.A(G110), .B(G122), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n587), .B(KEYINPUT8), .Z(new_n588));
  INV_X1    g402(.A(KEYINPUT5), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n229), .B2(new_n230), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n228), .A3(G116), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G113), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n233), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n512), .A2(new_n593), .ZN(new_n594));
  OR2_X1    g408(.A1(new_n590), .A2(new_n592), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n595), .A2(new_n233), .A3(new_n494), .A4(new_n489), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n588), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT83), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n242), .A2(G125), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n280), .B2(G125), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT82), .B(G224), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n258), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n604), .A2(KEYINPUT7), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n600), .B(new_n603), .C1(G125), .C2(new_n280), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n601), .A2(new_n606), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n586), .B1(new_n599), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n597), .B(KEYINPUT83), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n612), .A2(KEYINPUT84), .A3(new_n609), .A4(new_n608), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n234), .B(new_n501), .C1(new_n502), .C2(new_n503), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n596), .A3(new_n587), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n611), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(G210), .B1(G237), .B2(G902), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n614), .A2(new_n596), .ZN(new_n618));
  INV_X1    g432(.A(new_n587), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(KEYINPUT6), .A3(new_n615), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n605), .A2(new_n607), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT6), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n618), .A2(new_n623), .A3(new_n619), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n625), .A2(new_n379), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n616), .A2(new_n617), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n617), .B1(new_n616), .B2(new_n626), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(G214), .B1(G237), .B2(G902), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n585), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g447(.A(KEYINPUT85), .B(new_n631), .C1(new_n628), .C2(new_n629), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n476), .B(new_n584), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n330), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G101), .ZN(G3));
  NAND2_X1  g451(.A1(new_n326), .A2(new_n379), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n311), .B1(new_n638), .B2(G472), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n584), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n641), .B(KEYINPUT100), .Z(new_n642));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n384), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n374), .A2(KEYINPUT33), .A3(new_n375), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n331), .A2(G902), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n382), .A2(new_n331), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n463), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT102), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n616), .A2(new_n626), .ZN(new_n652));
  INV_X1    g466(.A(new_n617), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n655), .A3(new_n627), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n616), .A2(KEYINPUT101), .A3(new_n617), .A4(new_n626), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n657), .A2(new_n631), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n474), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n651), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n642), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT34), .B(G104), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT103), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n663), .B(new_n665), .ZN(G6));
  AND3_X1   g480(.A1(new_n457), .A2(new_n461), .A3(new_n458), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n461), .B1(new_n457), .B2(new_n458), .ZN(new_n668));
  AOI21_X1  g482(.A(G902), .B1(new_n441), .B2(new_n445), .ZN(new_n669));
  OAI22_X1  g483(.A1(new_n667), .A2(new_n668), .B1(new_n388), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n387), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n642), .A2(new_n660), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT35), .B(G107), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  OR2_X1    g488(.A1(new_n564), .A2(KEYINPUT36), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n563), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n576), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n580), .B2(new_n582), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n539), .A2(new_n679), .ZN(new_n680));
  AOI211_X1 g494(.A(new_n476), .B(new_n680), .C1(new_n633), .C2(new_n634), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n639), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT37), .B(G110), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G12));
  INV_X1    g498(.A(G900), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n471), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n470), .A2(new_n686), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n387), .A2(new_n670), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n689), .A2(new_n659), .A3(new_n680), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n293), .A2(KEYINPUT71), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n303), .B1(new_n302), .B2(new_n275), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n270), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n307), .A2(new_n309), .ZN(new_n694));
  OAI211_X1 g508(.A(KEYINPUT32), .B(new_n187), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n323), .A2(G472), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n311), .A2(KEYINPUT32), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n690), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G128), .ZN(G30));
  AOI21_X1  g514(.A(new_n268), .B1(new_n319), .B2(new_n248), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n379), .B1(new_n302), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(G472), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n329), .A2(new_n695), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n630), .B(KEYINPUT38), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n387), .A2(new_n463), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n631), .A3(new_n678), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT104), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n704), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n687), .B(KEYINPUT39), .Z(new_n714));
  NAND2_X1  g528(.A1(new_n539), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT106), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT40), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n712), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT107), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n208), .ZN(G45));
  NOR3_X1   g534(.A1(new_n649), .A2(new_n463), .A3(new_n687), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n722), .A2(new_n659), .A3(new_n680), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n697), .B2(new_n698), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G146), .ZN(G48));
  INV_X1    g539(.A(G469), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n536), .A2(new_n726), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n727), .A2(new_n477), .A3(new_n538), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n583), .B(new_n728), .C1(new_n697), .C2(new_n698), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT108), .B1(new_n729), .B2(new_n661), .ZN(new_n730));
  INV_X1    g544(.A(new_n583), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n324), .B2(new_n329), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n662), .A4(new_n728), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(KEYINPUT41), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G113), .ZN(G15));
  NAND2_X1  g551(.A1(new_n660), .A2(new_n671), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n729), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n227), .ZN(G18));
  INV_X1    g554(.A(new_n728), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n659), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n476), .A2(new_n678), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n742), .B(new_n743), .C1(new_n697), .C2(new_n698), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G119), .ZN(G21));
  AOI22_X1  g559(.A1(new_n308), .A2(KEYINPUT31), .B1(new_n269), .B2(new_n320), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n325), .A2(new_n746), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n638), .A2(G472), .B1(new_n187), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n727), .A2(new_n477), .A3(new_n538), .A4(new_n475), .ZN(new_n749));
  NOR4_X1   g563(.A1(new_n659), .A2(new_n463), .A3(new_n387), .A4(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n583), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G122), .ZN(G24));
  NAND2_X1  g566(.A1(new_n638), .A2(G472), .ZN(new_n753));
  AND4_X1   g567(.A1(new_n656), .A2(new_n721), .A3(new_n658), .A4(new_n728), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n747), .A2(new_n187), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n753), .A2(new_n754), .A3(new_n679), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  INV_X1    g571(.A(KEYINPUT42), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n628), .A2(new_n629), .A3(new_n632), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n511), .A2(new_n529), .A3(new_n534), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n514), .A2(KEYINPUT12), .A3(new_n505), .ZN(new_n761));
  INV_X1    g575(.A(new_n513), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n505), .B1(new_n762), .B2(new_n524), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n516), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n527), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  OAI211_X1 g579(.A(G469), .B(new_n760), .C1(new_n765), .C2(new_n534), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT110), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n519), .A2(new_n523), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n769), .A3(G469), .A4(new_n760), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(G469), .A2(G902), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT109), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n536), .B2(new_n537), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n478), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n759), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n583), .B(new_n777), .C1(new_n697), .C2(new_n698), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n758), .B1(new_n778), .B2(new_n722), .ZN(new_n779));
  OR3_X1    g593(.A1(new_n311), .A2(KEYINPUT111), .A3(KEYINPUT32), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT111), .B1(new_n311), .B2(KEYINPUT32), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n324), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n776), .A2(new_n722), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n758), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(new_n785), .A3(new_n583), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n779), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G131), .ZN(G33));
  AOI211_X1 g602(.A(new_n731), .B(new_n776), .C1(new_n324), .C2(new_n329), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n688), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  NOR2_X1   g605(.A1(new_n649), .A2(new_n670), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(KEYINPUT43), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n793), .A2(KEYINPUT113), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(KEYINPUT43), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n795), .B1(new_n793), .B2(KEYINPUT113), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n797), .A2(new_n639), .A3(new_n678), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n798), .A2(KEYINPUT44), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(KEYINPUT44), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n768), .A2(new_n760), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n726), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n802), .B2(new_n801), .ZN(new_n804));
  INV_X1    g618(.A(new_n773), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n806), .A2(new_n807), .A3(KEYINPUT46), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n806), .B2(KEYINPUT46), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n806), .A2(KEYINPUT46), .B1(new_n536), .B2(new_n537), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n477), .A3(new_n714), .ZN(new_n812));
  INV_X1    g626(.A(new_n759), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n799), .A2(new_n800), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G137), .ZN(G39));
  NAND2_X1  g630(.A1(new_n811), .A2(new_n477), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT47), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n330), .A2(new_n583), .A3(new_n722), .A4(new_n813), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G140), .ZN(G42));
  NAND2_X1  g636(.A1(new_n748), .A2(new_n583), .ZN(new_n823));
  INV_X1    g637(.A(new_n470), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n794), .B2(new_n796), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n706), .A2(new_n631), .A3(new_n741), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n828), .B(KEYINPUT50), .Z(new_n829));
  AND2_X1   g643(.A1(new_n727), .A2(new_n538), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(new_n478), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n759), .B(new_n826), .C1(new_n819), .C2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n704), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n813), .A2(new_n741), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n583), .A2(new_n833), .A3(new_n824), .A4(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n649), .A2(new_n463), .ZN(new_n836));
  AOI21_X1  g650(.A(G902), .B1(new_n305), .B2(new_n310), .ZN(new_n837));
  INV_X1    g651(.A(G472), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n679), .B(new_n755), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n824), .B(new_n834), .C1(new_n794), .C2(new_n796), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n835), .A2(new_n836), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n829), .A2(new_n832), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n829), .A2(new_n832), .A3(KEYINPUT51), .A4(new_n843), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n835), .A2(new_n651), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n826), .A2(new_n742), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n467), .A3(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n782), .A2(new_n583), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n842), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n852), .A2(KEYINPUT48), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(KEYINPUT48), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n846), .A2(new_n847), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n856), .B(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n769), .B1(new_n530), .B2(G469), .ZN(new_n859));
  INV_X1    g673(.A(new_n770), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n774), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI211_X1 g675(.A(new_n687), .B(new_n677), .C1(new_n580), .C2(new_n582), .ZN(new_n862));
  AND4_X1   g676(.A1(KEYINPUT116), .A2(new_n861), .A3(new_n862), .A4(new_n477), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT116), .B1(new_n775), .B2(new_n862), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n656), .A2(new_n707), .A3(new_n658), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n703), .B1(new_n311), .B2(KEYINPUT32), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n328), .B(new_n188), .C1(new_n305), .C2(new_n310), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n865), .B(new_n866), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n724), .A3(KEYINPUT52), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n699), .A2(new_n871), .A3(new_n756), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n656), .A2(new_n658), .ZN(new_n873));
  INV_X1    g687(.A(new_n680), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n874), .A3(new_n688), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n324), .B2(new_n329), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n873), .A2(new_n721), .A3(new_n728), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n839), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT115), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n870), .B1(new_n872), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n866), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n881), .A2(new_n864), .A3(new_n863), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n882), .A2(new_n704), .B1(new_n330), .B2(new_n723), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n876), .A2(new_n878), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT52), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT117), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n869), .A2(KEYINPUT52), .A3(new_n724), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n876), .A2(new_n878), .A3(KEYINPUT115), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n871), .B1(new_n699), .B2(new_n756), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT117), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT52), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n869), .A2(new_n724), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n699), .A2(new_n756), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n890), .A2(new_n891), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n886), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n387), .A2(new_n463), .ZN(new_n898));
  NOR4_X1   g712(.A1(new_n813), .A2(new_n680), .A3(new_n898), .A4(new_n687), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n330), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n900), .B1(new_n778), .B2(new_n689), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n475), .B1(new_n671), .B2(new_n650), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n633), .B2(new_n634), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n639), .A2(new_n904), .A3(new_n539), .A4(new_n583), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n636), .A2(new_n905), .A3(new_n682), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n840), .A2(KEYINPUT114), .A3(new_n783), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT114), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n784), .B2(new_n839), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n787), .A2(new_n902), .A3(new_n906), .A4(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n744), .B(new_n751), .C1(new_n729), .C2(new_n738), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n735), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT53), .B1(new_n897), .B2(new_n915), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n330), .A2(new_n635), .B1(new_n681), .B2(new_n639), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n910), .A2(new_n905), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n901), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT52), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n895), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n912), .B1(new_n734), .B2(new_n730), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n919), .A2(new_n921), .A3(new_n922), .A4(new_n787), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT53), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT54), .B1(new_n916), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n911), .A2(new_n914), .A3(new_n924), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n897), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT54), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n923), .A2(new_n924), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  OAI22_X1  g746(.A1(new_n858), .A2(new_n932), .B1(G952), .B2(G953), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n830), .B(KEYINPUT49), .ZN(new_n934));
  AND4_X1   g748(.A1(new_n477), .A2(new_n792), .A3(new_n583), .A4(new_n631), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n833), .A2(new_n705), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n936), .ZN(G75));
  NOR2_X1   g751(.A1(new_n258), .A2(G952), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n928), .A2(new_n930), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(G210), .A3(G902), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n621), .A2(new_n624), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(new_n622), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT55), .Z(new_n945));
  OR2_X1    g759(.A1(new_n945), .A2(KEYINPUT56), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n939), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT119), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT56), .B1(new_n941), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n948), .B2(new_n941), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n947), .B1(new_n950), .B2(new_n945), .ZN(G51));
  INV_X1    g765(.A(new_n940), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n952), .A2(new_n379), .A3(new_n804), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n773), .B(KEYINPUT57), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n929), .B1(new_n928), .B2(new_n930), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n533), .A2(new_n535), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT120), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n953), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n957), .A2(KEYINPUT120), .A3(new_n958), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n938), .B1(new_n961), .B2(new_n962), .ZN(G54));
  NAND4_X1  g777(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n964));
  INV_X1    g778(.A(new_n457), .ZN(new_n965));
  OAI21_X1  g779(.A(KEYINPUT121), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n938), .B1(new_n964), .B2(new_n965), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n964), .A2(KEYINPUT121), .A3(new_n965), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(G60));
  OR2_X1    g784(.A1(new_n955), .A2(new_n956), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n644), .A2(new_n645), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(G478), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT59), .Z(new_n975));
  NOR2_X1   g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n938), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n975), .B1(new_n926), .B2(new_n931), .ZN(new_n978));
  OAI21_X1  g792(.A(KEYINPUT122), .B1(new_n978), .B2(new_n972), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n978), .A2(KEYINPUT122), .A3(new_n972), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(G63));
  NAND2_X1  g796(.A1(G217), .A2(G902), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT60), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n952), .A2(new_n676), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n570), .B1(new_n952), .B2(new_n984), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n985), .A2(new_n939), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT61), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n985), .A2(new_n986), .A3(KEYINPUT61), .A4(new_n939), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(G66));
  INV_X1    g805(.A(new_n602), .ZN(new_n992));
  OAI21_X1  g806(.A(G953), .B1(new_n992), .B2(new_n472), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n922), .A2(new_n906), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n993), .B1(new_n994), .B2(G953), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n943), .B1(G898), .B2(new_n258), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT123), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n995), .B(new_n997), .ZN(G69));
  AND2_X1   g812(.A1(new_n298), .A2(new_n288), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n449), .A2(new_n450), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n812), .A2(new_n881), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n851), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n821), .A2(new_n790), .A3(new_n815), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n787), .ZN(new_n1005));
  INV_X1    g819(.A(new_n724), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1006), .B1(new_n879), .B2(new_n872), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n1004), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n1009), .A2(G953), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n685), .A2(G953), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1011), .B(KEYINPUT125), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1001), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1001), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n718), .A2(new_n1007), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1015), .A2(KEYINPUT62), .ZN(new_n1016));
  INV_X1    g830(.A(new_n715), .ZN(new_n1017));
  OR2_X1    g831(.A1(new_n671), .A2(new_n650), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n732), .A2(new_n1017), .A3(new_n759), .A4(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n821), .A2(new_n815), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  AND3_X1   g835(.A1(new_n1015), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1022));
  AOI21_X1  g836(.A(KEYINPUT124), .B1(new_n1015), .B2(KEYINPUT62), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1014), .B1(new_n1024), .B2(new_n258), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n258), .B1(G227), .B2(G900), .ZN(new_n1026));
  OR3_X1    g840(.A1(new_n1013), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1026), .B1(new_n1013), .B2(new_n1025), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(new_n1028), .ZN(G72));
  XNOR2_X1  g843(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n838), .A2(new_n379), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1030), .B(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1033), .B1(new_n1009), .B2(new_n994), .ZN(new_n1034));
  INV_X1    g848(.A(new_n313), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(new_n269), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n939), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g851(.A(new_n1021), .B(new_n994), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1038));
  AOI211_X1 g852(.A(new_n269), .B(new_n1035), .C1(new_n1038), .C2(new_n1032), .ZN(new_n1039));
  OR2_X1    g853(.A1(new_n916), .A2(new_n925), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1033), .B1(new_n314), .B2(new_n308), .ZN(new_n1041));
  XNOR2_X1  g855(.A(new_n1041), .B(KEYINPUT127), .ZN(new_n1042));
  AOI211_X1 g856(.A(new_n1037), .B(new_n1039), .C1(new_n1040), .C2(new_n1042), .ZN(G57));
endmodule


