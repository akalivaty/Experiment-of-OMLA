//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n189), .A2(KEYINPUT79), .A3(G104), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT3), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT80), .B(G101), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n189), .A2(G104), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n195), .A2(new_n189), .A3(KEYINPUT79), .A4(G104), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n191), .A2(new_n192), .A3(new_n194), .A4(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n189), .A2(G104), .ZN(new_n198));
  OAI21_X1  g012(.A(G101), .B1(new_n198), .B2(new_n193), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT64), .B1(new_n204), .B2(G146), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(G146), .ZN(new_n206));
  OAI211_X1 g020(.A(G128), .B(new_n203), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(G143), .B2(new_n202), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OR2_X1    g026(.A1(new_n205), .A2(new_n206), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(new_n203), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n200), .B1(new_n208), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n202), .A2(G143), .ZN(new_n216));
  OAI22_X1  g030(.A1(new_n210), .A2(new_n211), .B1(new_n206), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n215), .B1(new_n218), .B2(new_n200), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT11), .ZN(new_n220));
  INV_X1    g034(.A(G134), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G137), .ZN(new_n222));
  INV_X1    g036(.A(G137), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT11), .A3(G134), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(G137), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n222), .A2(new_n224), .A3(new_n228), .A4(new_n225), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n219), .A2(KEYINPUT12), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT12), .B1(new_n219), .B2(new_n230), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n197), .A2(KEYINPUT10), .A3(new_n199), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n215), .A2(new_n234), .B1(new_n218), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n197), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n191), .A2(new_n194), .A3(new_n196), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT81), .A3(G101), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n238), .A2(KEYINPUT81), .A3(KEYINPUT4), .A4(G101), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n245), .B(new_n203), .C1(new_n205), .C2(new_n206), .ZN(new_n246));
  OR2_X1    g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n244), .B(new_n247), .C1(new_n206), .C2(new_n216), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n246), .A2(new_n248), .A3(KEYINPUT69), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT69), .B1(new_n246), .B2(new_n248), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n243), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n236), .A2(new_n252), .A3(new_n229), .A4(new_n227), .ZN(new_n253));
  INV_X1    g067(.A(G953), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT70), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G227), .ZN(new_n259));
  XNOR2_X1  g073(.A(G110), .B(G140), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n259), .B(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n253), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n233), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n236), .A2(new_n252), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n230), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n261), .B1(new_n265), .B2(new_n253), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n187), .B(new_n188), .C1(new_n263), .C2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n187), .A2(new_n188), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n253), .B1(new_n231), .B2(new_n232), .ZN(new_n270));
  INV_X1    g084(.A(new_n261), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n265), .A2(new_n253), .A3(new_n261), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n267), .B(new_n269), .C1(new_n187), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G221), .ZN(new_n276));
  XOR2_X1   g090(.A(KEYINPUT9), .B(G234), .Z(new_n277));
  AOI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(new_n188), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT90), .ZN(new_n281));
  NOR2_X1   g095(.A1(G475), .A2(G902), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(KEYINPUT89), .ZN(new_n284));
  INV_X1    g098(.A(G237), .ZN(new_n285));
  AND4_X1   g099(.A1(G143), .A2(new_n258), .A3(G214), .A4(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(G237), .B1(new_n255), .B2(new_n257), .ZN(new_n287));
  AOI21_X1  g101(.A(G143), .B1(new_n287), .B2(G214), .ZN(new_n288));
  OAI21_X1  g102(.A(G131), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT17), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n258), .A2(G214), .A3(new_n285), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n204), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n287), .A2(G143), .A3(G214), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n228), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n289), .A2(new_n290), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(G125), .B(G140), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT16), .ZN(new_n297));
  INV_X1    g111(.A(G140), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G125), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n297), .B1(KEYINPUT16), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n202), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n297), .B(G146), .C1(KEYINPUT16), .C2(new_n299), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(KEYINPUT17), .B(G131), .C1(new_n286), .C2(new_n288), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n295), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(KEYINPUT18), .B(G131), .C1(new_n286), .C2(new_n288), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT18), .A2(G131), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n292), .A2(new_n293), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G125), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n299), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G146), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n296), .A2(new_n202), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n306), .A2(new_n308), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(G113), .B(G122), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(G104), .ZN(new_n317));
  XOR2_X1   g131(.A(new_n317), .B(KEYINPUT88), .Z(new_n318));
  NAND3_X1  g132(.A1(new_n305), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n306), .A2(new_n308), .A3(new_n314), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n311), .A2(KEYINPUT19), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT19), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n296), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n302), .B1(G146), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n289), .B2(new_n294), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n317), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  AOI211_X1 g141(.A(KEYINPUT20), .B(new_n284), .C1(new_n319), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n283), .A2(KEYINPUT89), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n319), .A2(new_n327), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n282), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n328), .A2(new_n329), .B1(new_n331), .B2(KEYINPUT20), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n305), .A2(new_n315), .A3(new_n318), .ZN(new_n333));
  INV_X1    g147(.A(new_n317), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n305), .B2(new_n315), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n188), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G475), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n281), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n254), .A2(G952), .ZN(new_n340));
  INV_X1    g154(.A(G234), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(new_n285), .ZN(new_n342));
  XOR2_X1   g156(.A(new_n342), .B(KEYINPUT95), .Z(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n258), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n345), .B(G902), .C1(new_n341), .C2(new_n285), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT96), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT21), .B(G898), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(KEYINPUT97), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n344), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT20), .ZN(new_n352));
  INV_X1    g166(.A(new_n284), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n330), .A2(new_n352), .A3(new_n329), .A4(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n283), .B1(new_n319), .B2(new_n327), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n354), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT90), .A3(new_n337), .ZN(new_n357));
  INV_X1    g171(.A(G478), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(KEYINPUT15), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n277), .A2(G217), .A3(new_n254), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n204), .A2(KEYINPUT13), .A3(G128), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT91), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n211), .A2(G143), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n204), .A2(KEYINPUT91), .A3(KEYINPUT13), .A4(G128), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT13), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n211), .B2(G143), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n363), .A2(new_n364), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT92), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(G134), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(G128), .B(G143), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n221), .ZN(new_n373));
  INV_X1    g187(.A(G116), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G122), .ZN(new_n375));
  INV_X1    g189(.A(G122), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G116), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n378), .A2(new_n189), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n189), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n373), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n369), .B1(new_n368), .B2(G134), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n371), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT93), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(new_n375), .B2(KEYINPUT14), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT14), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n386), .A2(new_n374), .A3(KEYINPUT93), .A4(G122), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n375), .A2(KEYINPUT14), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n385), .A2(new_n377), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G107), .ZN(new_n390));
  INV_X1    g204(.A(new_n379), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n372), .B(new_n221), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n360), .B1(new_n383), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n360), .ZN(new_n396));
  INV_X1    g210(.A(new_n382), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n370), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n393), .B(new_n396), .C1(new_n398), .C2(new_n381), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n359), .B1(new_n400), .B2(G902), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n395), .A2(new_n399), .ZN(new_n402));
  INV_X1    g216(.A(new_n359), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n188), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n401), .A2(KEYINPUT94), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT94), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n403), .B1(new_n402), .B2(new_n188), .ZN(new_n407));
  AOI211_X1 g221(.A(G902), .B(new_n359), .C1(new_n395), .C2(new_n399), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n339), .A2(new_n351), .A3(new_n357), .A4(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n280), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT87), .ZN(new_n413));
  OAI21_X1  g227(.A(G210), .B1(G237), .B2(G902), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(KEYINPUT86), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT66), .B1(new_n374), .B2(G119), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT66), .ZN(new_n417));
  INV_X1    g231(.A(G119), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(G116), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g234(.A1(KEYINPUT2), .A2(G113), .ZN(new_n421));
  NOR2_X1   g235(.A1(KEYINPUT2), .A2(G113), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT67), .B1(new_n418), .B2(G116), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT67), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n374), .A3(G119), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n420), .A2(new_n423), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT68), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n424), .A2(new_n426), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n430), .A2(KEYINPUT68), .A3(new_n423), .A4(new_n420), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT5), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n418), .A3(G116), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n420), .ZN(new_n435));
  OAI211_X1 g249(.A(G113), .B(new_n434), .C1(new_n435), .C2(new_n433), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n436), .A3(new_n200), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G122), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n239), .A2(new_n240), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n439), .A2(new_n197), .A3(new_n242), .ZN(new_n440));
  INV_X1    g254(.A(new_n423), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n429), .A2(new_n431), .B1(new_n441), .B2(new_n435), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n437), .B(new_n438), .C1(new_n440), .C2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n438), .B(KEYINPUT8), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n432), .A2(new_n200), .A3(new_n436), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n200), .B1(new_n432), .B2(new_n436), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n309), .B1(new_n246), .B2(new_n248), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT84), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT7), .ZN(new_n450));
  INV_X1    g264(.A(G224), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(G953), .ZN(new_n452));
  OAI22_X1  g266(.A1(new_n448), .A2(new_n449), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n217), .B(new_n309), .C1(new_n207), .C2(KEYINPUT1), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n246), .A2(new_n248), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(new_n309), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n453), .B(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n443), .A2(new_n447), .A3(new_n457), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n458), .A2(KEYINPUT85), .A3(new_n188), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT85), .B1(new_n458), .B2(new_n188), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n456), .B(new_n452), .Z(new_n462));
  INV_X1    g276(.A(new_n438), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n435), .A2(new_n441), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n241), .A2(new_n242), .B1(new_n432), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n463), .B1(new_n465), .B2(new_n445), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(KEYINPUT6), .A3(new_n443), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n468), .B(new_n463), .C1(new_n465), .C2(new_n445), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(KEYINPUT83), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT83), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n466), .A2(new_n443), .A3(new_n471), .A4(KEYINPUT6), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n462), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n415), .B1(new_n461), .B2(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n466), .A2(KEYINPUT6), .A3(new_n443), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n469), .A2(KEYINPUT83), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n462), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n458), .A2(new_n188), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n458), .A2(KEYINPUT85), .A3(new_n188), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n415), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n479), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n474), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G214), .B1(G237), .B2(G902), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n413), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n488), .ZN(new_n490));
  AOI211_X1 g304(.A(KEYINPUT87), .B(new_n490), .C1(new_n474), .C2(new_n486), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n412), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT98), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G217), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n495), .B1(G234), .B2(new_n188), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT24), .B(G110), .Z(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT76), .ZN(new_n498));
  XNOR2_X1  g312(.A(G119), .B(G128), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT77), .B1(new_n418), .B2(G128), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n500), .A2(KEYINPUT23), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(KEYINPUT23), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n501), .B(new_n502), .C1(G119), .C2(new_n211), .ZN(new_n503));
  OAI22_X1  g317(.A1(new_n498), .A2(new_n499), .B1(new_n503), .B2(G110), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n302), .A3(new_n313), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n301), .A2(new_n302), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(G110), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n498), .A2(new_n499), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n258), .A2(G221), .A3(G234), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT78), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT22), .B(G137), .Z(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n510), .A2(new_n514), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT25), .B1(new_n517), .B2(new_n188), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT25), .ZN(new_n519));
  AOI211_X1 g333(.A(new_n519), .B(G902), .C1(new_n515), .C2(new_n516), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n496), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n496), .A2(G902), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT74), .B(KEYINPUT32), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n230), .B1(new_n249), .B2(new_n250), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n221), .A2(G137), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT65), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT65), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n225), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n528), .B(G131), .C1(new_n530), .C2(new_n527), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n218), .A2(new_n229), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n526), .A2(new_n442), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT28), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n442), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n455), .A2(new_n230), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n526), .A2(new_n442), .A3(KEYINPUT28), .A4(new_n532), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n535), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n258), .A2(G210), .A3(new_n285), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT26), .B(G101), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n538), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n526), .A2(KEYINPUT30), .A3(new_n532), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n550), .A3(new_n536), .ZN(new_n551));
  XOR2_X1   g365(.A(new_n544), .B(new_n545), .Z(new_n552));
  INV_X1    g366(.A(KEYINPUT72), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n533), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT31), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n547), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n559));
  NOR2_X1   g373(.A1(G472), .A2(G902), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n559), .B1(new_n558), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n525), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n560), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n554), .A2(new_n555), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n554), .A2(new_n555), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n564), .B1(new_n567), .B2(new_n547), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT29), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n541), .A2(new_n552), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n551), .A2(new_n546), .A3(new_n533), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n569), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n526), .A2(new_n532), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n536), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(KEYINPUT75), .A3(new_n533), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT75), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n574), .A2(new_n577), .A3(new_n536), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n576), .A2(KEYINPUT28), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n535), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n552), .A2(KEYINPUT29), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n573), .B(new_n188), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n568), .A2(KEYINPUT32), .B1(new_n582), .B2(G472), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n524), .B1(new_n563), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n412), .B(KEYINPUT98), .C1(new_n489), .C2(new_n491), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n494), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n586), .B(new_n192), .Z(G3));
  INV_X1    g401(.A(new_n280), .ZN(new_n588));
  INV_X1    g402(.A(new_n524), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n558), .A2(new_n188), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(new_n561), .B2(new_n562), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT99), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n593), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT99), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n595), .A2(new_n588), .A3(new_n596), .A4(new_n589), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n414), .B1(new_n461), .B2(new_n473), .ZN(new_n600));
  INV_X1    g414(.A(new_n414), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n479), .A2(new_n484), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(new_n602), .A3(new_n488), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT100), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT100), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n600), .A2(new_n602), .A3(new_n605), .A4(new_n488), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n339), .A2(new_n357), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n400), .A2(KEYINPUT33), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n400), .A2(KEYINPUT33), .ZN(new_n610));
  OAI21_X1  g424(.A(G478), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n402), .A2(new_n358), .A3(new_n188), .ZN(new_n612));
  NAND2_X1  g426(.A1(G478), .A2(G902), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n350), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n599), .A2(new_n607), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT34), .B(G104), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  NAND2_X1  g433(.A1(new_n331), .A2(KEYINPUT20), .ZN(new_n620));
  OR2_X1    g434(.A1(new_n620), .A2(KEYINPUT101), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n330), .A2(new_n352), .A3(new_n282), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(KEYINPUT101), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n410), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n624), .A2(new_n351), .A3(new_n625), .A4(new_n337), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT102), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n599), .A2(new_n607), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT103), .B(KEYINPUT104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT36), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n514), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT105), .ZN(new_n636));
  OR2_X1    g450(.A1(new_n636), .A2(new_n510), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n510), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(new_n638), .A3(new_n522), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n521), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n633), .B1(new_n593), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n595), .A2(KEYINPUT106), .A3(new_n640), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n494), .A2(new_n585), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT37), .B(G110), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  INV_X1    g460(.A(G900), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n344), .B1(new_n347), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  AND4_X1   g463(.A1(new_n337), .A2(new_n624), .A3(new_n625), .A4(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n641), .B1(new_n563), .B2(new_n583), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n607), .A2(new_n588), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  XOR2_X1   g467(.A(new_n648), .B(KEYINPUT39), .Z(new_n654));
  NAND2_X1  g468(.A1(new_n588), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n487), .B(KEYINPUT38), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AOI221_X4 g472(.A(new_n281), .B1(new_n336), .B2(G475), .C1(new_n620), .C2(new_n354), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT90), .B1(new_n356), .B2(new_n337), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n625), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n656), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n568), .A2(KEYINPUT32), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n551), .A2(new_n533), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n552), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n576), .A2(new_n578), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n188), .B(new_n665), .C1(new_n666), .C2(new_n552), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G472), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n563), .A2(new_n663), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n641), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n490), .B1(new_n655), .B2(KEYINPUT40), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n662), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G143), .ZN(G45));
  NAND3_X1  g488(.A1(new_n608), .A2(new_n614), .A3(new_n649), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n607), .A2(new_n588), .A3(new_n651), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  OR2_X1    g492(.A1(new_n263), .A2(new_n266), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n187), .B1(new_n679), .B2(new_n188), .ZN(new_n680));
  INV_X1    g494(.A(new_n267), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n680), .A2(new_n278), .A3(new_n681), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n604), .A2(new_n606), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n584), .A3(new_n616), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n683), .A2(KEYINPUT107), .A3(new_n584), .A4(new_n616), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  NAND3_X1  g504(.A1(new_n627), .A2(new_n584), .A3(new_n683), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT108), .B(G116), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G18));
  INV_X1    g507(.A(new_n411), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n607), .A2(new_n694), .A3(new_n651), .A4(new_n682), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G119), .ZN(G21));
  AOI22_X1  g510(.A1(new_n565), .A2(new_n566), .B1(new_n580), .B2(new_n546), .ZN(new_n697));
  OR2_X1    g511(.A1(new_n697), .A2(new_n564), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n589), .A2(new_n592), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n682), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n350), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT109), .B1(new_n608), .B2(new_n625), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n704));
  AOI211_X1 g518(.A(new_n704), .B(new_n410), .C1(new_n339), .C2(new_n357), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n702), .B1(new_n607), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n661), .A2(new_n704), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n625), .B(KEYINPUT109), .C1(new_n659), .C2(new_n660), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(new_n604), .A3(new_n606), .A4(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(KEYINPUT110), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n699), .B(new_n701), .C1(new_n707), .C2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  NAND3_X1  g527(.A1(new_n640), .A2(new_n698), .A3(new_n592), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n675), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n683), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G125), .ZN(G27));
  NOR2_X1   g531(.A1(new_n487), .A2(new_n490), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n584), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT42), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n280), .B(KEYINPUT111), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n719), .A2(new_n720), .A3(new_n676), .A4(new_n721), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n568), .A2(KEYINPUT32), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n524), .B1(new_n583), .B2(new_n723), .ZN(new_n724));
  AND4_X1   g538(.A1(new_n676), .A2(new_n721), .A3(new_n724), .A4(new_n718), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n722), .B1(new_n725), .B2(new_n720), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n228), .ZN(G33));
  AND3_X1   g541(.A1(new_n719), .A2(new_n650), .A3(new_n721), .ZN(new_n728));
  XOR2_X1   g542(.A(KEYINPUT112), .B(G134), .Z(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G36));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n274), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n272), .A2(KEYINPUT45), .A3(new_n273), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(G469), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n268), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n738), .A2(KEYINPUT46), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n681), .B1(new_n738), .B2(KEYINPUT46), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n278), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n654), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT114), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n614), .A2(new_n339), .A3(new_n357), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT43), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(KEYINPUT43), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n593), .A3(new_n640), .A4(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n718), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n743), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g567(.A(KEYINPUT115), .B(G137), .Z(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G39));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n739), .A2(new_n740), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n756), .B1(new_n757), .B2(new_n278), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n741), .A2(KEYINPUT47), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n761));
  INV_X1    g575(.A(new_n718), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n563), .A2(new_n583), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n762), .A2(new_n763), .A3(new_n589), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n760), .A2(new_n761), .A3(new_n676), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n741), .A2(KEYINPUT47), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n756), .B(new_n278), .C1(new_n739), .C2(new_n740), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n676), .B(new_n764), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT116), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n680), .A2(new_n681), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n758), .B(new_n759), .C1(new_n279), .C2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n745), .A2(new_n699), .A3(new_n344), .A4(new_n746), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n775), .A2(new_n718), .A3(new_n777), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n776), .A2(new_n488), .A3(new_n657), .A4(new_n700), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n745), .A2(new_n746), .ZN(new_n783));
  INV_X1    g597(.A(new_n714), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n762), .A2(new_n700), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n344), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n781), .A2(new_n782), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n669), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n785), .A2(new_n589), .A3(new_n788), .A4(new_n344), .ZN(new_n789));
  OR3_X1    g603(.A1(new_n789), .A2(new_n608), .A3(new_n614), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n772), .B1(new_n778), .B2(new_n791), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n789), .A2(new_n615), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n775), .A2(new_n718), .A3(new_n777), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n794), .A2(KEYINPUT51), .A3(new_n787), .A4(new_n790), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n792), .A2(new_n340), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n783), .A2(new_n344), .A3(new_n724), .A4(new_n785), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n797), .B(KEYINPUT48), .Z(new_n798));
  NOR2_X1   g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n652), .A2(new_n677), .A3(new_n716), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n280), .A2(new_n648), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n671), .B(new_n801), .C1(new_n707), .C2(new_n711), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n800), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n803), .B1(new_n800), .B2(new_n802), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n688), .A2(new_n712), .A3(new_n691), .A4(new_n695), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n726), .ZN(new_n808));
  INV_X1    g622(.A(new_n489), .ZN(new_n809));
  INV_X1    g623(.A(new_n491), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n350), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n407), .A2(new_n408), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n608), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n811), .A2(new_n594), .A3(new_n597), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n644), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n615), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n811), .A2(new_n594), .A3(new_n597), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n586), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT117), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n586), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n815), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n721), .A2(new_n592), .A3(new_n676), .A4(new_n698), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n338), .A2(new_n648), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n624), .A2(new_n812), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n280), .B1(new_n825), .B2(KEYINPUT118), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n826), .B(new_n763), .C1(KEYINPUT118), .C2(new_n825), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n641), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n728), .B1(new_n828), .B2(new_n718), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n806), .A2(new_n808), .A3(new_n822), .A4(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n815), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n586), .A2(new_n817), .A3(new_n820), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n820), .B1(new_n586), .B2(new_n817), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n829), .B(new_n833), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n801), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n607), .A2(new_n706), .A3(new_n702), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n710), .A2(KEYINPUT110), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n670), .B(new_n837), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n652), .A2(new_n677), .A3(new_n716), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT52), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n800), .A2(new_n802), .A3(new_n803), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n836), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT53), .B1(new_n845), .B2(new_n808), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT54), .B1(new_n832), .B2(new_n846), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n807), .A2(KEYINPUT119), .A3(new_n726), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT119), .B1(new_n807), .B2(new_n726), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n845), .A2(KEYINPUT53), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n830), .A2(new_n831), .ZN(new_n851));
  XNOR2_X1  g665(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT121), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n799), .A2(new_n847), .A3(new_n853), .A4(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n777), .A2(new_n683), .ZN(new_n858));
  OAI22_X1  g672(.A1(new_n857), .A2(new_n858), .B1(G952), .B2(G953), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n589), .B1(new_n774), .B2(KEYINPUT49), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(KEYINPUT49), .B2(new_n774), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n744), .A2(new_n490), .A3(new_n278), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(new_n658), .A3(new_n788), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n863), .ZN(G75));
  AOI21_X1  g678(.A(new_n188), .B1(new_n850), .B2(new_n851), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(G210), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT56), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n477), .B(new_n462), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT55), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n869), .B1(new_n866), .B2(new_n867), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n258), .A2(G952), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(G51));
  NAND2_X1  g687(.A1(new_n269), .A2(KEYINPUT57), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n269), .A2(KEYINPUT57), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n852), .B1(new_n850), .B2(new_n851), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n874), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n679), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n865), .A2(new_n737), .A3(new_n736), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n872), .B1(new_n879), .B2(new_n880), .ZN(G54));
  NAND3_X1  g695(.A1(new_n865), .A2(KEYINPUT58), .A3(G475), .ZN(new_n882));
  INV_X1    g696(.A(new_n330), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n884), .A2(new_n885), .A3(new_n872), .ZN(G60));
  NOR2_X1   g700(.A1(new_n609), .A2(new_n610), .ZN(new_n887));
  XNOR2_X1  g701(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(new_n613), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n887), .B(new_n889), .C1(new_n876), .C2(new_n877), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n891));
  INV_X1    g705(.A(new_n872), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n891), .B1(new_n890), .B2(new_n892), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n856), .A2(new_n847), .A3(new_n853), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n887), .B1(new_n895), .B2(new_n889), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(G63));
  XNOR2_X1  g711(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n850), .A2(new_n851), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n637), .A2(new_n638), .ZN(new_n900));
  NAND2_X1  g714(.A1(G217), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT60), .Z(new_n902));
  NAND3_X1  g716(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n892), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n517), .B1(new_n899), .B2(new_n902), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n898), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT125), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n904), .A2(new_n905), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT61), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n910), .B(new_n898), .C1(new_n904), .C2(new_n905), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n907), .A2(new_n909), .A3(new_n911), .ZN(G66));
  INV_X1    g726(.A(new_n822), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n913), .A2(new_n807), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n349), .A2(new_n451), .ZN(new_n915));
  AOI22_X1  g729(.A1(new_n914), .A2(new_n258), .B1(G953), .B2(new_n915), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n470), .B(new_n472), .C1(G898), .C2(new_n258), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n916), .B(new_n917), .Z(G69));
  NOR2_X1   g732(.A1(new_n258), .A2(G900), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n549), .A2(new_n550), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT126), .Z(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n324), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n724), .B1(new_n707), .B2(new_n711), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n751), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n726), .B1(new_n743), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n728), .A2(new_n841), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n770), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI211_X1 g741(.A(new_n919), .B(new_n922), .C1(new_n927), .C2(new_n258), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n673), .A2(new_n800), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT62), .Z(new_n930));
  INV_X1    g744(.A(new_n813), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n655), .B1(new_n615), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n719), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n770), .A2(new_n930), .A3(new_n753), .A4(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n934), .A2(new_n258), .A3(new_n922), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT127), .B1(new_n928), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n922), .B1(new_n927), .B2(new_n258), .ZN(new_n937));
  INV_X1    g751(.A(new_n919), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n934), .A2(new_n258), .A3(new_n922), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(G227), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n345), .B1(new_n943), .B2(new_n647), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n936), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n944), .B1(new_n936), .B2(new_n942), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(G72));
  OR2_X1    g761(.A1(new_n832), .A2(new_n846), .ZN(new_n948));
  NAND2_X1  g762(.A1(G472), .A2(G902), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT63), .Z(new_n950));
  NAND4_X1  g764(.A1(new_n948), .A2(new_n571), .A3(new_n665), .A4(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n950), .B1(new_n934), .B2(new_n914), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n952), .A2(new_n552), .A3(new_n664), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n950), .B1(new_n927), .B2(new_n914), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n872), .B1(new_n954), .B2(new_n572), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n951), .A2(new_n953), .A3(new_n955), .ZN(G57));
endmodule


