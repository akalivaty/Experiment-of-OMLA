//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G116), .ZN(new_n213));
  INV_X1    g0013(.A(G270), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AND2_X1   g0015(.A1(G68), .A2(G238), .ZN(new_n216));
  AND2_X1   g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  NOR4_X1   g0017(.A1(new_n212), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n203), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n207), .B(new_n228), .C1(new_n231), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n214), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  OAI211_X1 g0057(.A(G1), .B(G13), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n252), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n260));
  OR2_X1    g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n260), .B1(new_n263), .B2(G77), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G222), .ZN(new_n266));
  INV_X1    g0066(.A(G223), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(new_n265), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n255), .B1(new_n220), .B2(new_n259), .C1(new_n264), .C2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G169), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G179), .B2(new_n273), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n229), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n251), .A2(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G50), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(G50), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G150), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR3_X1   g0089(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n287), .A2(new_n289), .B1(new_n290), .B2(new_n230), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n224), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(KEYINPUT66), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n256), .A2(G20), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n283), .B(new_n286), .C1(new_n296), .C2(new_n279), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n276), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G238), .A2(G1698), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n263), .B(new_n301), .C1(new_n225), .C2(G1698), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n302), .B(new_n260), .C1(G107), .C2(new_n263), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n303), .B(new_n255), .C1(new_n222), .C2(new_n259), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n274), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G20), .A2(G77), .ZN(new_n306));
  XOR2_X1   g0106(.A(KEYINPUT15), .B(G87), .Z(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n295), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n306), .B1(new_n293), .B2(new_n289), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n284), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n310), .A2(new_n278), .B1(new_n221), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n282), .A2(G77), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n305), .B(new_n314), .C1(G179), .C2(new_n304), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT68), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n317), .A2(KEYINPUT9), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(KEYINPUT9), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n297), .A2(KEYINPUT67), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n297), .A2(KEYINPUT67), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n318), .B(new_n319), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n291), .ZN(new_n323));
  INV_X1    g0123(.A(new_n294), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n309), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n285), .B1(new_n325), .B2(new_n278), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT67), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(new_n283), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n297), .A2(KEYINPUT67), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n328), .A2(new_n317), .A3(KEYINPUT9), .A4(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT69), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n273), .A2(new_n332), .A3(G200), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n332), .B1(new_n273), .B2(G200), .ZN(new_n334));
  INV_X1    g0134(.A(G190), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n333), .A2(new_n334), .B1(new_n335), .B2(new_n273), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n316), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  AOI211_X1 g0138(.A(KEYINPUT10), .B(new_n336), .C1(new_n322), .C2(new_n330), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n300), .B(new_n315), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT16), .ZN(new_n341));
  INV_X1    g0141(.A(G68), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n261), .A2(new_n230), .A3(new_n262), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT7), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n230), .A4(new_n262), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n342), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n224), .A2(new_n342), .ZN(new_n348));
  NOR2_X1   g0148(.A1(G58), .A2(G68), .ZN(new_n349));
  OAI21_X1  g0149(.A(G20), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n288), .A2(G159), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n341), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT7), .B1(new_n271), .B2(new_n230), .ZN(new_n354));
  INV_X1    g0154(.A(new_n346), .ZN(new_n355));
  OAI21_X1  g0155(.A(G68), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n352), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(KEYINPUT16), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(new_n358), .A3(new_n278), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n324), .A2(new_n284), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n294), .A2(new_n281), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G179), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n255), .B1(new_n259), .B2(new_n225), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT71), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n267), .A2(new_n265), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n220), .A2(G1698), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n368), .B(new_n369), .C1(new_n269), .C2(new_n270), .ZN(new_n370));
  AND3_X1   g0170(.A1(KEYINPUT70), .A2(G33), .A3(G87), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT70), .B1(G33), .B2(G87), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n367), .B1(new_n374), .B2(new_n260), .ZN(new_n375));
  AOI211_X1 g0175(.A(KEYINPUT71), .B(new_n258), .C1(new_n370), .C2(new_n373), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n364), .B(new_n366), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n258), .B1(new_n370), .B2(new_n373), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n274), .B1(new_n365), .B2(new_n378), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n363), .A2(new_n380), .A3(KEYINPUT18), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT18), .B1(new_n363), .B2(new_n380), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n359), .A2(new_n362), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n335), .B(new_n366), .C1(new_n375), .C2(new_n376), .ZN(new_n385));
  INV_X1    g0185(.A(G200), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n365), .B2(new_n378), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n384), .A2(KEYINPUT17), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n362), .A3(new_n359), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT17), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n383), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n314), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n304), .A2(G200), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n395), .B(new_n396), .C1(new_n335), .C2(new_n304), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT13), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n225), .A2(G1698), .ZN(new_n400));
  OAI221_X1 g0200(.A(new_n400), .B1(G226), .B2(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G97), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n254), .B1(new_n403), .B2(new_n260), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n258), .A2(G238), .A3(new_n252), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n399), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n258), .B1(new_n401), .B2(new_n402), .ZN(new_n408));
  NOR4_X1   g0208(.A1(new_n408), .A2(KEYINPUT13), .A3(new_n405), .A4(new_n254), .ZN(new_n409));
  OAI21_X1  g0209(.A(G169), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT14), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n407), .A2(new_n409), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G179), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(G169), .C1(new_n407), .C2(new_n409), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n411), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n309), .A2(new_n221), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n289), .A2(new_n219), .B1(new_n230), .B2(G68), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n278), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  XOR2_X1   g0219(.A(new_n419), .B(KEYINPUT11), .Z(new_n420));
  NOR2_X1   g0220(.A1(new_n281), .A2(new_n342), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n311), .A2(new_n342), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT12), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n420), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n416), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n412), .A2(G190), .ZN(new_n429));
  OAI21_X1  g0229(.A(G200), .B1(new_n407), .B2(new_n409), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n425), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NOR4_X1   g0232(.A1(new_n340), .A2(new_n398), .A3(new_n428), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT23), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n230), .B2(G107), .ZN(new_n435));
  INV_X1    g0235(.A(G107), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(KEYINPUT23), .A3(G20), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n295), .A2(G116), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n230), .B(G87), .C1(new_n269), .C2(new_n270), .ZN(new_n440));
  NAND2_X1  g0240(.A1(KEYINPUT81), .A2(KEYINPUT22), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n438), .B(new_n439), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OR2_X1    g0243(.A1(KEYINPUT81), .A2(KEYINPUT22), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(new_n444), .A3(new_n441), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(KEYINPUT24), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT24), .ZN(new_n447));
  INV_X1    g0247(.A(new_n445), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n447), .B1(new_n448), .B2(new_n442), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n278), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n251), .A2(G33), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n284), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(new_n278), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G107), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n284), .A2(G107), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n455), .B(KEYINPUT25), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n450), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  OR2_X1    g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  NAND2_X1  g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G1), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(G264), .B(new_n258), .C1(new_n460), .C2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n251), .A2(G45), .A3(G274), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n261), .A2(new_n262), .B1(new_n211), .B2(G1698), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n209), .A2(new_n265), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n467), .A2(new_n468), .B1(G33), .B2(G294), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n464), .B(new_n466), .C1(new_n469), .C2(new_n258), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n335), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n457), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(G200), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n470), .A2(G169), .ZN(new_n475));
  OAI221_X1 g0275(.A(new_n468), .B1(G257), .B2(new_n265), .C1(new_n269), .C2(new_n270), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G294), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n256), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n260), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n480), .A2(G179), .A3(new_n466), .A4(new_n464), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT82), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n475), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n482), .B1(new_n475), .B2(new_n481), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n457), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n474), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n345), .A2(new_n346), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT73), .B1(new_n487), .B2(G107), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT73), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n489), .B(new_n436), .C1(new_n345), .C2(new_n346), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492));
  AND2_X1   g0292(.A1(G97), .A2(G107), .ZN(new_n493));
  NOR2_X1   g0293(.A1(G97), .A2(G107), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n436), .A2(KEYINPUT6), .A3(G97), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n230), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n289), .A2(new_n221), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT72), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT72), .ZN(new_n500));
  INV_X1    g0300(.A(new_n498), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n436), .A2(KEYINPUT6), .A3(G97), .ZN(new_n502));
  XNOR2_X1  g0302(.A(G97), .B(G107), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(new_n492), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n500), .B(new_n501), .C1(new_n504), .C2(new_n230), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n279), .B1(new_n491), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n284), .A2(G97), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n453), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(new_n210), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT76), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(G107), .B1(new_n354), .B2(new_n355), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n489), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n487), .A2(KEYINPUT73), .A3(G107), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n514), .A2(new_n505), .A3(new_n499), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n278), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT76), .ZN(new_n518));
  INV_X1    g0318(.A(new_n511), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n512), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n222), .A2(G1698), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n269), .B2(new_n270), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT4), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n522), .B(KEYINPUT4), .C1(new_n270), .C2(new_n269), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G283), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT74), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT74), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(G33), .A3(G283), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(G250), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n525), .A2(new_n526), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n260), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n258), .A2(new_n458), .A3(new_n459), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n258), .A2(new_n463), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G257), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n534), .A2(new_n466), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(G179), .ZN(new_n540));
  AND4_X1   g0340(.A1(KEYINPUT75), .A2(new_n534), .A3(new_n466), .A4(new_n538), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n460), .A2(new_n465), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n533), .B2(new_n260), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT75), .B1(new_n543), .B2(new_n538), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n540), .B1(new_n545), .B2(new_n274), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT75), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n543), .A2(KEYINPUT75), .A3(new_n538), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(G190), .B1(G200), .B2(new_n539), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n507), .A2(new_n511), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n521), .A2(new_n546), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n214), .B1(new_n535), .B2(new_n536), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n265), .A2(G257), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G264), .A2(G1698), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n555), .B(new_n556), .C1(new_n269), .C2(new_n270), .ZN(new_n557));
  INV_X1    g0357(.A(G303), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n261), .A2(new_n558), .A3(new_n262), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n260), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT79), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT79), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n557), .A2(new_n559), .A3(new_n562), .A4(new_n260), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n554), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n274), .B1(new_n564), .B2(new_n466), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT20), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n230), .B1(new_n210), .B2(G33), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n530), .B2(new_n528), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n278), .B1(new_n230), .B2(G116), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n567), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n531), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n277), .A2(new_n229), .B1(G20), .B2(new_n213), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(KEYINPUT20), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n311), .A2(new_n213), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n452), .A2(new_n213), .A3(new_n278), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AND4_X1   g0378(.A1(KEYINPUT80), .A2(new_n575), .A3(new_n576), .A4(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n577), .B1(new_n570), .B2(new_n574), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT80), .B1(new_n580), .B2(new_n576), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n565), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT21), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n561), .A2(new_n563), .ZN(new_n585));
  INV_X1    g0385(.A(new_n554), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n466), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(new_n364), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n581), .B2(new_n579), .ZN(new_n589));
  OAI211_X1 g0389(.A(KEYINPUT21), .B(new_n565), .C1(new_n579), .C2(new_n581), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n580), .A2(new_n576), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT80), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n587), .A2(G200), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n580), .A2(KEYINPUT80), .A3(new_n576), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n564), .A2(G190), .A3(new_n466), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n593), .A2(new_n594), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n584), .A2(new_n589), .A3(new_n590), .A4(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT78), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n258), .A2(new_n463), .A3(G250), .ZN(new_n600));
  XNOR2_X1  g0400(.A(new_n465), .B(KEYINPUT77), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n222), .A2(G1698), .ZN(new_n603));
  OAI221_X1 g0403(.A(new_n603), .B1(G238), .B2(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n604));
  NAND2_X1  g0404(.A1(G33), .A2(G116), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n600), .B(new_n602), .C1(new_n606), .C2(new_n258), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n599), .B1(new_n607), .B2(new_n335), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(G200), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n258), .B1(new_n604), .B2(new_n605), .ZN(new_n610));
  INV_X1    g0410(.A(new_n600), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n610), .A2(new_n611), .A3(new_n601), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(KEYINPUT78), .A3(G190), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n307), .A2(new_n284), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n452), .A2(new_n208), .A3(new_n278), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n263), .A2(new_n230), .A3(G68), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n494), .A2(new_n208), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n402), .A2(new_n230), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(KEYINPUT19), .A3(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n402), .A2(G20), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n616), .B(new_n619), .C1(KEYINPUT19), .C2(new_n620), .ZN(new_n621));
  AOI211_X1 g0421(.A(new_n614), .B(new_n615), .C1(new_n621), .C2(new_n278), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n608), .A2(new_n609), .A3(new_n613), .A4(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n614), .B1(new_n621), .B2(new_n278), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n308), .B2(new_n510), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n607), .A2(new_n274), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n612), .A2(new_n364), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n598), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n433), .A2(new_n486), .A3(new_n553), .A4(new_n630), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n631), .B(KEYINPUT83), .ZN(G372));
  NAND2_X1  g0432(.A1(new_n609), .A2(new_n622), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n633), .A2(KEYINPUT84), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n633), .A2(KEYINPUT84), .B1(G190), .B2(new_n612), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n475), .A2(new_n481), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n457), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n584), .A2(new_n589), .A3(new_n590), .A4(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n548), .A2(new_n274), .A3(new_n549), .ZN(new_n640));
  INV_X1    g0440(.A(new_n540), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n518), .B1(new_n517), .B2(new_n519), .ZN(new_n642));
  AOI211_X1 g0442(.A(KEYINPUT76), .B(new_n511), .C1(new_n516), .C2(new_n278), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n539), .A2(G200), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n552), .B(new_n645), .C1(new_n335), .C2(new_n545), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n639), .A2(new_n644), .A3(new_n474), .A4(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  INV_X1    g0448(.A(new_n552), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n640), .A2(KEYINPUT85), .A3(new_n641), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT85), .B1(new_n640), .B2(new_n641), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n648), .B(new_n649), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n636), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n623), .A2(new_n628), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n521), .A2(new_n655), .A3(new_n546), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT26), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n628), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n433), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n427), .B1(new_n432), .B2(new_n315), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n390), .B(KEYINPUT17), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n383), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n338), .A2(new_n339), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n300), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n659), .A2(new_n665), .ZN(G369));
  INV_X1    g0466(.A(G13), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G20), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n251), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n457), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n474), .A2(new_n485), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g0476(.A(new_n676), .B(KEYINPUT86), .Z(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n638), .ZN(new_n678));
  INV_X1    g0478(.A(new_n674), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n639), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n485), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n674), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G330), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n679), .B1(new_n593), .B2(new_n595), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n598), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n584), .A2(new_n589), .A3(new_n590), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n685), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n684), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n680), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n204), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G1), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n494), .A2(new_n208), .A3(new_n213), .ZN(new_n696));
  OAI22_X1  g0496(.A1(new_n695), .A2(new_n696), .B1(new_n232), .B2(new_n694), .ZN(new_n697));
  XOR2_X1   g0497(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n698));
  XNOR2_X1  g0498(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n628), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n644), .A2(new_n474), .A3(new_n646), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n584), .A2(new_n485), .A3(new_n589), .A4(new_n590), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n700), .B1(new_n634), .B2(new_n635), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n700), .B1(new_n702), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n640), .A2(new_n641), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT85), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n552), .B1(new_n710), .B2(new_n650), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n648), .B1(new_n634), .B2(new_n635), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n656), .A2(new_n648), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n674), .B1(new_n707), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n679), .B1(new_n654), .B2(new_n658), .ZN(new_n717));
  XOR2_X1   g0517(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n718));
  AOI22_X1  g0518(.A1(new_n716), .A2(KEYINPUT29), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n481), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n564), .A2(new_n612), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n720), .B(new_n721), .C1(new_n541), .C2(new_n544), .ZN(new_n722));
  XNOR2_X1  g0522(.A(KEYINPUT89), .B(KEYINPUT30), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT92), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n587), .A2(KEYINPUT90), .A3(new_n364), .A4(new_n607), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n470), .A3(new_n539), .ZN(new_n730));
  AOI21_X1  g0530(.A(G179), .B1(new_n564), .B2(new_n466), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT90), .B1(new_n731), .B2(new_n607), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n722), .A2(KEYINPUT92), .A3(new_n723), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n726), .A2(new_n728), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n674), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g0538(.A(KEYINPUT88), .B(KEYINPUT31), .Z(new_n739));
  OAI22_X1  g0539(.A1(new_n722), .A2(new_n727), .B1(new_n730), .B2(new_n732), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n722), .A2(new_n723), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n674), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT91), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n630), .A2(new_n553), .A3(new_n486), .A4(new_n679), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n728), .A2(new_n733), .A3(new_n724), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n746), .A2(KEYINPUT91), .A3(new_n674), .A4(new_n739), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n738), .A2(new_n744), .A3(new_n745), .A4(new_n747), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n748), .A2(G330), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n719), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n699), .B1(new_n750), .B2(G1), .ZN(G364));
  OAI21_X1  g0551(.A(G20), .B1(KEYINPUT94), .B2(G169), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(KEYINPUT94), .A2(G169), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n229), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n335), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G326), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n271), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n230), .B1(new_n761), .B2(G190), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n760), .B1(G294), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n756), .A2(G190), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT33), .B(G317), .Z(new_n767));
  NOR2_X1   g0567(.A1(new_n230), .A2(new_n335), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n386), .A2(G179), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n764), .B1(new_n766), .B2(new_n767), .C1(new_n558), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n364), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n768), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n230), .A2(G190), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n769), .ZN(new_n780));
  INV_X1    g0580(.A(G283), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n775), .A2(new_n779), .ZN(new_n783));
  INV_X1    g0583(.A(G311), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n779), .A2(new_n761), .ZN(new_n785));
  INV_X1    g0585(.A(G329), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n783), .A2(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR4_X1   g0587(.A1(new_n774), .A2(new_n778), .A3(new_n782), .A4(new_n787), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n766), .A2(new_n342), .B1(new_n762), .B2(new_n210), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT96), .ZN(new_n790));
  INV_X1    g0590(.A(new_n776), .ZN(new_n791));
  INV_X1    g0591(.A(new_n783), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G58), .A2(new_n791), .B1(new_n792), .B2(G77), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n773), .B2(new_n208), .ZN(new_n794));
  INV_X1    g0594(.A(new_n785), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G159), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT32), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n263), .B1(new_n780), .B2(new_n436), .C1(new_n758), .C2(new_n219), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n790), .A2(new_n794), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n755), .B1(new_n788), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n692), .A2(new_n271), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G355), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n246), .A2(new_n461), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n692), .A2(new_n263), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(G45), .B2(new_n232), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n802), .B1(G116), .B2(new_n204), .C1(new_n803), .C2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G13), .A2(G33), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G20), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n755), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n686), .A2(new_n688), .ZN(new_n812));
  INV_X1    g0612(.A(new_n809), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n800), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n695), .B1(G45), .B2(new_n668), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n815), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n812), .A2(G330), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(new_n689), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT97), .Z(G396));
  NOR2_X1   g0621(.A1(new_n755), .A2(new_n807), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT98), .Z(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n397), .B1(new_n395), .B2(new_n679), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n315), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n315), .A2(new_n674), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n815), .B1(G77), .B2(new_n824), .C1(new_n829), .C2(new_n808), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n773), .A2(new_n436), .B1(new_n210), .B2(new_n762), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n758), .A2(new_n558), .B1(new_n783), .B2(new_n213), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G283), .B2(new_n765), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT99), .Z(new_n834));
  AOI211_X1 g0634(.A(new_n831), .B(new_n834), .C1(G294), .C2(new_n791), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n795), .A2(G311), .ZN(new_n836));
  INV_X1    g0636(.A(new_n780), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(G87), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n835), .A2(new_n271), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT100), .Z(new_n840));
  AOI22_X1  g0640(.A1(new_n791), .A2(G143), .B1(G150), .B2(new_n765), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  INV_X1    g0642(.A(G159), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n841), .B1(new_n842), .B2(new_n758), .C1(new_n843), .C2(new_n783), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n845), .A2(KEYINPUT34), .B1(new_n846), .B2(new_n785), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G58), .B2(new_n763), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n837), .A2(G68), .ZN(new_n849));
  INV_X1    g0649(.A(new_n773), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(G50), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n271), .B1(new_n845), .B2(KEYINPUT34), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n848), .A2(new_n849), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n840), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n830), .B1(new_n854), .B2(new_n755), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n717), .A2(new_n828), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n679), .B(new_n829), .C1(new_n654), .C2(new_n658), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(new_n749), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n855), .B1(new_n859), .B2(new_n817), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G384));
  INV_X1    g0661(.A(new_n504), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n213), .B1(new_n862), .B2(KEYINPUT35), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n863), .B(new_n231), .C1(KEYINPUT35), .C2(new_n862), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT36), .ZN(new_n865));
  OAI21_X1  g0665(.A(G77), .B1(new_n224), .B2(new_n342), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n866), .A2(new_n232), .B1(G50), .B2(new_n342), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(G1), .A3(new_n667), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT101), .Z(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT106), .B1(new_n719), .B2(new_n433), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n717), .A2(new_n718), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n628), .B1(new_n701), .B2(new_n705), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n711), .A2(new_n712), .B1(new_n656), .B2(new_n648), .ZN(new_n874));
  OAI211_X1 g0674(.A(KEYINPUT29), .B(new_n679), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  AND4_X1   g0675(.A1(KEYINPUT106), .A2(new_n872), .A3(new_n433), .A4(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n665), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT37), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT103), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n881), .B(new_n341), .C1(new_n347), .C2(new_n352), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n341), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n356), .A2(new_n357), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n882), .A2(new_n278), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n362), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n384), .A2(new_n388), .B1(new_n886), .B2(new_n380), .ZN(new_n887));
  INV_X1    g0687(.A(new_n672), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n880), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n363), .A2(new_n380), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n363), .A2(new_n888), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n891), .A2(new_n892), .A3(new_n880), .A4(new_n390), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT18), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n363), .A2(new_n380), .A3(KEYINPUT18), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n889), .B1(new_n661), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n879), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n886), .A2(new_n380), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n889), .A2(new_n902), .A3(new_n390), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT37), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n893), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n905), .B(KEYINPUT38), .C1(new_n394), .C2(new_n889), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n901), .A2(KEYINPUT104), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT104), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n908), .B(new_n879), .C1(new_n895), .C2(new_n900), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n878), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n392), .B(new_n389), .C1(new_n381), .C2(new_n382), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT105), .ZN(new_n913));
  INV_X1    g0713(.A(new_n892), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n913), .B1(new_n912), .B2(new_n914), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n891), .A2(new_n892), .A3(new_n390), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n919), .A2(new_n893), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n906), .B1(new_n921), .B2(KEYINPUT38), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n878), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT102), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n416), .A2(new_n924), .A3(new_n426), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n924), .B1(new_n416), .B2(new_n426), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n925), .A2(new_n926), .A3(new_n674), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n911), .A2(new_n923), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n426), .A2(new_n674), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n431), .B(new_n929), .C1(new_n925), .C2(new_n926), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n428), .A2(new_n674), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n857), .B2(new_n827), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n909), .A3(new_n907), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n899), .A2(new_n888), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n928), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n877), .B(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n722), .A2(KEYINPUT92), .A3(new_n723), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT92), .B1(new_n722), .B2(new_n723), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n740), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n679), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n940), .B(new_n745), .C1(new_n945), .C2(new_n739), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n433), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(KEYINPUT107), .B(KEYINPUT108), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  INV_X1    g0750(.A(new_n917), .ZN(new_n951));
  INV_X1    g0751(.A(new_n920), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n952), .A3(new_n915), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n879), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n950), .B1(new_n954), .B2(new_n906), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n828), .B1(new_n930), .B2(new_n931), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n946), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n907), .A2(new_n946), .A3(new_n909), .A4(new_n956), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n955), .A2(new_n957), .B1(new_n958), .B2(new_n950), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n949), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(G330), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n939), .B(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n668), .A2(new_n251), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n870), .B1(new_n962), .B2(new_n963), .ZN(G367));
  OAI21_X1  g0764(.A(new_n553), .B1(new_n552), .B2(new_n679), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n687), .A2(new_n679), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n677), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT42), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n711), .A2(new_n674), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT109), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n971), .A2(new_n681), .B1(new_n546), .B2(new_n521), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n968), .B1(new_n972), .B2(new_n674), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n622), .A2(new_n679), .ZN(new_n974));
  MUX2_X1   g0774(.A(new_n704), .B(new_n700), .S(new_n974), .Z(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n690), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n971), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT110), .Z(new_n981));
  XNOR2_X1  g0781(.A(new_n979), .B(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n977), .B(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n693), .B(KEYINPUT41), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n680), .A2(new_n553), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(KEYINPUT111), .B2(KEYINPUT44), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT111), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT44), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(new_n680), .C2(new_n553), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n987), .B(new_n990), .C1(new_n988), .C2(new_n989), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n680), .A2(new_n970), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT45), .Z(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n978), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n991), .A2(new_n993), .A3(new_n690), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n683), .A2(new_n689), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n690), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n998), .A2(new_n687), .A3(new_n679), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n690), .A3(new_n966), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n750), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n995), .A2(new_n996), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n985), .B1(new_n1004), .B2(new_n750), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n251), .B1(new_n668), .B2(G45), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n983), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n763), .A2(G68), .B1(G159), .B2(new_n765), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1009), .B(new_n263), .C1(new_n773), .C2(new_n224), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G150), .A2(new_n791), .B1(new_n795), .B2(G137), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n219), .B2(new_n783), .C1(new_n221), .C2(new_n780), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(G143), .C2(new_n757), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n780), .A2(new_n210), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n762), .A2(new_n436), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n766), .A2(new_n478), .B1(new_n758), .B2(new_n784), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(G317), .C2(new_n795), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n792), .A2(G283), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n850), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT46), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n773), .B2(new_n213), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1014), .B(new_n1022), .C1(G303), .C2(new_n791), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1013), .B1(new_n1023), .B2(new_n271), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT47), .Z(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n755), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n975), .A2(new_n813), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n804), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n810), .B1(new_n204), .B2(new_n308), .C1(new_n242), .C2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1026), .A2(new_n815), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1008), .A2(new_n1030), .ZN(G387));
  OR2_X1    g0831(.A1(new_n1001), .A2(new_n750), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(new_n1002), .A3(new_n693), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1028), .B1(new_n239), .B2(G45), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n696), .B2(new_n801), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n293), .A2(G50), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT50), .Z(new_n1037));
  NOR2_X1   g0837(.A1(new_n342), .A2(new_n221), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1037), .A2(G45), .A3(new_n1038), .A4(new_n696), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1035), .A2(new_n1039), .B1(G107), .B2(new_n204), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n810), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n815), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n683), .A2(new_n813), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n758), .A2(new_n843), .B1(new_n780), .B2(new_n210), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n773), .A2(new_n221), .B1(new_n342), .B2(new_n783), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(G150), .C2(new_n795), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n294), .A2(new_n765), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n308), .A2(new_n762), .B1(new_n219), .B2(new_n776), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT112), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1046), .A2(new_n263), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n791), .A2(G317), .B1(G311), .B2(new_n765), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n558), .B2(new_n783), .C1(new_n777), .C2(new_n758), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT48), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n781), .B2(new_n762), .C1(new_n478), .C2(new_n773), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT49), .Z(new_n1055));
  OAI221_X1 g0855(.A(new_n271), .B1(new_n785), .B2(new_n759), .C1(new_n213), .C2(new_n780), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1050), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1042), .B(new_n1043), .C1(new_n755), .C2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1033), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(KEYINPUT113), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT113), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1033), .A2(new_n1062), .A3(new_n1059), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(G393));
  OR2_X1    g0864(.A1(new_n971), .A2(new_n813), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n791), .A2(G311), .B1(G317), .B2(new_n757), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT52), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1067), .A2(new_n263), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n781), .B2(new_n773), .C1(new_n478), .C2(new_n783), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n762), .A2(new_n213), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n766), .A2(new_n558), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n780), .A2(new_n436), .B1(new_n785), .B2(new_n777), .ZN(new_n1072));
  NOR4_X1   g0872(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n758), .A2(new_n287), .B1(new_n776), .B2(new_n843), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n795), .A2(G143), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1075), .A2(new_n263), .A3(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n762), .A2(new_n221), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n773), .A2(new_n342), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n838), .B1(new_n293), .B2(new_n783), .C1(new_n766), .C2(new_n219), .ZN(new_n1080));
  NOR4_X1   g0880(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n755), .B1(new_n1073), .B2(new_n1081), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n810), .B1(new_n210), .B2(new_n204), .C1(new_n249), .C2(new_n1028), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1065), .A2(new_n815), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n995), .A2(new_n996), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1084), .B1(new_n1085), .B2(new_n1006), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n694), .B1(new_n1085), .B2(new_n1002), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1086), .B1(new_n1004), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(G390));
  NOR3_X1   g0889(.A1(new_n895), .A2(new_n900), .A3(new_n879), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n953), .B2(new_n879), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1091), .A2(KEYINPUT39), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1092), .A2(new_n910), .B1(new_n934), .B2(new_n927), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT115), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n679), .B(new_n826), .C1(new_n873), .C2(new_n874), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n827), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1091), .B1(new_n1096), .B2(new_n932), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n927), .A2(KEYINPUT114), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT114), .ZN(new_n1099));
  NOR4_X1   g0899(.A1(new_n925), .A2(new_n926), .A3(new_n1099), .A4(new_n674), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1094), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n933), .B1(new_n1095), .B2(new_n827), .ZN(new_n1104));
  NOR4_X1   g0904(.A1(new_n1104), .A2(new_n1091), .A3(KEYINPUT115), .A4(new_n1101), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1093), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT116), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n946), .A2(G330), .A3(new_n956), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT117), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT117), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n946), .A2(new_n956), .A3(new_n1110), .A4(G330), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1107), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1106), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(KEYINPUT116), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n748), .A2(G330), .A3(new_n829), .A4(new_n932), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1093), .B1(new_n1114), .B2(new_n1115), .C1(new_n1103), .C2(new_n1105), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1096), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n946), .A2(G330), .A3(new_n829), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n933), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1120), .A2(new_n1115), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n744), .B1(new_n945), .B2(KEYINPUT31), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n745), .A2(new_n747), .ZN(new_n1123));
  OAI211_X1 g0923(.A(G330), .B(new_n829), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n933), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1125), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n857), .A2(new_n827), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1118), .A2(new_n1121), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(KEYINPUT118), .B1(new_n947), .B2(new_n684), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT118), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n433), .A2(new_n1130), .A3(new_n946), .A4(G330), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1132), .B(new_n665), .C1(new_n871), .C2(new_n876), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n694), .B1(new_n1117), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1134), .A2(new_n1113), .A3(new_n1116), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n807), .B1(new_n1092), .B2(new_n910), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT53), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n850), .B2(G150), .ZN(new_n1141));
  XOR2_X1   g0941(.A(KEYINPUT54), .B(G143), .Z(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n792), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n795), .A2(G125), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n763), .A2(G159), .B1(G128), .B2(new_n757), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n842), .B2(new_n766), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n271), .B(new_n1146), .C1(G132), .C2(new_n791), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n850), .A2(new_n1140), .A3(G150), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1143), .A2(new_n1144), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G50), .B2(new_n837), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1078), .B1(new_n850), .B2(G87), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1151), .B(new_n271), .C1(new_n781), .C2(new_n758), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n776), .A2(new_n213), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n785), .A2(new_n478), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n849), .B1(new_n210), .B2(new_n783), .C1(new_n766), .C2(new_n436), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n755), .B1(new_n1150), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n823), .A2(new_n324), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1139), .A2(new_n815), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n1117), .B2(new_n1006), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1138), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(G378));
  INV_X1    g0962(.A(KEYINPUT57), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1133), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1137), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT120), .ZN(new_n1166));
  XOR2_X1   g0966(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n663), .B2(new_n299), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n320), .A2(new_n321), .A3(new_n672), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1167), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n300), .B(new_n1170), .C1(new_n338), .C2(new_n339), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1169), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n959), .B2(G330), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n958), .A2(new_n950), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n922), .A2(KEYINPUT40), .A3(new_n956), .A4(new_n946), .ZN(new_n1177));
  AND4_X1   g0977(.A1(G330), .A2(new_n1176), .A3(new_n1174), .A4(new_n1177), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1175), .A2(new_n1178), .A3(new_n938), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(G330), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1174), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1176), .A2(new_n1174), .A3(new_n1177), .A4(G330), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n910), .B1(new_n878), .B2(new_n922), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n936), .B1(new_n1184), .B2(new_n927), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1182), .A2(new_n1183), .B1(new_n1185), .B2(new_n935), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1166), .B1(new_n1179), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n938), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1182), .A2(new_n1185), .A3(new_n935), .A4(new_n1183), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n1189), .A3(KEYINPUT120), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1163), .B1(new_n1165), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT121), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1137), .A2(new_n1164), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1179), .A2(new_n1186), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(KEYINPUT57), .A3(new_n1196), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1197), .A2(new_n693), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1190), .A3(new_n1187), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(KEYINPUT121), .A3(new_n1163), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1194), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1188), .A2(KEYINPUT120), .A3(new_n1189), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT120), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n1007), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n817), .B1(new_n1174), .B2(new_n807), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n822), .A2(new_n219), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n219), .B1(new_n269), .B2(G41), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n850), .A2(new_n1142), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n791), .A2(G128), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n792), .A2(G137), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n763), .A2(G150), .B1(G132), .B2(new_n765), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G125), .B2(new_n757), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT59), .ZN(new_n1215));
  AOI21_X1  g1015(.A(G33), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(G41), .B1(new_n795), .B2(G124), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(new_n843), .C2(new_n780), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1208), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n773), .A2(new_n221), .B1(new_n342), .B2(new_n762), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n780), .A2(new_n224), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n257), .B1(new_n766), .B2(new_n210), .C1(new_n213), .C2(new_n758), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n271), .B1(new_n785), .B2(new_n781), .ZN(new_n1224));
  NOR4_X1   g1024(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n436), .B2(new_n776), .C1(new_n308), .C2(new_n783), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT58), .Z(new_n1227));
  OAI21_X1  g1027(.A(new_n755), .B1(new_n1220), .B2(new_n1227), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT119), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1206), .A2(new_n1207), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1205), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1201), .A2(new_n1232), .ZN(G375));
  NOR2_X1   g1033(.A1(new_n824), .A2(G68), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n780), .A2(new_n224), .B1(new_n762), .B2(new_n219), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n271), .B(new_n1235), .C1(G128), .C2(new_n795), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n287), .B2(new_n783), .C1(new_n843), .C2(new_n773), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT122), .Z(new_n1238));
  OAI22_X1  g1038(.A1(new_n758), .A2(new_n846), .B1(new_n776), .B2(new_n842), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n765), .B2(new_n1142), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n308), .A2(new_n762), .B1(new_n478), .B2(new_n758), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n766), .A2(new_n213), .B1(new_n780), .B2(new_n221), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n783), .A2(new_n436), .B1(new_n785), .B2(new_n558), .ZN(new_n1244));
  NOR4_X1   g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n263), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1245), .B1(new_n210), .B2(new_n773), .C1(new_n781), .C2(new_n776), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1241), .A2(new_n1246), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT123), .Z(new_n1248));
  AOI211_X1 g1048(.A(new_n817), .B(new_n1234), .C1(new_n1248), .C2(new_n755), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n933), .A2(new_n807), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1128), .B2(new_n1006), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1252), .B(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1135), .A2(new_n984), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(G381));
  NAND3_X1  g1057(.A1(new_n1201), .A2(new_n1161), .A3(new_n1232), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1258), .A2(G384), .A3(G381), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1088), .A2(new_n1008), .A3(new_n1030), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(G393), .A2(G396), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1259), .A2(new_n1261), .A3(new_n1262), .ZN(G407));
  OAI211_X1 g1063(.A(G407), .B(G213), .C1(G343), .C2(new_n1258), .ZN(G409));
  INV_X1    g1064(.A(G213), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(G343), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1204), .A2(new_n984), .A3(new_n1195), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1196), .A2(new_n1007), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1161), .A2(new_n1268), .A3(new_n1230), .A4(new_n1269), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1193), .B(KEYINPUT57), .C1(new_n1204), .C2(new_n1195), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT121), .B1(new_n1199), .B2(new_n1163), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1231), .B1(new_n1273), .B2(new_n1198), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1267), .B(new_n1270), .C1(new_n1274), .C2(new_n1161), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1266), .A2(G2897), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1255), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1128), .A2(new_n1133), .A3(KEYINPUT60), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1278), .A2(new_n1135), .A3(new_n693), .A4(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1254), .A2(G384), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(G384), .B1(new_n1254), .B2(new_n1280), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1276), .B1(new_n1284), .B2(KEYINPUT126), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(KEYINPUT126), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT126), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1276), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1287), .B(new_n1288), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1285), .A2(new_n1286), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT61), .B1(new_n1275), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1197), .A2(new_n693), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1271), .A2(new_n1272), .A3(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(G378), .B1(new_n1293), .B2(new_n1231), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1294), .A2(new_n1267), .A3(new_n1270), .A4(new_n1284), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(KEYINPUT62), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1161), .B1(new_n1201), .B2(new_n1232), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1297), .A2(new_n1266), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT62), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1270), .A4(new_n1284), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1291), .A2(new_n1296), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(G387), .A2(G390), .ZN(new_n1302));
  INV_X1    g1102(.A(G396), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(G393), .B(new_n1303), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1302), .A2(new_n1260), .A3(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1304), .B1(new_n1302), .B2(new_n1260), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1301), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1270), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1284), .ZN(new_n1310));
  NOR4_X1   g1110(.A1(new_n1297), .A2(new_n1309), .A3(new_n1266), .A4(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(KEYINPUT63), .B1(new_n1311), .B2(KEYINPUT125), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1307), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT125), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1295), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1312), .A2(new_n1313), .A3(new_n1291), .A4(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1308), .A2(new_n1317), .ZN(G405));
  INV_X1    g1118(.A(new_n1258), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1310), .B1(new_n1319), .B2(new_n1297), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1294), .A2(new_n1258), .A3(new_n1284), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1307), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(KEYINPUT127), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1313), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT127), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1320), .A2(new_n1307), .A3(new_n1326), .A4(new_n1321), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1323), .A2(new_n1325), .A3(new_n1327), .ZN(G402));
endmodule


