

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745;

  NOR2_X1 U376 ( .A1(n614), .A2(n710), .ZN(n617) );
  INV_X1 U377 ( .A(G146), .ZN(n403) );
  XNOR2_X1 U378 ( .A(n403), .B(G125), .ZN(n488) );
  NOR2_X1 U379 ( .A1(n632), .A2(n710), .ZN(n634) );
  NOR2_X1 U380 ( .A1(n627), .A2(n710), .ZN(n628) );
  AND2_X4 U381 ( .A1(n611), .A2(n642), .ZN(n706) );
  NAND2_X2 U382 ( .A1(n564), .A2(n659), .ZN(n561) );
  XNOR2_X2 U383 ( .A(n407), .B(n460), .ZN(n564) );
  XNOR2_X2 U384 ( .A(n470), .B(KEYINPUT4), .ZN(n446) );
  XNOR2_X2 U385 ( .A(n414), .B(n413), .ZN(n470) );
  XNOR2_X2 U386 ( .A(n588), .B(KEYINPUT41), .ZN(n674) );
  NOR2_X1 U387 ( .A1(n623), .A2(n710), .ZN(n624) );
  NOR2_X1 U388 ( .A1(n556), .A2(n523), .ZN(n679) );
  NOR2_X1 U389 ( .A1(n745), .A2(n743), .ZN(n401) );
  INV_X1 U390 ( .A(n525), .ZN(n500) );
  XNOR2_X1 U391 ( .A(n380), .B(n379), .ZN(n722) );
  INV_X1 U392 ( .A(G143), .ZN(n413) );
  XNOR2_X1 U393 ( .A(n370), .B(n397), .ZN(n419) );
  NOR2_X1 U394 ( .A1(n679), .A2(n536), .ZN(n537) );
  XNOR2_X1 U395 ( .A(n393), .B(KEYINPUT32), .ZN(n741) );
  XNOR2_X1 U396 ( .A(n501), .B(KEYINPUT22), .ZN(n375) );
  NAND2_X1 U397 ( .A1(n500), .A2(n499), .ZN(n501) );
  NOR2_X1 U398 ( .A1(n516), .A2(n647), .ZN(n517) );
  OR2_X1 U399 ( .A1(n646), .A2(n559), .ZN(n516) );
  INV_X1 U400 ( .A(n527), .ZN(n653) );
  AND2_X1 U401 ( .A1(n661), .A2(n498), .ZN(n499) );
  XNOR2_X1 U402 ( .A(n448), .B(n447), .ZN(n527) );
  XNOR2_X1 U403 ( .A(n574), .B(KEYINPUT1), .ZN(n647) );
  XNOR2_X1 U404 ( .A(n429), .B(n430), .ZN(n441) );
  XNOR2_X1 U405 ( .A(n442), .B(n722), .ZN(n453) );
  XNOR2_X1 U406 ( .A(G119), .B(G116), .ZN(n430) );
  XNOR2_X1 U407 ( .A(G104), .B(G110), .ZN(n380) );
  INV_X2 U408 ( .A(G953), .ZN(n735) );
  XNOR2_X1 U409 ( .A(n517), .B(n355), .ZN(n673) );
  XOR2_X1 U410 ( .A(KEYINPUT102), .B(KEYINPUT33), .Z(n355) );
  NOR2_X2 U411 ( .A1(n374), .A2(n467), .ZN(n469) );
  XNOR2_X2 U412 ( .A(n561), .B(n462), .ZN(n374) );
  XNOR2_X1 U413 ( .A(n446), .B(n445), .ZN(n450) );
  XNOR2_X1 U414 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U415 ( .A(G134), .B(G131), .ZN(n444) );
  XNOR2_X1 U416 ( .A(n434), .B(KEYINPUT67), .ZN(n442) );
  XNOR2_X1 U417 ( .A(G101), .B(KEYINPUT68), .ZN(n434) );
  NOR2_X1 U418 ( .A1(G902), .A2(n703), .ZN(n456) );
  XOR2_X1 U419 ( .A(G137), .B(G140), .Z(n507) );
  XNOR2_X1 U420 ( .A(n450), .B(n449), .ZN(n728) );
  NAND2_X1 U421 ( .A1(n688), .A2(n741), .ZN(n544) );
  NOR2_X1 U422 ( .A1(n583), .A2(n691), .ZN(n371) );
  OR2_X1 U423 ( .A1(G902), .A2(G237), .ZN(n461) );
  XNOR2_X1 U424 ( .A(n358), .B(n438), .ZN(n384) );
  XOR2_X1 U425 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n438) );
  XNOR2_X1 U426 ( .A(G137), .B(G146), .ZN(n439) );
  XNOR2_X1 U427 ( .A(n488), .B(n402), .ZN(n506) );
  INV_X1 U428 ( .A(KEYINPUT10), .ZN(n402) );
  AND2_X1 U429 ( .A1(n419), .A2(n603), .ZN(n638) );
  NOR2_X1 U430 ( .A1(n653), .A2(n391), .ZN(n387) );
  NAND2_X1 U431 ( .A1(n653), .A2(n389), .ZN(n388) );
  NOR2_X1 U432 ( .A1(n390), .A2(n565), .ZN(n389) );
  AND2_X1 U433 ( .A1(n573), .A2(n653), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n513), .B(n512), .ZN(n644) );
  XNOR2_X1 U435 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U436 ( .A(G128), .B(G110), .ZN(n502) );
  NAND2_X1 U437 ( .A1(n735), .A2(G234), .ZN(n475) );
  XNOR2_X1 U438 ( .A(n506), .B(n507), .ZN(n727) );
  XNOR2_X1 U439 ( .A(n420), .B(KEYINPUT81), .ZN(n610) );
  XNOR2_X1 U440 ( .A(n585), .B(KEYINPUT39), .ZN(n592) );
  AND2_X1 U441 ( .A1(n584), .A2(n658), .ZN(n585) );
  INV_X1 U442 ( .A(KEYINPUT19), .ZN(n462) );
  XNOR2_X1 U443 ( .A(n421), .B(n728), .ZN(n703) );
  XNOR2_X1 U444 ( .A(n453), .B(n507), .ZN(n454) );
  NOR2_X1 U445 ( .A1(G952), .A2(n735), .ZN(n710) );
  NOR2_X1 U446 ( .A1(G953), .A2(G237), .ZN(n481) );
  INV_X1 U447 ( .A(n659), .ZN(n390) );
  XNOR2_X1 U448 ( .A(G122), .B(n411), .ZN(n410) );
  INV_X1 U449 ( .A(KEYINPUT16), .ZN(n411) );
  XNOR2_X1 U450 ( .A(G122), .B(G113), .ZN(n484) );
  XNOR2_X1 U451 ( .A(G140), .B(G143), .ZN(n489) );
  XOR2_X1 U452 ( .A(G104), .B(G131), .Z(n490) );
  NOR2_X1 U453 ( .A1(n541), .A2(n540), .ZN(n543) );
  INV_X1 U454 ( .A(KEYINPUT83), .ZN(n542) );
  XNOR2_X1 U455 ( .A(n432), .B(n362), .ZN(n378) );
  INV_X1 U456 ( .A(KEYINPUT48), .ZN(n397) );
  NAND2_X1 U457 ( .A1(G237), .A2(G234), .ZN(n463) );
  XNOR2_X1 U458 ( .A(n442), .B(n440), .ZN(n382) );
  NAND2_X1 U459 ( .A1(n396), .A2(n408), .ZN(n720) );
  NAND2_X1 U460 ( .A1(n441), .A2(n409), .ZN(n408) );
  NAND2_X1 U461 ( .A1(n412), .A2(n410), .ZN(n396) );
  XNOR2_X1 U462 ( .A(KEYINPUT16), .B(G122), .ZN(n409) );
  XOR2_X1 U463 ( .A(G122), .B(G116), .Z(n472) );
  XNOR2_X1 U464 ( .A(G134), .B(G107), .ZN(n471) );
  AND2_X1 U465 ( .A1(G227), .A2(n735), .ZN(n451) );
  XNOR2_X1 U466 ( .A(n377), .B(n376), .ZN(n457) );
  XNOR2_X1 U467 ( .A(n453), .B(n446), .ZN(n376) );
  XNOR2_X1 U468 ( .A(n720), .B(n369), .ZN(n377) );
  XNOR2_X1 U469 ( .A(n378), .B(n433), .ZN(n369) );
  BUF_X1 U470 ( .A(n564), .Z(n593) );
  XNOR2_X1 U471 ( .A(n570), .B(n569), .ZN(n584) );
  NAND2_X1 U472 ( .A1(n568), .A2(n385), .ZN(n570) );
  NOR2_X1 U473 ( .A1(n576), .A2(n575), .ZN(n589) );
  INV_X1 U474 ( .A(KEYINPUT28), .ZN(n372) );
  INV_X1 U475 ( .A(n653), .ZN(n415) );
  XOR2_X1 U476 ( .A(n527), .B(KEYINPUT6), .Z(n559) );
  INV_X1 U477 ( .A(G107), .ZN(n379) );
  XNOR2_X1 U478 ( .A(n404), .B(n727), .ZN(n626) );
  XNOR2_X1 U479 ( .A(n406), .B(n405), .ZN(n404) );
  XNOR2_X1 U480 ( .A(n505), .B(n360), .ZN(n405) );
  XNOR2_X1 U481 ( .A(n521), .B(n520), .ZN(n739) );
  NOR2_X1 U482 ( .A1(n519), .A2(n572), .ZN(n520) );
  XNOR2_X1 U483 ( .A(n395), .B(n394), .ZN(n704) );
  XNOR2_X1 U484 ( .A(n703), .B(n702), .ZN(n394) );
  AND2_X1 U485 ( .A1(n556), .A2(n415), .ZN(n356) );
  AND2_X1 U486 ( .A1(n565), .A2(n390), .ZN(n357) );
  AND2_X1 U487 ( .A1(G210), .A2(n481), .ZN(n358) );
  NOR2_X1 U488 ( .A1(n577), .A2(n374), .ZN(n359) );
  XNOR2_X1 U489 ( .A(KEYINPUT23), .B(G119), .ZN(n360) );
  AND2_X1 U490 ( .A1(n676), .A2(n424), .ZN(n361) );
  AND2_X1 U491 ( .A1(G224), .A2(n735), .ZN(n362) );
  XOR2_X1 U492 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n363) );
  OR2_X1 U493 ( .A1(n646), .A2(n527), .ZN(n364) );
  AND2_X1 U494 ( .A1(n603), .A2(KEYINPUT2), .ZN(n365) );
  NOR2_X1 U495 ( .A1(n647), .A2(n364), .ZN(n366) );
  OR2_X1 U496 ( .A1(n392), .A2(n357), .ZN(n367) );
  NAND2_X1 U497 ( .A1(n368), .A2(n398), .ZN(n370) );
  XNOR2_X1 U498 ( .A(n401), .B(n422), .ZN(n368) );
  NOR2_X1 U499 ( .A1(n387), .A2(n367), .ZN(n386) );
  AND2_X1 U500 ( .A1(n388), .A2(n386), .ZN(n385) );
  NAND2_X1 U501 ( .A1(n544), .A2(KEYINPUT44), .ZN(n515) );
  INV_X1 U502 ( .A(n488), .ZN(n432) );
  NOR2_X2 U503 ( .A1(n375), .A2(n597), .ZN(n522) );
  NAND2_X1 U504 ( .A1(n359), .A2(n663), .ZN(n578) );
  XNOR2_X1 U505 ( .A(n371), .B(n400), .ZN(n399) );
  XNOR2_X1 U506 ( .A(n373), .B(n372), .ZN(n576) );
  NAND2_X1 U507 ( .A1(n504), .A2(G221), .ZN(n406) );
  OR2_X1 U508 ( .A1(n375), .A2(n418), .ZN(n393) );
  XNOR2_X2 U509 ( .A(n456), .B(n455), .ZN(n574) );
  XNOR2_X1 U510 ( .A(n450), .B(n381), .ZN(n629) );
  XNOR2_X1 U511 ( .A(n383), .B(n382), .ZN(n381) );
  XNOR2_X1 U512 ( .A(n441), .B(n384), .ZN(n383) );
  INV_X1 U513 ( .A(n565), .ZN(n391) );
  INV_X1 U514 ( .A(n566), .ZN(n392) );
  NAND2_X1 U515 ( .A1(n706), .A2(G469), .ZN(n395) );
  NAND2_X1 U516 ( .A1(n457), .A2(n604), .ZN(n407) );
  XNOR2_X1 U517 ( .A(n454), .B(n452), .ZN(n421) );
  AND2_X1 U518 ( .A1(n399), .A2(n699), .ZN(n398) );
  INV_X1 U519 ( .A(KEYINPUT71), .ZN(n400) );
  INV_X1 U520 ( .A(n441), .ZN(n412) );
  XNOR2_X2 U521 ( .A(G128), .B(KEYINPUT64), .ZN(n414) );
  NAND2_X1 U522 ( .A1(n416), .A2(n356), .ZN(n688) );
  XNOR2_X1 U523 ( .A(n522), .B(n417), .ZN(n416) );
  INV_X1 U524 ( .A(KEYINPUT101), .ZN(n417) );
  NAND2_X1 U525 ( .A1(n514), .A2(n556), .ZN(n418) );
  NAND2_X1 U526 ( .A1(n419), .A2(n365), .ZN(n420) );
  XNOR2_X2 U527 ( .A(n469), .B(n468), .ZN(n525) );
  XNOR2_X1 U528 ( .A(KEYINPUT46), .B(KEYINPUT82), .ZN(n422) );
  AND2_X1 U529 ( .A1(n674), .A2(n673), .ZN(n423) );
  NOR2_X1 U530 ( .A1(n675), .A2(n423), .ZN(n424) );
  INV_X1 U531 ( .A(n558), .ZN(n498) );
  INV_X1 U532 ( .A(n701), .ZN(n602) );
  INV_X1 U533 ( .A(KEYINPUT69), .ZN(n443) );
  NOR2_X1 U534 ( .A1(n700), .A2(n602), .ZN(n603) );
  XNOR2_X1 U535 ( .A(n459), .B(n458), .ZN(n460) );
  BUF_X1 U536 ( .A(n638), .Z(n732) );
  XNOR2_X1 U537 ( .A(n451), .B(G146), .ZN(n452) );
  INV_X1 U538 ( .A(KEYINPUT63), .ZN(n633) );
  XNOR2_X1 U539 ( .A(n678), .B(n677), .ZN(G75) );
  INV_X1 U540 ( .A(G113), .ZN(n425) );
  NAND2_X1 U541 ( .A1(KEYINPUT3), .A2(n425), .ZN(n428) );
  INV_X1 U542 ( .A(KEYINPUT3), .ZN(n426) );
  NAND2_X1 U543 ( .A1(n426), .A2(G113), .ZN(n427) );
  NAND2_X1 U544 ( .A1(n428), .A2(n427), .ZN(n429) );
  XNOR2_X1 U545 ( .A(KEYINPUT74), .B(KEYINPUT18), .ZN(n431) );
  XNOR2_X1 U546 ( .A(n363), .B(n431), .ZN(n433) );
  XOR2_X1 U547 ( .A(KEYINPUT54), .B(KEYINPUT114), .Z(n436) );
  XNOR2_X1 U548 ( .A(KEYINPUT84), .B(KEYINPUT55), .ZN(n435) );
  XNOR2_X1 U549 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U550 ( .A(n457), .B(n437), .Z(n613) );
  XNOR2_X1 U551 ( .A(n439), .B(KEYINPUT92), .ZN(n440) );
  NOR2_X1 U552 ( .A1(G902), .A2(n629), .ZN(n448) );
  XNOR2_X1 U553 ( .A(KEYINPUT94), .B(G472), .ZN(n447) );
  INV_X1 U554 ( .A(KEYINPUT89), .ZN(n449) );
  XNOR2_X1 U555 ( .A(KEYINPUT70), .B(G469), .ZN(n455) );
  INV_X1 U556 ( .A(n647), .ZN(n597) );
  XNOR2_X1 U557 ( .A(G902), .B(KEYINPUT15), .ZN(n604) );
  NAND2_X1 U558 ( .A1(n461), .A2(G210), .ZN(n459) );
  XNOR2_X1 U559 ( .A(KEYINPUT75), .B(KEYINPUT86), .ZN(n458) );
  NAND2_X1 U560 ( .A1(G214), .A2(n461), .ZN(n659) );
  XNOR2_X1 U561 ( .A(n463), .B(KEYINPUT14), .ZN(n465) );
  NAND2_X1 U562 ( .A1(G952), .A2(n465), .ZN(n672) );
  NOR2_X1 U563 ( .A1(G953), .A2(n672), .ZN(n464) );
  XOR2_X1 U564 ( .A(KEYINPUT87), .B(n464), .Z(n552) );
  XOR2_X1 U565 ( .A(KEYINPUT88), .B(G898), .Z(n714) );
  NAND2_X1 U566 ( .A1(G953), .A2(n714), .ZN(n723) );
  NAND2_X1 U567 ( .A1(G902), .A2(n465), .ZN(n550) );
  NOR2_X1 U568 ( .A1(n723), .A2(n550), .ZN(n466) );
  NOR2_X1 U569 ( .A1(n552), .A2(n466), .ZN(n467) );
  INV_X1 U570 ( .A(KEYINPUT0), .ZN(n468) );
  INV_X1 U571 ( .A(n470), .ZN(n474) );
  XNOR2_X1 U572 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U573 ( .A(n474), .B(n473), .ZN(n479) );
  XOR2_X1 U574 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n477) );
  XOR2_X1 U575 ( .A(KEYINPUT8), .B(n475), .Z(n504) );
  NAND2_X1 U576 ( .A1(G217), .A2(n504), .ZN(n476) );
  XNOR2_X1 U577 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U578 ( .A(n479), .B(n478), .ZN(n705) );
  NOR2_X1 U579 ( .A1(G902), .A2(n705), .ZN(n480) );
  XOR2_X1 U580 ( .A(G478), .B(n480), .Z(n531) );
  XNOR2_X1 U581 ( .A(KEYINPUT13), .B(G475), .ZN(n495) );
  XOR2_X1 U582 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n483) );
  NAND2_X1 U583 ( .A1(n481), .A2(G214), .ZN(n482) );
  XNOR2_X1 U584 ( .A(n483), .B(n482), .ZN(n487) );
  XOR2_X1 U585 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n485) );
  XNOR2_X1 U586 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U587 ( .A(n487), .B(n486), .Z(n493) );
  XNOR2_X1 U588 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U589 ( .A(n506), .B(n491), .ZN(n492) );
  XNOR2_X1 U590 ( .A(n493), .B(n492), .ZN(n618) );
  NOR2_X1 U591 ( .A1(G902), .A2(n618), .ZN(n494) );
  XNOR2_X1 U592 ( .A(n495), .B(n494), .ZN(n532) );
  NOR2_X1 U593 ( .A1(n531), .A2(n532), .ZN(n661) );
  NAND2_X1 U594 ( .A1(G234), .A2(n604), .ZN(n496) );
  XNOR2_X1 U595 ( .A(KEYINPUT20), .B(n496), .ZN(n508) );
  NAND2_X1 U596 ( .A1(n508), .A2(G221), .ZN(n497) );
  XNOR2_X1 U597 ( .A(n497), .B(KEYINPUT21), .ZN(n558) );
  XOR2_X1 U598 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n503) );
  XNOR2_X1 U599 ( .A(n503), .B(n502), .ZN(n505) );
  NOR2_X1 U600 ( .A1(n626), .A2(G902), .ZN(n513) );
  NAND2_X1 U601 ( .A1(n508), .A2(G217), .ZN(n511) );
  XNOR2_X1 U602 ( .A(KEYINPUT91), .B(KEYINPUT25), .ZN(n509) );
  XNOR2_X1 U603 ( .A(n509), .B(KEYINPUT73), .ZN(n510) );
  INV_X1 U604 ( .A(n644), .ZN(n556) );
  AND2_X1 U605 ( .A1(n559), .A2(n597), .ZN(n514) );
  XNOR2_X1 U606 ( .A(KEYINPUT65), .B(n515), .ZN(n541) );
  INV_X1 U607 ( .A(KEYINPUT35), .ZN(n521) );
  NAND2_X1 U608 ( .A1(n531), .A2(n532), .ZN(n572) );
  NAND2_X1 U609 ( .A1(n498), .A2(n644), .ZN(n646) );
  INV_X1 U610 ( .A(n525), .ZN(n528) );
  NAND2_X1 U611 ( .A1(n673), .A2(n528), .ZN(n518) );
  XNOR2_X1 U612 ( .A(n518), .B(KEYINPUT34), .ZN(n519) );
  NAND2_X1 U613 ( .A1(KEYINPUT44), .A2(n739), .ZN(n539) );
  NAND2_X1 U614 ( .A1(n559), .A2(n522), .ZN(n523) );
  NOR2_X2 U615 ( .A1(n574), .A2(n646), .ZN(n567) );
  NAND2_X1 U616 ( .A1(n415), .A2(n567), .ZN(n524) );
  NOR2_X1 U617 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U618 ( .A(KEYINPUT95), .B(n526), .Z(n684) );
  NAND2_X1 U619 ( .A1(n366), .A2(n528), .ZN(n530) );
  XNOR2_X1 U620 ( .A(KEYINPUT31), .B(KEYINPUT96), .ZN(n529) );
  XNOR2_X1 U621 ( .A(n530), .B(n529), .ZN(n696) );
  NOR2_X1 U622 ( .A1(n684), .A2(n696), .ZN(n535) );
  INV_X1 U623 ( .A(n531), .ZN(n533) );
  NAND2_X1 U624 ( .A1(n532), .A2(n533), .ZN(n681) );
  NOR2_X1 U625 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U626 ( .A(n534), .B(KEYINPUT99), .ZN(n683) );
  NAND2_X1 U627 ( .A1(n681), .A2(n683), .ZN(n663) );
  XOR2_X1 U628 ( .A(KEYINPUT78), .B(n663), .Z(n579) );
  NOR2_X1 U629 ( .A1(n535), .A2(n579), .ZN(n536) );
  XNOR2_X1 U630 ( .A(n537), .B(KEYINPUT100), .ZN(n538) );
  NAND2_X1 U631 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U632 ( .A(n543), .B(n542), .ZN(n548) );
  INV_X1 U633 ( .A(n544), .ZN(n546) );
  NOR2_X1 U634 ( .A1(n739), .A2(KEYINPUT44), .ZN(n545) );
  NAND2_X1 U635 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U636 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X2 U637 ( .A(n549), .B(KEYINPUT45), .ZN(n716) );
  NOR2_X1 U638 ( .A1(G900), .A2(n550), .ZN(n551) );
  NAND2_X1 U639 ( .A1(n551), .A2(G953), .ZN(n554) );
  INV_X1 U640 ( .A(n552), .ZN(n553) );
  NAND2_X1 U641 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U642 ( .A(n555), .B(KEYINPUT76), .ZN(n566) );
  NAND2_X1 U643 ( .A1(n556), .A2(n566), .ZN(n557) );
  NOR2_X1 U644 ( .A1(n558), .A2(n557), .ZN(n573) );
  NOR2_X1 U645 ( .A1(n559), .A2(n681), .ZN(n560) );
  NAND2_X1 U646 ( .A1(n573), .A2(n560), .ZN(n594) );
  NOR2_X1 U647 ( .A1(n561), .A2(n594), .ZN(n562) );
  XNOR2_X1 U648 ( .A(KEYINPUT36), .B(n562), .ZN(n563) );
  NAND2_X1 U649 ( .A1(n563), .A2(n597), .ZN(n699) );
  XOR2_X1 U650 ( .A(KEYINPUT30), .B(KEYINPUT105), .Z(n565) );
  XNOR2_X1 U651 ( .A(n567), .B(KEYINPUT104), .ZN(n568) );
  INV_X1 U652 ( .A(KEYINPUT72), .ZN(n569) );
  NAND2_X1 U653 ( .A1(n593), .A2(n584), .ZN(n571) );
  NOR2_X1 U654 ( .A1(n572), .A2(n571), .ZN(n691) );
  XNOR2_X1 U655 ( .A(n574), .B(KEYINPUT106), .ZN(n575) );
  INV_X1 U656 ( .A(n589), .ZN(n577) );
  NAND2_X1 U657 ( .A1(n578), .A2(KEYINPUT47), .ZN(n582) );
  NOR2_X1 U658 ( .A1(KEYINPUT47), .A2(n579), .ZN(n580) );
  NAND2_X1 U659 ( .A1(n580), .A2(n359), .ZN(n581) );
  NAND2_X1 U660 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U661 ( .A(KEYINPUT38), .B(n593), .Z(n658) );
  NOR2_X1 U662 ( .A1(n681), .A2(n592), .ZN(n586) );
  XNOR2_X1 U663 ( .A(n586), .B(KEYINPUT40), .ZN(n745) );
  XOR2_X1 U664 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n591) );
  NAND2_X1 U665 ( .A1(n659), .A2(n658), .ZN(n587) );
  XNOR2_X1 U666 ( .A(KEYINPUT107), .B(n587), .ZN(n664) );
  NAND2_X1 U667 ( .A1(n664), .A2(n661), .ZN(n588) );
  NAND2_X1 U668 ( .A1(n589), .A2(n674), .ZN(n590) );
  XNOR2_X1 U669 ( .A(n591), .B(n590), .ZN(n743) );
  NOR2_X1 U670 ( .A1(n683), .A2(n592), .ZN(n700) );
  INV_X1 U671 ( .A(n593), .ZN(n601) );
  XNOR2_X1 U672 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n599) );
  INV_X1 U673 ( .A(n594), .ZN(n595) );
  NAND2_X1 U674 ( .A1(n595), .A2(n659), .ZN(n596) );
  NOR2_X1 U675 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U676 ( .A(n599), .B(n598), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n601), .A2(n600), .ZN(n701) );
  INV_X1 U678 ( .A(n604), .ZN(n606) );
  AND2_X1 U679 ( .A1(n638), .A2(n606), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n716), .A2(n605), .ZN(n609) );
  XNOR2_X1 U681 ( .A(n606), .B(KEYINPUT80), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n607), .A2(KEYINPUT2), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n610), .A2(n716), .ZN(n642) );
  NAND2_X1 U685 ( .A1(n706), .A2(G210), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n613), .B(n612), .ZN(n614) );
  INV_X1 U687 ( .A(KEYINPUT115), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n615), .B(KEYINPUT56), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n617), .B(n616), .ZN(G51) );
  XOR2_X1 U690 ( .A(KEYINPUT59), .B(KEYINPUT116), .Z(n620) );
  XNOR2_X1 U691 ( .A(n618), .B(KEYINPUT66), .ZN(n619) );
  XNOR2_X1 U692 ( .A(n620), .B(n619), .ZN(n622) );
  NAND2_X1 U693 ( .A1(n706), .A2(G475), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U695 ( .A(n624), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U696 ( .A1(G217), .A2(n706), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n628), .B(KEYINPUT118), .ZN(G66) );
  XNOR2_X1 U699 ( .A(n629), .B(KEYINPUT62), .ZN(n631) );
  NAND2_X1 U700 ( .A1(G472), .A2(n706), .ZN(n630) );
  XNOR2_X1 U701 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U702 ( .A(n634), .B(n633), .ZN(G57) );
  INV_X1 U703 ( .A(n716), .ZN(n636) );
  XOR2_X1 U704 ( .A(KEYINPUT2), .B(KEYINPUT77), .Z(n639) );
  INV_X1 U705 ( .A(n639), .ZN(n635) );
  NAND2_X1 U706 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U707 ( .A(n637), .B(KEYINPUT79), .ZN(n641) );
  NOR2_X1 U708 ( .A1(n732), .A2(n639), .ZN(n640) );
  NOR2_X1 U709 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U710 ( .A1(n643), .A2(n642), .ZN(n676) );
  NOR2_X1 U711 ( .A1(n498), .A2(n644), .ZN(n645) );
  XNOR2_X1 U712 ( .A(KEYINPUT49), .B(n645), .ZN(n651) );
  NAND2_X1 U713 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U714 ( .A(n648), .B(KEYINPUT50), .ZN(n649) );
  XNOR2_X1 U715 ( .A(KEYINPUT110), .B(n649), .ZN(n650) );
  NAND2_X1 U716 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U717 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U718 ( .A(KEYINPUT111), .B(n654), .Z(n655) );
  NOR2_X1 U719 ( .A1(n366), .A2(n655), .ZN(n656) );
  XNOR2_X1 U720 ( .A(KEYINPUT51), .B(n656), .ZN(n657) );
  NAND2_X1 U721 ( .A1(n657), .A2(n674), .ZN(n669) );
  OR2_X1 U722 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U723 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U724 ( .A(n662), .B(KEYINPUT112), .ZN(n666) );
  NAND2_X1 U725 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U726 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U727 ( .A1(n667), .A2(n673), .ZN(n668) );
  NAND2_X1 U728 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U729 ( .A(KEYINPUT52), .B(n670), .Z(n671) );
  NOR2_X1 U730 ( .A1(n672), .A2(n671), .ZN(n675) );
  NAND2_X1 U731 ( .A1(n735), .A2(n361), .ZN(n678) );
  XNOR2_X1 U732 ( .A(KEYINPUT113), .B(KEYINPUT53), .ZN(n677) );
  XNOR2_X1 U733 ( .A(G101), .B(n679), .ZN(n680) );
  XNOR2_X1 U734 ( .A(n680), .B(KEYINPUT109), .ZN(G3) );
  INV_X1 U735 ( .A(n681), .ZN(n693) );
  NAND2_X1 U736 ( .A1(n693), .A2(n684), .ZN(n682) );
  XNOR2_X1 U737 ( .A(G104), .B(n682), .ZN(G6) );
  XOR2_X1 U738 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n686) );
  INV_X1 U739 ( .A(n683), .ZN(n695) );
  NAND2_X1 U740 ( .A1(n684), .A2(n695), .ZN(n685) );
  XNOR2_X1 U741 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U742 ( .A(G107), .B(n687), .ZN(G9) );
  XNOR2_X1 U743 ( .A(G110), .B(n688), .ZN(G12) );
  XOR2_X1 U744 ( .A(G128), .B(KEYINPUT29), .Z(n690) );
  NAND2_X1 U745 ( .A1(n359), .A2(n695), .ZN(n689) );
  XNOR2_X1 U746 ( .A(n690), .B(n689), .ZN(G30) );
  XOR2_X1 U747 ( .A(G143), .B(n691), .Z(G45) );
  NAND2_X1 U748 ( .A1(n359), .A2(n693), .ZN(n692) );
  XNOR2_X1 U749 ( .A(n692), .B(G146), .ZN(G48) );
  NAND2_X1 U750 ( .A1(n696), .A2(n693), .ZN(n694) );
  XNOR2_X1 U751 ( .A(n694), .B(G113), .ZN(G15) );
  NAND2_X1 U752 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U753 ( .A(n697), .B(G116), .ZN(G18) );
  XOR2_X1 U754 ( .A(G125), .B(KEYINPUT37), .Z(n698) );
  XNOR2_X1 U755 ( .A(n699), .B(n698), .ZN(G27) );
  XOR2_X1 U756 ( .A(G134), .B(n700), .Z(G36) );
  XNOR2_X1 U757 ( .A(G140), .B(n701), .ZN(G42) );
  XOR2_X1 U758 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n702) );
  NOR2_X1 U759 ( .A1(n710), .A2(n704), .ZN(G54) );
  XOR2_X1 U760 ( .A(n705), .B(KEYINPUT117), .Z(n708) );
  NAND2_X1 U761 ( .A1(n706), .A2(G478), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U763 ( .A1(n710), .A2(n709), .ZN(G63) );
  NAND2_X1 U764 ( .A1(G224), .A2(G953), .ZN(n711) );
  XNOR2_X1 U765 ( .A(n711), .B(KEYINPUT61), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n712), .B(KEYINPUT119), .ZN(n713) );
  NOR2_X1 U767 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n715), .B(KEYINPUT120), .ZN(n718) );
  AND2_X1 U769 ( .A1(n716), .A2(n735), .ZN(n717) );
  NOR2_X1 U770 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U771 ( .A(n719), .B(KEYINPUT121), .Z(n726) );
  XOR2_X1 U772 ( .A(n720), .B(G101), .Z(n721) );
  XNOR2_X1 U773 ( .A(n722), .B(n721), .ZN(n724) );
  NAND2_X1 U774 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U775 ( .A(n726), .B(n725), .ZN(G69) );
  XNOR2_X1 U776 ( .A(n728), .B(n727), .ZN(n733) );
  XOR2_X1 U777 ( .A(G227), .B(n733), .Z(n729) );
  NAND2_X1 U778 ( .A1(n729), .A2(G900), .ZN(n730) );
  NAND2_X1 U779 ( .A1(G953), .A2(n730), .ZN(n731) );
  XOR2_X1 U780 ( .A(KEYINPUT123), .B(n731), .Z(n738) );
  XNOR2_X1 U781 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U782 ( .A(n734), .B(KEYINPUT122), .ZN(n736) );
  NAND2_X1 U783 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U784 ( .A1(n738), .A2(n737), .ZN(G72) );
  XOR2_X1 U785 ( .A(G122), .B(n739), .Z(n740) );
  XNOR2_X1 U786 ( .A(KEYINPUT124), .B(n740), .ZN(G24) );
  XOR2_X1 U787 ( .A(G119), .B(n741), .Z(n742) );
  XNOR2_X1 U788 ( .A(KEYINPUT125), .B(n742), .ZN(G21) );
  XOR2_X1 U789 ( .A(G137), .B(n743), .Z(n744) );
  XNOR2_X1 U790 ( .A(KEYINPUT126), .B(n744), .ZN(G39) );
  XOR2_X1 U791 ( .A(G131), .B(n745), .Z(G33) );
endmodule

