//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT0), .B(G128), .Z(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n193), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G134), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n205), .B1(new_n204), .B2(new_n206), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n206), .A2(new_n199), .A3(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n200), .A2(new_n202), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G137), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n198), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n204), .A2(new_n206), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n215), .A2(new_n198), .A3(new_n212), .A4(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n197), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n192), .A2(KEYINPUT1), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n222), .A2(G128), .B1(new_n189), .B2(new_n191), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n204), .B1(G134), .B2(new_n203), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n217), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  OR2_X1    g042(.A1(KEYINPUT68), .A2(KEYINPUT30), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT68), .A2(KEYINPUT30), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n219), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n197), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n215), .A2(new_n212), .A3(new_n216), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G131), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n232), .B1(new_n234), .B2(new_n217), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n217), .A2(new_n225), .A3(new_n227), .ZN(new_n236));
  OAI211_X1 g050(.A(KEYINPUT68), .B(KEYINPUT30), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT66), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G116), .ZN(new_n244));
  INV_X1    g058(.A(G116), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n245), .A2(KEYINPUT67), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(KEYINPUT67), .ZN(new_n247));
  OAI21_X1  g061(.A(G119), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT2), .B(G113), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n250), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n244), .A2(new_n248), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n219), .A2(new_n255), .A3(new_n228), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n219), .A2(KEYINPUT69), .A3(new_n255), .A4(new_n228), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n238), .A2(new_n254), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT31), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT70), .B(G953), .ZN(new_n262));
  INV_X1    g076(.A(G237), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(G210), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT72), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G101), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n260), .A2(new_n261), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n256), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n219), .A2(new_n228), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n254), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n235), .A2(new_n236), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT69), .B1(new_n277), .B2(new_n255), .ZN(new_n278));
  NOR4_X1   g092(.A1(new_n235), .A2(new_n236), .A3(new_n257), .A4(new_n254), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n276), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n274), .B1(new_n280), .B2(KEYINPUT28), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n271), .B1(new_n281), .B2(new_n270), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n283));
  AOI211_X1 g097(.A(new_n283), .B(new_n261), .C1(new_n260), .C2(new_n270), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n238), .A2(new_n254), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n258), .A2(new_n259), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(new_n270), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT73), .B1(new_n287), .B2(KEYINPUT31), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n282), .A2(new_n284), .A3(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(G472), .A2(G902), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n187), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n278), .A2(new_n279), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n255), .B1(new_n231), .B2(new_n237), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n293), .A2(new_n269), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n283), .B1(new_n295), .B2(new_n261), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n258), .A2(new_n259), .B1(new_n254), .B2(new_n275), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n273), .B1(new_n297), .B2(new_n272), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n269), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n287), .A2(KEYINPUT73), .A3(KEYINPUT31), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n296), .A2(new_n299), .A3(new_n271), .A4(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT32), .A3(new_n290), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n297), .B2(new_n272), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n280), .A2(KEYINPUT74), .A3(KEYINPUT28), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n273), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n270), .A2(KEYINPUT29), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n303), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n298), .A2(new_n270), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n260), .A2(new_n269), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT29), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G472), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n292), .A2(new_n302), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G221), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT9), .B(G234), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT80), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n315), .B1(new_n317), .B2(new_n303), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G110), .B(G140), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT81), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n262), .A2(G227), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G107), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(G104), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n327));
  INV_X1    g141(.A(G104), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(G107), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n326), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT84), .B(G101), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT3), .B1(new_n328), .B2(G107), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT83), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n325), .A2(G104), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(KEYINPUT83), .A3(KEYINPUT3), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n330), .A2(new_n331), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n329), .A2(new_n327), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n328), .A2(G107), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n334), .A2(new_n336), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n337), .A2(KEYINPUT4), .B1(new_n340), .B2(G101), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n340), .A2(KEYINPUT4), .A3(G101), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n197), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT85), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT85), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n345), .B(new_n197), .C1(new_n341), .C2(new_n342), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n234), .A2(new_n217), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G101), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(new_n335), .B2(new_n339), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(KEYINPUT86), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT86), .ZN(new_n353));
  AOI211_X1 g167(.A(new_n353), .B(new_n350), .C1(new_n335), .C2(new_n339), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT87), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n220), .B1(new_n222), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n189), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n193), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n355), .B(new_n337), .C1(new_n221), .C2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n355), .A2(new_n337), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n363), .A2(new_n361), .A3(new_n224), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n347), .A2(new_n349), .A3(new_n362), .A4(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n364), .B1(new_n344), .B2(new_n346), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n349), .B1(new_n368), .B2(new_n362), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n324), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n337), .ZN(new_n371));
  OAI21_X1  g185(.A(G101), .B1(new_n329), .B2(new_n326), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n353), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n351), .A2(KEYINPUT86), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n224), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n360), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n348), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT89), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n377), .A2(new_n348), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT12), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n377), .A2(new_n348), .A3(new_n384), .A4(new_n378), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n380), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n366), .A3(new_n323), .ZN(new_n387));
  AOI211_X1 g201(.A(G469), .B(G902), .C1(new_n370), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n366), .ZN(new_n389));
  XOR2_X1   g203(.A(new_n323), .B(KEYINPUT82), .Z(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n347), .A2(new_n362), .A3(new_n365), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n348), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n366), .A3(new_n323), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(G469), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G469), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(new_n303), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n319), .B1(new_n388), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G214), .B1(G237), .B2(G902), .ZN(new_n401));
  INV_X1    g215(.A(G125), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n225), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n197), .A2(G125), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G953), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G224), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n405), .B(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n254), .B1(new_n341), .B2(new_n342), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT90), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n244), .A2(new_n248), .A3(KEYINPUT5), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT5), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n243), .A2(new_n413), .A3(G116), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n414), .A3(G113), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n415), .A2(new_n253), .A3(new_n337), .A4(new_n355), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT90), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n254), .B(new_n417), .C1(new_n341), .C2(new_n342), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n411), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(G110), .B(G122), .Z(new_n420));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(KEYINPUT91), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n422), .B1(new_n419), .B2(new_n420), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n411), .A2(new_n418), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT92), .ZN(new_n428));
  INV_X1    g242(.A(new_n420), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .A4(new_n416), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n411), .A2(new_n429), .A3(new_n416), .A4(new_n418), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT92), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(KEYINPUT6), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n409), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n415), .A2(new_n253), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n363), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(KEYINPUT94), .A3(new_n416), .ZN(new_n437));
  OR3_X1    g251(.A1(new_n435), .A2(KEYINPUT94), .A3(new_n363), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT93), .B(KEYINPUT8), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n420), .B(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT95), .B(KEYINPUT7), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n403), .B(new_n404), .C1(new_n408), .C2(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n405), .A2(KEYINPUT7), .A3(new_n407), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT96), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n445), .B(new_n446), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n431), .A2(KEYINPUT92), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n431), .A2(KEYINPUT92), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n444), .B(new_n447), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n303), .ZN(new_n451));
  OAI21_X1  g265(.A(G210), .B1(G237), .B2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n434), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n409), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n448), .A2(new_n449), .A3(new_n421), .ZN(new_n456));
  INV_X1    g270(.A(new_n425), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n423), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n455), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n441), .A2(new_n443), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n460), .B1(new_n430), .B2(new_n432), .ZN(new_n461));
  AOI21_X1  g275(.A(G902), .B1(new_n461), .B2(new_n447), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n452), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n401), .B1(new_n454), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n400), .B1(new_n464), .B2(KEYINPUT97), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT22), .B(G137), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n243), .A2(KEYINPUT23), .A3(G128), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n239), .A2(G128), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(new_n243), .B2(G128), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(KEYINPUT23), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G110), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT24), .B(G110), .Z(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT75), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n471), .ZN(new_n476));
  XNOR2_X1  g290(.A(G125), .B(G140), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT16), .ZN(new_n478));
  INV_X1    g292(.A(G140), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G125), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n480), .A2(KEYINPUT16), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(G146), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(G146), .B1(new_n478), .B2(new_n481), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n473), .B(new_n476), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT76), .ZN(new_n486));
  OAI22_X1  g300(.A1(new_n472), .A2(G110), .B1(new_n475), .B2(new_n471), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n402), .A2(G140), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT77), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT77), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n477), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n492), .A3(new_n188), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n487), .A2(new_n482), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n468), .B1(new_n486), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OR2_X1    g310(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n486), .A2(new_n494), .A3(new_n468), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n496), .A2(new_n303), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n500));
  INV_X1    g314(.A(new_n498), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(new_n495), .ZN(new_n502));
  NAND2_X1  g316(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n502), .A2(new_n303), .A3(new_n503), .A4(new_n497), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n303), .A2(G234), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n500), .A2(new_n504), .A3(G217), .A4(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT79), .ZN(new_n507));
  AOI21_X1  g321(.A(G902), .B1(new_n505), .B2(G217), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n502), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n507), .B1(new_n502), .B2(new_n508), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(KEYINPUT70), .A2(G953), .ZN(new_n514));
  NOR2_X1   g328(.A1(KEYINPUT70), .A2(G953), .ZN(new_n515));
  OAI211_X1 g329(.A(G214), .B(new_n263), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n190), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n262), .A2(G143), .A3(G214), .A4(new_n263), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G131), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n518), .A3(new_n198), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n483), .A2(new_n484), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(KEYINPUT17), .A3(G131), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n493), .B1(new_n188), .B2(new_n477), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT98), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT18), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(new_n198), .ZN(new_n530));
  OAI221_X1 g344(.A(new_n527), .B1(new_n519), .B2(new_n530), .C1(new_n520), .C2(new_n529), .ZN(new_n531));
  XNOR2_X1  g345(.A(G113), .B(G122), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT100), .B(G104), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n526), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT101), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT101), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n526), .A2(new_n531), .A3(new_n537), .A4(new_n534), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n534), .B1(new_n526), .B2(new_n531), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n540), .A2(KEYINPUT104), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(KEYINPUT104), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n303), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT105), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n543), .A2(KEYINPUT105), .A3(new_n303), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(G475), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n520), .A2(new_n522), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT19), .B1(new_n490), .B2(KEYINPUT99), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n491), .B1(KEYINPUT99), .B2(KEYINPUT19), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n489), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n188), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(new_n482), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n534), .B1(new_n531), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n539), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(G475), .A2(G902), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT20), .B1(new_n558), .B2(KEYINPUT102), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(KEYINPUT102), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n557), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT103), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n560), .B1(new_n539), .B2(new_n556), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT103), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n559), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n557), .A2(new_n558), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT20), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n563), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G952), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(G953), .ZN(new_n571));
  NAND2_X1  g385(.A1(G234), .A2(G237), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT108), .ZN(new_n574));
  INV_X1    g388(.A(new_n262), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(G902), .A3(new_n572), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT21), .B(G898), .Z(new_n577));
  OAI21_X1  g391(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G478), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(KEYINPUT15), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(G122), .B1(new_n246), .B2(new_n247), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n582), .A2(KEYINPUT14), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT106), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(G122), .ZN(new_n585));
  INV_X1    g399(.A(G122), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(KEYINPUT106), .ZN(new_n587));
  OAI21_X1  g401(.A(G116), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n582), .B2(KEYINPUT14), .ZN(new_n589));
  OAI21_X1  g403(.A(G107), .B1(new_n583), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n211), .ZN(new_n591));
  XOR2_X1   g405(.A(G128), .B(G143), .Z(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n582), .A2(new_n588), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n590), .B(new_n593), .C1(G107), .C2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(G107), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n591), .B2(new_n592), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT13), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n190), .A3(G128), .ZN(new_n599));
  OAI211_X1 g413(.A(G134), .B(new_n599), .C1(new_n592), .C2(new_n598), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n600), .B(KEYINPUT107), .Z(new_n601));
  OAI21_X1  g415(.A(new_n595), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n317), .A2(G217), .A3(new_n406), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n581), .B1(new_n606), .B2(new_n303), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n303), .B(new_n581), .C1(new_n604), .C2(new_n605), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n548), .A2(new_n569), .A3(new_n578), .A4(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n401), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n453), .B1(new_n434), .B2(new_n451), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n459), .A2(new_n462), .A3(new_n452), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n611), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n314), .A2(new_n465), .A3(new_n513), .A4(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(new_n331), .Z(G3));
  NAND2_X1  g433(.A1(new_n301), .A2(new_n303), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n620), .A2(G472), .B1(new_n290), .B2(new_n301), .ZN(new_n621));
  INV_X1    g435(.A(new_n400), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n513), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n548), .A2(new_n569), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  OR3_X1    g439(.A1(new_n604), .A2(new_n605), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n625), .B1(new_n604), .B2(new_n605), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n579), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n579), .B(new_n303), .C1(new_n604), .C2(new_n605), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n579), .A2(new_n303), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n628), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n624), .A2(new_n632), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n401), .B(new_n578), .C1(new_n454), .C2(new_n463), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n623), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT34), .B(G104), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  INV_X1    g451(.A(new_n610), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n567), .B(KEYINPUT20), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n548), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n623), .A2(new_n634), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT35), .B(G107), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NAND2_X1  g457(.A1(new_n486), .A2(new_n494), .ZN(new_n644));
  INV_X1    g458(.A(new_n468), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n644), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n508), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n506), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n465), .A2(new_n617), .A3(new_n621), .A4(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  XNOR2_X1  g466(.A(new_n574), .B(KEYINPUT109), .ZN(new_n653));
  INV_X1    g467(.A(G900), .ZN(new_n654));
  INV_X1    g468(.A(new_n576), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n640), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n400), .B1(new_n506), .B2(new_n648), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n314), .A2(new_n615), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  XNOR2_X1  g474(.A(KEYINPUT111), .B(KEYINPUT39), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n656), .B(new_n661), .Z(new_n662));
  NOR2_X1   g476(.A1(new_n400), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT40), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n287), .B(G472), .C1(new_n297), .C2(new_n270), .ZN(new_n666));
  NAND2_X1  g480(.A1(G472), .A2(G902), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT110), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n292), .A2(new_n670), .A3(new_n302), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n624), .A2(new_n401), .A3(new_n638), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n613), .A2(new_n614), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT38), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n665), .A2(new_n671), .A3(new_n673), .A4(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n664), .A2(KEYINPUT40), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n676), .A2(new_n649), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n190), .ZN(G45));
  INV_X1    g493(.A(new_n656), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n543), .A2(KEYINPUT105), .A3(new_n303), .ZN(new_n681));
  AOI21_X1  g495(.A(KEYINPUT105), .B1(new_n543), .B2(new_n303), .ZN(new_n682));
  INV_X1    g496(.A(G475), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n565), .B1(new_n564), .B2(new_n559), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n555), .B1(new_n536), .B2(new_n538), .ZN(new_n686));
  INV_X1    g500(.A(new_n559), .ZN(new_n687));
  NOR4_X1   g501(.A1(new_n686), .A2(KEYINPUT103), .A3(new_n687), .A4(new_n560), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT20), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n557), .B2(new_n558), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n685), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n632), .B(new_n680), .C1(new_n684), .C2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n314), .A2(new_n615), .A3(new_n658), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT112), .B(G146), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G48));
  NOR2_X1   g510(.A1(new_n634), .A2(new_n633), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n323), .B1(new_n393), .B2(new_n366), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n386), .A2(new_n366), .A3(new_n323), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n303), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(G469), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n370), .A2(new_n387), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n396), .A3(new_n303), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n701), .A2(new_n319), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n314), .A2(new_n697), .A3(new_n513), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  INV_X1    g522(.A(new_n640), .ZN(new_n709));
  INV_X1    g523(.A(new_n578), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n512), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n464), .A2(new_n704), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n314), .A2(new_n709), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  INV_X1    g528(.A(new_n611), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n314), .A2(new_n715), .A3(new_n649), .A4(new_n712), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n716), .A2(KEYINPUT113), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(KEYINPUT113), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  NAND2_X1  g534(.A1(new_n287), .A2(KEYINPUT31), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT114), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n307), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n269), .B1(new_n307), .B2(new_n722), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n271), .B(new_n721), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n725), .A2(new_n290), .B1(G472), .B2(new_n620), .ZN(new_n726));
  INV_X1    g540(.A(new_n674), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n672), .A2(new_n727), .A3(new_n710), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n726), .A2(new_n728), .A3(new_n513), .A4(new_n705), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  NAND2_X1  g544(.A1(new_n692), .A2(KEYINPUT115), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n624), .A2(new_n732), .A3(new_n632), .A4(new_n680), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n726), .A2(new_n734), .A3(new_n649), .A4(new_n712), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  AND3_X1   g550(.A1(new_n301), .A2(KEYINPUT32), .A3(new_n290), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT32), .B1(new_n301), .B2(new_n290), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n512), .B1(new_n739), .B2(new_n313), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT116), .B1(new_n388), .B2(new_n399), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n703), .A2(new_n742), .A3(new_n398), .A4(new_n395), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n741), .A2(new_n743), .A3(new_n319), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n613), .A2(new_n614), .A3(new_n401), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n740), .A2(KEYINPUT42), .A3(new_n734), .A4(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n734), .A2(new_n314), .A3(new_n746), .A4(new_n513), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  NAND4_X1  g566(.A1(new_n314), .A2(new_n746), .A3(new_n513), .A4(new_n657), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G134), .ZN(G36));
  NOR2_X1   g568(.A1(new_n684), .A2(new_n691), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n632), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT43), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n758), .A3(new_n632), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n621), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n649), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n745), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n760), .A2(KEYINPUT44), .A3(new_n761), .A4(new_n649), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n391), .A2(new_n394), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n391), .A2(KEYINPUT45), .A3(new_n394), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(G469), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n398), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n703), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT46), .B1(new_n772), .B2(new_n398), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n319), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(new_n662), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n767), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(KEYINPUT117), .B(G137), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G39));
  AND2_X1   g594(.A1(new_n776), .A2(KEYINPUT47), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n782), .B(new_n319), .C1(new_n774), .C2(new_n775), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  OR3_X1    g598(.A1(new_n781), .A2(new_n692), .A3(new_n784), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n785), .A2(new_n314), .A3(new_n513), .A4(new_n745), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n479), .ZN(G42));
  AND2_X1   g601(.A1(new_n701), .A2(new_n703), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n789), .A2(KEYINPUT49), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(KEYINPUT49), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n513), .A3(new_n791), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n792), .A2(new_n612), .A3(new_n675), .ZN(new_n793));
  INV_X1    g607(.A(new_n671), .ZN(new_n794));
  INV_X1    g608(.A(new_n756), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n793), .A2(new_n319), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n726), .A2(new_n513), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n757), .A2(new_n653), .A3(new_n759), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n675), .A2(new_n401), .A3(new_n704), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(KEYINPUT119), .A2(KEYINPUT50), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n799), .B(new_n800), .C1(KEYINPUT119), .C2(KEYINPUT50), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI22_X1  g619(.A1(new_n781), .A2(new_n784), .B1(new_n319), .B2(new_n789), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n765), .A3(new_n799), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n725), .A2(new_n290), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n620), .A2(G472), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n808), .A2(new_n809), .A3(new_n649), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n757), .A2(new_n653), .A3(new_n759), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n745), .A2(new_n704), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n512), .A2(new_n574), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n794), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n815), .A2(new_n624), .A3(new_n632), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n805), .A2(new_n807), .A3(new_n813), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n811), .A2(new_n740), .A3(new_n812), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT121), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n811), .A2(new_n740), .A3(new_n823), .A4(new_n812), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT122), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n822), .A2(KEYINPUT122), .A3(new_n824), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(KEYINPUT48), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n816), .B1(new_n803), .B2(new_n804), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(KEYINPUT51), .A3(new_n813), .A4(new_n807), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n799), .A2(new_n712), .ZN(new_n831));
  INV_X1    g645(.A(new_n633), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n794), .A2(new_n832), .A3(new_n812), .A4(new_n814), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(new_n571), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT120), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n831), .A2(new_n836), .A3(new_n571), .A4(new_n833), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT48), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n835), .A2(new_n837), .B1(new_n825), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n820), .A2(new_n828), .A3(new_n830), .A4(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n618), .A2(new_n650), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n633), .B1(new_n610), .B2(new_n624), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n464), .A2(KEYINPUT97), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n615), .A2(new_n616), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n578), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n623), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n610), .A2(new_n548), .A3(new_n639), .A4(new_n680), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n314), .A2(new_n658), .A3(new_n765), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n753), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n751), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n706), .A2(new_n713), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n716), .A2(KEYINPUT113), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n716), .A2(KEYINPUT113), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n854), .B(new_n729), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n810), .A2(new_n858), .A3(new_n734), .A4(new_n746), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n734), .A2(new_n746), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n808), .A2(new_n809), .A3(new_n649), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT118), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n853), .A2(new_n857), .A3(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n659), .A2(new_n694), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n744), .A2(new_n727), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n649), .A2(new_n656), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n671), .A2(new_n867), .A3(new_n673), .A4(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n865), .A2(new_n866), .A3(new_n735), .A4(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n735), .A2(new_n869), .A3(new_n659), .A4(new_n694), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT52), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT53), .B1(new_n864), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n729), .A2(new_n706), .A3(new_n713), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n717), .B2(new_n718), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n851), .A2(new_n842), .A3(new_n847), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n859), .A2(new_n862), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n877), .A2(new_n751), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n880), .A2(new_n881), .A3(new_n873), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n841), .B1(new_n875), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n864), .A2(KEYINPUT53), .A3(new_n874), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n881), .B1(new_n880), .B2(new_n873), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT54), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n840), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n570), .A2(new_n406), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT123), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n796), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(KEYINPUT124), .B(new_n796), .C1(new_n887), .C2(new_n889), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(G75));
  AOI21_X1  g708(.A(new_n303), .B1(new_n884), .B2(new_n885), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(G210), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n456), .A2(new_n458), .A3(new_n455), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n434), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT55), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n896), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n896), .B2(new_n897), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n262), .A2(G952), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(G51));
  NAND2_X1  g718(.A1(new_n398), .A2(KEYINPUT57), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n883), .A2(new_n886), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n398), .A2(KEYINPUT57), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n702), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n895), .A2(G469), .A3(new_n770), .A4(new_n771), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(G54));
  NAND3_X1  g724(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n911), .A2(new_n686), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n686), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n912), .A2(new_n913), .A3(new_n903), .ZN(G60));
  XOR2_X1   g728(.A(new_n631), .B(KEYINPUT59), .Z(new_n915));
  NAND3_X1  g729(.A1(new_n883), .A2(new_n886), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n626), .A2(new_n627), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n916), .A2(KEYINPUT125), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n903), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n916), .B2(new_n917), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT125), .B1(new_n916), .B2(new_n917), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n918), .A2(new_n920), .A3(new_n921), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n884), .B2(new_n885), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n925), .A2(new_n502), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n903), .B1(new_n925), .B2(new_n647), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n926), .A2(KEYINPUT61), .A3(new_n927), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(G66));
  AOI21_X1  g746(.A(new_n406), .B1(new_n577), .B2(G224), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n877), .A2(new_n848), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n934), .B2(new_n262), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n426), .B(new_n433), .C1(G898), .C2(new_n262), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n935), .B(new_n936), .Z(G69));
  AOI21_X1  g751(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT127), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n550), .A2(new_n552), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n238), .B(new_n940), .Z(new_n941));
  NAND2_X1  g755(.A1(new_n575), .A2(G900), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n865), .A2(new_n735), .A3(new_n753), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n786), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n672), .A2(new_n727), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n740), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n767), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n777), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n944), .A2(new_n949), .A3(new_n751), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n941), .B(new_n942), .C1(new_n950), .C2(new_n575), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n939), .B1(new_n951), .B2(KEYINPUT126), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n865), .A2(new_n735), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(new_n678), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n786), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n740), .A2(new_n663), .A3(new_n765), .A4(new_n843), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n778), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n575), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n951), .B1(new_n960), .B2(new_n941), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n952), .A2(new_n961), .ZN(new_n962));
  OAI221_X1 g776(.A(new_n951), .B1(KEYINPUT126), .B2(new_n939), .C1(new_n960), .C2(new_n941), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(G72));
  XOR2_X1   g778(.A(new_n667), .B(KEYINPUT63), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n957), .A2(new_n959), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(new_n934), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n260), .A2(new_n269), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n965), .B1(new_n950), .B2(new_n934), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n970), .A2(new_n269), .A3(new_n260), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n884), .A2(new_n885), .ZN(new_n972));
  INV_X1    g786(.A(new_n968), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n972), .A2(new_n311), .A3(new_n965), .A4(new_n973), .ZN(new_n974));
  AND4_X1   g788(.A1(new_n919), .A2(new_n969), .A3(new_n971), .A4(new_n974), .ZN(G57));
endmodule


