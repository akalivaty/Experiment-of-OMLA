//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995;
  INV_X1    g000(.A(G197gat), .ZN(new_n202));
  INV_X1    g001(.A(G204gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  NAND2_X1  g005(.A1(G211gat), .A2(G218gat), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(G211gat), .A2(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT72), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(new_n207), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n210), .B1(new_n209), .B2(new_n207), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n208), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT73), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n204), .A2(new_n205), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n207), .A2(new_n206), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G211gat), .B(G218gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT72), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n220), .A3(new_n211), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n214), .A2(new_n215), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n218), .A2(new_n220), .A3(KEYINPUT73), .A4(new_n211), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT2), .ZN(new_n229));
  OR2_X1    g028(.A1(G141gat), .A2(G148gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT75), .ZN(new_n233));
  AND2_X1   g032(.A1(G155gat), .A2(G162gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G155gat), .ZN(new_n237));
  INV_X1    g036(.A(G162gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(KEYINPUT75), .A3(new_n228), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n232), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n234), .A2(new_n235), .ZN(new_n242));
  AND2_X1   g041(.A1(G141gat), .A2(G148gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(G141gat), .A2(G148gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n242), .A2(new_n245), .A3(KEYINPUT75), .A4(new_n229), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n227), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT76), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n250), .B1(new_n247), .B2(new_n226), .ZN(new_n251));
  AOI211_X1 g050(.A(KEYINPUT76), .B(KEYINPUT3), .C1(new_n241), .C2(new_n246), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n223), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n222), .A2(new_n224), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G228gat), .A2(G233gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n249), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT82), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n253), .A2(KEYINPUT82), .A3(new_n254), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n214), .A2(new_n221), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n223), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n247), .B1(new_n263), .B2(new_n226), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n260), .A2(new_n261), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n258), .B1(new_n266), .B2(new_n256), .ZN(new_n267));
  INV_X1    g066(.A(G22gat), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT85), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT85), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT82), .B1(new_n253), .B2(new_n254), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(new_n264), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n257), .B1(new_n272), .B2(new_n261), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n270), .B(G22gat), .C1(new_n273), .C2(new_n258), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT86), .ZN(new_n276));
  XOR2_X1   g075(.A(KEYINPUT83), .B(G22gat), .Z(new_n277));
  NAND3_X1  g076(.A1(new_n267), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G78gat), .B(G106gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT31), .B(G50gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  NAND3_X1  g080(.A1(new_n249), .A2(new_n255), .A3(new_n257), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n253), .A2(KEYINPUT82), .A3(new_n254), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n283), .A2(new_n271), .A3(new_n264), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n277), .B(new_n282), .C1(new_n284), .C2(new_n257), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n281), .B1(new_n285), .B2(KEYINPUT86), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n275), .A2(new_n278), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT84), .ZN(new_n288));
  INV_X1    g087(.A(new_n277), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(new_n273), .B2(new_n258), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n285), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n281), .B(KEYINPUT81), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n288), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  AOI211_X1 g093(.A(KEYINPUT84), .B(new_n292), .C1(new_n290), .C2(new_n285), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n287), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  NAND2_X1  g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G183gat), .ZN(new_n302));
  INV_X1    g101(.A(G190gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT24), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  OR2_X1    g106(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n302), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT23), .ZN(new_n313));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(G169gat), .B2(G176gat), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n311), .A2(KEYINPUT25), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n304), .A2(new_n306), .B1(new_n302), .B2(new_n303), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(G169gat), .B2(G176gat), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n312), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(KEYINPUT65), .B(G190gat), .Z(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT27), .B(G183gat), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n328), .A2(KEYINPUT28), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT28), .B1(new_n328), .B2(new_n329), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n327), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n301), .B1(new_n333), .B2(new_n223), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n300), .B1(new_n323), .B2(new_n332), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n254), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n329), .A2(new_n308), .A3(new_n309), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n328), .A2(KEYINPUT28), .A3(new_n329), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n341), .A2(new_n327), .B1(new_n318), .B2(new_n322), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n300), .B1(new_n342), .B2(KEYINPUT29), .ZN(new_n343));
  INV_X1    g142(.A(new_n254), .ZN(new_n344));
  INV_X1    g143(.A(new_n335), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n299), .B1(new_n336), .B2(new_n346), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n334), .A2(new_n254), .A3(new_n335), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n344), .B1(new_n343), .B2(new_n345), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n299), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT30), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n347), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n336), .A2(new_n346), .A3(KEYINPUT30), .A4(new_n299), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n354), .A2(new_n355), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n353), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT5), .ZN(new_n359));
  AND2_X1   g158(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n361));
  INV_X1    g160(.A(G120gat), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(G113gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT69), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT69), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT68), .B(G113gat), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n367), .B(new_n364), .C1(new_n368), .C2(new_n362), .ZN(new_n369));
  XOR2_X1   g168(.A(G127gat), .B(G134gat), .Z(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(KEYINPUT1), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n366), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT66), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G127gat), .B(G134gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT66), .ZN(new_n376));
  INV_X1    g175(.A(G113gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G120gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n364), .A2(new_n378), .A3(KEYINPUT67), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT67), .B1(new_n364), .B2(new_n378), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n374), .B(new_n376), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n372), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n248), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n372), .A2(new_n383), .A3(new_n247), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n359), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n384), .B(new_n391), .C1(new_n251), .C2(new_n252), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n386), .A2(KEYINPUT4), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n392), .B(new_n388), .C1(KEYINPUT77), .C2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n372), .A2(new_n383), .A3(new_n395), .A4(new_n247), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n393), .A2(KEYINPUT77), .A3(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n390), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT0), .ZN(new_n400));
  XNOR2_X1  g199(.A(G57gat), .B(G85gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  NAND3_X1  g201(.A1(new_n393), .A2(KEYINPUT78), .A3(new_n396), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT78), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n404), .A3(KEYINPUT4), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n392), .A2(new_n359), .A3(new_n388), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT79), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n405), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT79), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n410), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n398), .B(new_n402), .C1(new_n409), .C2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT80), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n398), .B1(new_n409), .B2(new_n412), .ZN(new_n416));
  INV_X1    g215(.A(new_n402), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n406), .A2(new_n408), .A3(KEYINPUT79), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n411), .B1(new_n410), .B2(new_n407), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n422), .A2(KEYINPUT80), .A3(new_n402), .A4(new_n398), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n415), .A2(new_n418), .A3(new_n419), .A4(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n416), .A2(KEYINPUT6), .A3(new_n417), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n358), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n333), .A2(new_n372), .A3(new_n383), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n342), .A2(new_n384), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT32), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(new_n429), .B2(new_n430), .ZN(new_n433));
  XOR2_X1   g232(.A(G15gat), .B(G43gat), .Z(new_n434));
  XNOR2_X1  g233(.A(G71gat), .B(G99gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n436), .ZN(new_n439));
  OAI221_X1 g238(.A(KEYINPUT32), .B1(new_n432), .B2(new_n439), .C1(new_n429), .C2(new_n430), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT34), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n429), .A2(KEYINPUT70), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n429), .A2(KEYINPUT70), .B1(G227gat), .B2(G233gat), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n442), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT71), .B1(new_n429), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n429), .A2(KEYINPUT71), .A3(new_n447), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI22_X1  g250(.A1(new_n438), .A2(new_n441), .B1(new_n445), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n443), .A2(new_n444), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT34), .ZN(new_n455));
  INV_X1    g254(.A(new_n450), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(new_n448), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n455), .A2(new_n457), .A3(new_n437), .A4(new_n440), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n296), .A2(new_n426), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT35), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n452), .A2(new_n458), .A3(KEYINPUT90), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT90), .B1(new_n452), .B2(new_n458), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n402), .B(KEYINPUT87), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n416), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n415), .A2(new_n469), .A3(new_n419), .A4(new_n423), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n425), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT35), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n353), .B(new_n472), .C1(new_n356), .C2(new_n357), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n466), .A2(new_n296), .A3(new_n471), .A4(new_n474), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n452), .A2(new_n458), .A3(KEYINPUT36), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT36), .B1(new_n452), .B2(new_n458), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n424), .A2(new_n425), .ZN(new_n479));
  INV_X1    g278(.A(new_n358), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n273), .A2(new_n289), .A3(new_n258), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n266), .A2(new_n256), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n277), .B1(new_n483), .B2(new_n282), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n293), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT84), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n291), .A2(new_n288), .A3(new_n293), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n285), .A2(KEYINPUT86), .ZN(new_n488));
  INV_X1    g287(.A(new_n281), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n488), .A2(new_n489), .A3(new_n278), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n486), .A2(new_n487), .B1(new_n490), .B2(new_n275), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n478), .B1(new_n481), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT37), .B1(new_n348), .B2(new_n349), .ZN(new_n493));
  INV_X1    g292(.A(new_n299), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n494), .A2(KEYINPUT37), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n493), .B1(new_n347), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT89), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT38), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n497), .B1(new_n496), .B2(KEYINPUT38), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n343), .A2(new_n500), .A3(new_n345), .A4(new_n344), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT37), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n502), .B1(new_n350), .B2(KEYINPUT88), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT38), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n336), .A2(new_n346), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n504), .B(new_n494), .C1(new_n505), .C2(KEYINPUT37), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n351), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n498), .A2(new_n499), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(new_n425), .A3(new_n470), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n406), .A2(new_n392), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n389), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n467), .B1(new_n511), .B2(KEYINPUT39), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT40), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT39), .B1(new_n387), .B2(new_n389), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n514), .B1(new_n510), .B2(new_n389), .ZN(new_n515));
  OR3_X1    g314(.A1(new_n512), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n513), .B1(new_n512), .B2(new_n515), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n516), .A2(new_n469), .A3(new_n517), .A4(new_n358), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n296), .A2(new_n509), .A3(new_n518), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n462), .A2(new_n475), .B1(new_n492), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT92), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(G1gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT16), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT93), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n521), .A2(new_n522), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n521), .A2(new_n522), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n524), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT94), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G8gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT93), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n523), .A2(new_n534), .A3(new_n525), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n528), .A2(new_n531), .A3(new_n524), .A4(new_n529), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n527), .A2(new_n533), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(G8gat), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n526), .A2(new_n530), .A3(new_n532), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NOR3_X1   g341(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n543));
  INV_X1    g342(.A(G29gat), .ZN(new_n544));
  INV_X1    g343(.A(G36gat), .ZN(new_n545));
  OAI22_X1  g344(.A1(new_n542), .A2(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G43gat), .B(G50gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(KEYINPUT15), .A3(new_n547), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n547), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(KEYINPUT15), .B2(new_n547), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n543), .A2(KEYINPUT91), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n543), .A2(KEYINPUT91), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n542), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n548), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT17), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n556), .B(new_n548), .C1(new_n550), .C2(new_n553), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n538), .A2(new_n540), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n539), .B1(new_n537), .B2(G8gat), .ZN(new_n561));
  INV_X1    g360(.A(new_n554), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n559), .B(new_n560), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT18), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n560), .B(KEYINPUT13), .Z(new_n565));
  AOI21_X1  g364(.A(new_n562), .B1(new_n538), .B2(new_n540), .ZN(new_n566));
  AOI211_X1 g365(.A(new_n554), .B(new_n539), .C1(new_n537), .C2(G8gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT95), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g369(.A(KEYINPUT95), .B(new_n565), .C1(new_n566), .C2(new_n567), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n564), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(G197gat), .ZN(new_n575));
  XOR2_X1   g374(.A(KEYINPUT11), .B(G169gat), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(KEYINPUT12), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT18), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n566), .B1(new_n561), .B2(new_n558), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(KEYINPUT18), .A3(new_n560), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n572), .A2(new_n580), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n579), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n520), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n479), .ZN(new_n589));
  XNOR2_X1  g388(.A(G190gat), .B(G218gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT98), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT97), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT7), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT7), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT97), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n594), .A2(new_n596), .A3(G85gat), .A4(G92gat), .ZN(new_n597));
  INV_X1    g396(.A(G99gat), .ZN(new_n598));
  INV_X1    g397(.A(G106gat), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT8), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(G85gat), .A2(G92gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(G85gat), .A2(G92gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(KEYINPUT97), .A3(new_n595), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n597), .A2(new_n600), .A3(new_n601), .A4(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G99gat), .B(G106gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n558), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n606), .ZN(new_n608));
  AND2_X1   g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n608), .A2(new_n554), .B1(KEYINPUT41), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n592), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n609), .A2(KEYINPUT41), .ZN(new_n613));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n607), .A2(new_n592), .A3(new_n610), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n612), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n612), .B2(new_n616), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G57gat), .B(G64gat), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(G71gat), .A2(G78gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(G71gat), .A2(G78gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT96), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(KEYINPUT96), .A3(new_n624), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n622), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n625), .B(new_n626), .C1(new_n620), .C2(new_n621), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT21), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n561), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n629), .A2(new_n630), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT21), .ZN(new_n635));
  NAND2_X1  g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  OAI211_X1 g436(.A(G231gat), .B(G233gat), .C1(new_n631), .C2(KEYINPUT21), .ZN(new_n638));
  INV_X1    g437(.A(G127gat), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n639), .B1(new_n637), .B2(new_n638), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n633), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n561), .B(new_n632), .C1(new_n640), .C2(new_n641), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(new_n237), .ZN(new_n646));
  XNOR2_X1  g445(.A(G183gat), .B(G211gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  AND3_X1   g447(.A1(new_n643), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n643), .B2(new_n644), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT99), .B1(new_n619), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n651), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n617), .A2(new_n618), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(G120gat), .B(G148gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT101), .ZN(new_n658));
  XNOR2_X1  g457(.A(G176gat), .B(G204gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n658), .B(new_n659), .Z(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(G230gat), .ZN(new_n662));
  INV_X1    g461(.A(G233gat), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n606), .A2(new_n634), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT10), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n604), .A2(new_n605), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n604), .A2(new_n605), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n631), .A3(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n665), .A2(KEYINPUT100), .A3(new_n666), .A4(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n608), .A2(KEYINPUT10), .A3(new_n631), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n665), .A2(new_n666), .A3(new_n669), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n664), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n665), .A2(new_n669), .ZN(new_n678));
  INV_X1    g477(.A(new_n664), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n661), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n674), .A2(new_n675), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n679), .B1(new_n682), .B2(new_n672), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n683), .B(new_n660), .C1(new_n679), .C2(new_n678), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(KEYINPUT102), .B(new_n661), .C1(new_n677), .C2(new_n680), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n652), .A2(new_n656), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n588), .A2(new_n589), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G1gat), .ZN(G1324gat));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n588), .A2(new_n358), .A3(new_n690), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT16), .B(G8gat), .Z(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n693), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n694), .A2(new_n696), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(G8gat), .B2(new_n694), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n699), .B2(new_n693), .ZN(G1325gat));
  NAND2_X1  g499(.A1(new_n588), .A2(new_n690), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n476), .A2(new_n477), .ZN(new_n702));
  OAI21_X1  g501(.A(G15gat), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(G15gat), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n588), .A2(new_n704), .A3(new_n466), .A4(new_n690), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT103), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT103), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n703), .A2(new_n708), .A3(new_n705), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(G1326gat));
  NOR2_X1   g509(.A1(new_n701), .A2(new_n296), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT43), .B(G22gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  NAND2_X1  g512(.A1(new_n462), .A2(new_n475), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n492), .A2(new_n519), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n655), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n688), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n587), .A2(new_n653), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n479), .A2(G29gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(KEYINPUT45), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n723));
  INV_X1    g522(.A(new_n721), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n719), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n520), .B2(new_n655), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n474), .B1(new_n464), .B2(new_n465), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n491), .A2(new_n728), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n729), .A2(new_n471), .B1(new_n461), .B2(KEYINPUT35), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n296), .A2(new_n509), .A3(new_n518), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n702), .B1(new_n296), .B2(new_n426), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g532(.A(KEYINPUT44), .B(new_n619), .C1(new_n730), .C2(new_n733), .ZN(new_n734));
  AND4_X1   g533(.A1(new_n589), .A2(new_n727), .A3(new_n718), .A4(new_n734), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n722), .B(new_n725), .C1(new_n735), .C2(new_n544), .ZN(G1328gat));
  NOR2_X1   g535(.A1(new_n480), .A2(G36gat), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  OR3_X1    g537(.A1(new_n719), .A2(KEYINPUT46), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT46), .B1(new_n719), .B2(new_n738), .ZN(new_n740));
  AND4_X1   g539(.A1(new_n358), .A2(new_n727), .A3(new_n718), .A4(new_n734), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n739), .B(new_n740), .C1(new_n741), .C2(new_n545), .ZN(G1329gat));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n718), .A3(new_n734), .ZN(new_n743));
  OAI21_X1  g542(.A(G43gat), .B1(new_n743), .B2(new_n702), .ZN(new_n744));
  INV_X1    g543(.A(G43gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n720), .A2(new_n745), .A3(new_n466), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n744), .A2(KEYINPUT47), .A3(new_n746), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(G1330gat));
  OR3_X1    g550(.A1(new_n719), .A2(G50gat), .A3(new_n296), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n727), .A2(new_n491), .A3(new_n734), .A4(new_n718), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G50gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT48), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n752), .A2(new_n754), .A3(KEYINPUT48), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1331gat));
  NAND4_X1  g558(.A1(new_n587), .A2(new_n652), .A3(new_n656), .A4(new_n717), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT104), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n714), .A2(new_n715), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n479), .B(KEYINPUT105), .Z(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g566(.A(new_n480), .B(new_n763), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n768));
  NOR2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1333gat));
  NAND3_X1  g569(.A1(new_n761), .A2(new_n762), .A3(new_n466), .ZN(new_n771));
  AOI21_X1  g570(.A(G71gat), .B1(new_n771), .B2(KEYINPUT106), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n761), .A2(new_n762), .A3(new_n773), .A4(new_n466), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n764), .A2(G71gat), .A3(new_n478), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT50), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n775), .A2(new_n779), .A3(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1334gat));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n491), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g582(.A1(new_n587), .A2(new_n651), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n688), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n727), .A2(new_n734), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786), .B2(new_n479), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n479), .A2(G85gat), .A3(new_n688), .ZN(new_n788));
  INV_X1    g587(.A(new_n784), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT51), .B1(new_n716), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  NOR4_X1   g590(.A1(new_n520), .A2(new_n791), .A3(new_n655), .A4(new_n784), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n788), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n787), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n787), .A2(new_n793), .A3(KEYINPUT107), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(G1336gat));
  NAND4_X1  g597(.A1(new_n727), .A2(new_n358), .A3(new_n734), .A4(new_n785), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G92gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n688), .A2(new_n480), .A3(G92gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n790), .B2(new_n792), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n802), .A3(KEYINPUT108), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT52), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n800), .A2(new_n802), .A3(KEYINPUT108), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1337gat));
  OAI21_X1  g606(.A(G99gat), .B1(new_n786), .B2(new_n702), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n466), .A2(new_n598), .A3(new_n717), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT109), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n790), .B2(new_n792), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(G1338gat));
  NAND4_X1  g611(.A1(new_n727), .A2(new_n491), .A3(new_n734), .A4(new_n785), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G106gat), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n491), .A2(new_n599), .A3(new_n717), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n790), .B2(new_n792), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(new_n817), .A3(KEYINPUT110), .ZN(new_n818));
  XNOR2_X1  g617(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n814), .A2(new_n817), .A3(KEYINPUT110), .A4(new_n819), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1339gat));
  NOR2_X1   g622(.A1(new_n689), .A2(new_n586), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n583), .A2(new_n560), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n566), .A2(new_n567), .A3(new_n565), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n577), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n585), .A2(new_n687), .A3(new_n686), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n655), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n676), .A2(new_n664), .A3(new_n671), .A4(new_n670), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n683), .A2(KEYINPUT54), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n833), .B(new_n679), .C1(new_n682), .C2(new_n672), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n832), .A2(KEYINPUT55), .A3(new_n661), .A4(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n835), .A2(new_n684), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n832), .A2(new_n661), .A3(new_n834), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n579), .A2(new_n585), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n830), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n837), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n585), .A2(new_n841), .A3(new_n828), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n835), .A2(new_n684), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n619), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n651), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n825), .B1(new_n840), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n296), .A2(new_n460), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n847), .A3(new_n765), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT113), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n846), .A2(new_n850), .A3(new_n847), .A4(new_n765), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n480), .A3(new_n851), .ZN(new_n852));
  OR3_X1    g651(.A1(new_n852), .A2(new_n368), .A3(new_n587), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n466), .A2(new_n296), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n479), .A2(new_n358), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(G113gat), .B1(new_n857), .B2(new_n587), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n853), .B1(new_n860), .B2(new_n861), .ZN(G1340gat));
  NAND4_X1  g661(.A1(new_n849), .A2(new_n480), .A3(new_n717), .A4(new_n851), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n362), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n855), .A2(G120gat), .A3(new_n717), .A4(new_n856), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n864), .A2(KEYINPUT114), .A3(new_n865), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1341gat));
  NAND4_X1  g669(.A1(new_n855), .A2(G127gat), .A3(new_n653), .A4(new_n856), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT115), .Z(new_n872));
  INV_X1    g671(.A(new_n852), .ZN(new_n873));
  AOI21_X1  g672(.A(G127gat), .B1(new_n873), .B2(new_n653), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n874), .ZN(G1342gat));
  INV_X1    g674(.A(G134gat), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n619), .A2(new_n876), .ZN(new_n877));
  OR3_X1    g676(.A1(new_n852), .A2(KEYINPUT56), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G134gat), .B1(new_n857), .B2(new_n655), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT56), .B1(new_n852), .B2(new_n877), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G1343gat));
  NAND2_X1  g680(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n882));
  OR2_X1    g681(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n846), .A2(new_n491), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n585), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n580), .B1(new_n564), .B2(new_n572), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n836), .B(new_n841), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n655), .A3(new_n829), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n836), .A2(new_n585), .A3(new_n841), .A4(new_n828), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n653), .B1(new_n889), .B2(new_n619), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n824), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g690(.A(KEYINPUT116), .B(KEYINPUT57), .C1(new_n891), .C2(new_n296), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n478), .A2(new_n479), .A3(new_n358), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n884), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G141gat), .B1(new_n894), .B2(new_n587), .ZN(new_n895));
  OR2_X1    g694(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n846), .A2(new_n765), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n491), .A2(new_n702), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n898), .A2(KEYINPUT117), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(KEYINPUT117), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n480), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n587), .A2(G141gat), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n902), .A2(new_n903), .B1(KEYINPUT118), .B2(KEYINPUT58), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n895), .A2(new_n896), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n896), .B1(new_n895), .B2(new_n904), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(G1344gat));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT57), .B1(new_n491), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(new_n846), .B2(new_n491), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n891), .A2(new_n909), .A3(new_n296), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n893), .A2(new_n717), .ZN(new_n914));
  OAI211_X1 g713(.A(KEYINPUT59), .B(G148gat), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n884), .A2(new_n892), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n893), .A2(new_n917), .A3(new_n717), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n902), .B2(new_n717), .ZN(new_n919));
  OAI221_X1 g718(.A(new_n915), .B1(new_n916), .B2(new_n918), .C1(G148gat), .C2(new_n919), .ZN(G1345gat));
  OAI21_X1  g719(.A(G155gat), .B1(new_n894), .B2(new_n651), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n902), .A2(new_n237), .A3(new_n653), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1346gat));
  NOR3_X1   g722(.A1(new_n894), .A2(new_n238), .A3(new_n655), .ZN(new_n924));
  AOI21_X1  g723(.A(G162gat), .B1(new_n902), .B2(new_n619), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n765), .A2(new_n480), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n855), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(G169gat), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n928), .A2(new_n929), .A3(new_n587), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n846), .A2(KEYINPUT120), .A3(new_n479), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT120), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n932), .B1(new_n891), .B2(new_n589), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n847), .A2(new_n358), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n586), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n930), .B1(new_n937), .B2(new_n929), .ZN(G1348gat));
  INV_X1    g737(.A(G176gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n936), .A2(new_n939), .A3(new_n717), .ZN(new_n940));
  OAI21_X1  g739(.A(G176gat), .B1(new_n928), .B2(new_n688), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1349gat));
  NAND4_X1  g741(.A1(new_n934), .A2(new_n329), .A3(new_n653), .A4(new_n935), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n927), .A2(new_n846), .A3(new_n653), .A4(new_n854), .ZN(new_n944));
  AOI22_X1  g743(.A1(new_n944), .A2(G183gat), .B1(KEYINPUT121), .B2(KEYINPUT60), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g745(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n946), .B(new_n947), .ZN(G1350gat));
  NAND3_X1  g747(.A1(new_n855), .A2(new_n619), .A3(new_n927), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT123), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n949), .A2(G190gat), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n951), .B1(new_n949), .B2(G190gat), .ZN(new_n953));
  OAI22_X1  g752(.A1(new_n952), .A2(new_n953), .B1(KEYINPUT123), .B2(new_n950), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n619), .A2(new_n328), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n936), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n955), .B1(new_n936), .B2(new_n956), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G1351gat));
  INV_X1    g758(.A(new_n898), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n934), .A2(new_n358), .A3(new_n586), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n927), .A2(new_n702), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n846), .A2(new_n491), .A3(new_n910), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n909), .B1(new_n891), .B2(new_n296), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n587), .A2(new_n202), .ZN(new_n966));
  AOI22_X1  g765(.A1(new_n961), .A2(new_n202), .B1(new_n965), .B2(new_n966), .ZN(G1352gat));
  AOI21_X1  g766(.A(new_n203), .B1(new_n965), .B2(new_n717), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n688), .A2(new_n480), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n934), .A2(new_n203), .A3(new_n969), .A4(new_n960), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n971), .A2(KEYINPUT124), .A3(new_n972), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT124), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n975), .B1(new_n970), .B2(KEYINPUT62), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n974), .B2(new_n976), .ZN(G1353gat));
  NOR3_X1   g776(.A1(new_n765), .A2(new_n480), .A3(new_n478), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n653), .B(new_n978), .C1(new_n911), .C2(new_n912), .ZN(new_n979));
  NAND2_X1  g778(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n979), .A2(G211gat), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n980), .B1(new_n979), .B2(G211gat), .ZN(new_n982));
  OAI22_X1  g781(.A1(new_n981), .A2(new_n982), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n651), .A2(G211gat), .ZN(new_n984));
  NAND4_X1  g783(.A1(new_n934), .A2(new_n358), .A3(new_n960), .A4(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT125), .ZN(new_n986));
  XNOR2_X1  g785(.A(new_n985), .B(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n983), .A2(new_n987), .ZN(G1354gat));
  NAND4_X1  g787(.A1(new_n934), .A2(new_n358), .A3(new_n619), .A4(new_n960), .ZN(new_n989));
  INV_X1    g788(.A(G218gat), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n989), .A2(KEYINPUT127), .A3(new_n990), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n655), .A2(new_n990), .ZN(new_n995));
  AOI22_X1  g794(.A1(new_n993), .A2(new_n994), .B1(new_n965), .B2(new_n995), .ZN(G1355gat));
endmodule


