//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004;
  INV_X1    g000(.A(G141gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G148gat), .ZN(new_n203));
  INV_X1    g002(.A(G148gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G141gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT77), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n206), .A2(new_n207), .B1(KEYINPUT2), .B2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT77), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n208), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT76), .B1(G155gat), .B2(G162gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n211), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n214), .A2(new_n208), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT79), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT78), .B1(new_n202), .B2(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT78), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(new_n204), .A3(G141gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n228), .A3(new_n203), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT79), .A3(new_n208), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n224), .A2(new_n225), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n220), .A2(new_n221), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n231), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n218), .B1(new_n209), .B2(new_n210), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT3), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G113gat), .B(G120gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n237));
  XOR2_X1   g036(.A(G127gat), .B(G134gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n232), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G225gat), .A2(G233gat), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n242), .B(KEYINPUT80), .Z(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n220), .A2(KEYINPUT81), .A3(new_n231), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT81), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(new_n233), .B2(new_n234), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(KEYINPUT4), .A3(new_n239), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n233), .A2(new_n234), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n239), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n245), .A2(new_n250), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT5), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n251), .B(new_n239), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(new_n243), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n252), .A2(KEYINPUT4), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n246), .A2(new_n248), .A3(new_n253), .A4(new_n239), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT82), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n241), .A2(new_n256), .A3(new_n244), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n264), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n260), .A2(new_n261), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT82), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n259), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G1gat), .B(G29gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT0), .ZN(new_n271));
  XNOR2_X1  g070(.A(G57gat), .B(G85gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n269), .A2(KEYINPUT6), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(new_n269), .B2(new_n274), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n263), .B1(new_n262), .B2(new_n264), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n266), .A2(KEYINPUT82), .A3(new_n267), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n278), .A2(new_n279), .B1(new_n255), .B2(new_n258), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(new_n273), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n275), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT75), .ZN(new_n283));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n286), .A2(KEYINPUT64), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(KEYINPUT64), .ZN(new_n288));
  NAND3_X1  g087(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(G183gat), .B2(G190gat), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n287), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G169gat), .ZN(new_n292));
  INV_X1    g091(.A(G176gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT23), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(G169gat), .B2(G176gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n291), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n285), .B1(new_n299), .B2(KEYINPUT25), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301));
  OAI211_X1 g100(.A(KEYINPUT65), .B(new_n301), .C1(new_n291), .C2(new_n298), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n286), .A2(new_n303), .ZN(new_n304));
  OR2_X1    g103(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(G183gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n286), .A2(new_n303), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n304), .A2(new_n289), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n298), .A2(new_n301), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT68), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT68), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n314), .A3(new_n311), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n300), .A2(new_n302), .A3(new_n313), .A4(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n305), .A2(new_n307), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT27), .B(G183gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT69), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(KEYINPUT69), .A3(KEYINPUT28), .ZN(new_n323));
  NOR2_X1   g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(KEYINPUT26), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n297), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n324), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n322), .A2(new_n323), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n284), .B1(new_n316), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G197gat), .B(G204gat), .ZN(new_n331));
  INV_X1    g130(.A(G211gat), .ZN(new_n332));
  INV_X1    g131(.A(G218gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n331), .B1(KEYINPUT22), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G211gat), .B(G218gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT73), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n334), .A2(KEYINPUT22), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n339), .A2(new_n340), .A3(new_n336), .A4(new_n331), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n336), .A2(KEYINPUT72), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n336), .A2(KEYINPUT72), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n335), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT29), .B1(new_n316), .B2(new_n328), .ZN(new_n347));
  INV_X1    g146(.A(new_n284), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n330), .B(new_n346), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n313), .A2(new_n302), .A3(new_n315), .ZN(new_n350));
  OR3_X1    g149(.A1(new_n287), .A2(new_n288), .A3(new_n290), .ZN(new_n351));
  INV_X1    g150(.A(new_n298), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT65), .B1(new_n353), .B2(new_n301), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n328), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n348), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT74), .B1(new_n357), .B2(new_n329), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(new_n347), .B2(new_n348), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n283), .B(new_n349), .C1(new_n361), .C2(new_n346), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n346), .B1(new_n358), .B2(new_n360), .ZN(new_n363));
  INV_X1    g162(.A(new_n349), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT75), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G8gat), .B(G36gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(G64gat), .B(G92gat), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n366), .B(new_n367), .Z(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n362), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT30), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n363), .A2(new_n364), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(new_n368), .ZN(new_n373));
  NOR4_X1   g172(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT30), .A4(new_n369), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n282), .B(new_n370), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G228gat), .A2(G233gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n338), .A2(KEYINPUT83), .A3(new_n341), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n335), .A2(new_n337), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT83), .B1(new_n338), .B2(new_n341), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n356), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n249), .B1(new_n221), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n232), .A2(new_n356), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT84), .ZN(new_n384));
  INV_X1    g183(.A(new_n346), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n376), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n251), .A2(new_n376), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT29), .B1(new_n342), .B2(new_n345), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT85), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n221), .B1(new_n390), .B2(new_n391), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n383), .A2(new_n385), .B1(new_n384), .B2(new_n376), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(KEYINPUT87), .A2(G22gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n388), .A2(new_n396), .A3(new_n398), .ZN(new_n401));
  XNOR2_X1  g200(.A(G78gat), .B(G106gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT31), .B(G50gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n400), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  OR2_X1    g205(.A1(KEYINPUT86), .A2(G22gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(KEYINPUT86), .A2(G22gat), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n388), .A2(new_n396), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n381), .A2(new_n221), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n386), .B1(new_n410), .B2(new_n249), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n411), .A2(new_n376), .B1(new_n394), .B2(new_n395), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n409), .B(new_n404), .C1(new_n412), .C2(new_n407), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n406), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n355), .A2(new_n240), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n316), .A2(new_n239), .A3(new_n328), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G227gat), .A2(G233gat), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT70), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT34), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(KEYINPUT70), .B(KEYINPUT34), .C1(new_n417), .C2(new_n419), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XOR2_X1   g223(.A(G15gat), .B(G43gat), .Z(new_n425));
  XNOR2_X1  g224(.A(G71gat), .B(G99gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n418), .B1(new_n415), .B2(new_n416), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(KEYINPUT33), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT32), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AOI221_X4 g231(.A(new_n430), .B1(KEYINPUT33), .B2(new_n427), .C1(new_n417), .C2(new_n419), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n424), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n355), .A2(new_n240), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n239), .B1(new_n316), .B2(new_n328), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n419), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT32), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n440), .A3(new_n427), .ZN(new_n441));
  INV_X1    g240(.A(new_n427), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n437), .B(KEYINPUT32), .C1(new_n439), .C2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n441), .A2(new_n423), .A3(new_n422), .A4(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n414), .A2(new_n434), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT35), .B1(new_n375), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT91), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT91), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n448), .B(KEYINPUT35), .C1(new_n375), .C2(new_n445), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT71), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n444), .A3(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n424), .B(KEYINPUT71), .C1(new_n432), .C2(new_n433), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n349), .B(new_n368), .C1(new_n361), .C2(new_n346), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT30), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n372), .A2(new_n371), .A3(new_n368), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(new_n370), .A3(new_n414), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT88), .B1(new_n280), .B2(new_n273), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT6), .B1(new_n280), .B2(new_n273), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n269), .A2(new_n463), .A3(new_n274), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n465), .A2(new_n275), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n466), .A2(KEYINPUT35), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n447), .A2(new_n449), .B1(new_n460), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT36), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n469), .A3(new_n452), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n434), .A2(new_n444), .A3(KEYINPUT36), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n406), .A2(new_n413), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n375), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT38), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n330), .B1(new_n347), .B2(new_n348), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT37), .B1(new_n477), .B2(new_n346), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n385), .B1(new_n358), .B2(new_n360), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT37), .ZN(new_n481));
  OR3_X1    g280(.A1(new_n480), .A2(new_n481), .A3(new_n368), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n466), .A2(new_n482), .A3(KEYINPUT90), .A4(new_n455), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n362), .A2(KEYINPUT37), .A3(new_n365), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n481), .A2(new_n368), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT38), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT90), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n465), .A2(new_n275), .A3(new_n455), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n480), .A2(new_n481), .A3(new_n368), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n483), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n244), .B1(new_n267), .B2(new_n241), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT39), .B1(new_n257), .B2(new_n243), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT39), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n494), .A2(new_n273), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n461), .B(new_n464), .C1(new_n497), .C2(KEYINPUT40), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n494), .A2(KEYINPUT40), .A3(new_n273), .A4(new_n496), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT89), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n499), .A2(KEYINPUT89), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n458), .A2(new_n370), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n473), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n475), .B1(new_n491), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n468), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(G197gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT11), .B(G169gat), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n508), .B(new_n509), .Z(new_n510));
  XOR2_X1   g309(.A(new_n510), .B(KEYINPUT12), .Z(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G229gat), .A2(G233gat), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(KEYINPUT13), .Z(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G8gat), .ZN(new_n516));
  INV_X1    g315(.A(G22gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(G15gat), .ZN(new_n518));
  INV_X1    g317(.A(G15gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(G22gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT16), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n518), .B(new_n520), .C1(new_n521), .C2(G1gat), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n516), .B1(new_n522), .B2(KEYINPUT94), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n522), .B1(G1gat), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  OAI221_X1 g325(.A(new_n522), .B1(KEYINPUT94), .B2(new_n516), .C1(G1gat), .C2(new_n524), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT96), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(KEYINPUT96), .A3(new_n527), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G50gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G43gat), .ZN(new_n534));
  INV_X1    g333(.A(G43gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(G50gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(new_n536), .A3(KEYINPUT15), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT15), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(KEYINPUT92), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT92), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(G43gat), .ZN(new_n542));
  AOI21_X1  g341(.A(G50gat), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT93), .B1(new_n533), .B2(G43gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT93), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n545), .A2(new_n535), .A3(G50gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n539), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT14), .B(G29gat), .ZN(new_n549));
  INV_X1    g348(.A(G36gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G29gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n538), .B1(new_n548), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n537), .B1(new_n551), .B2(new_n553), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n532), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n530), .A2(new_n557), .A3(new_n531), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n515), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n548), .A2(new_n554), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n537), .ZN(new_n563));
  INV_X1    g362(.A(new_n556), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n563), .A2(KEYINPUT95), .A3(KEYINPUT17), .A4(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(KEYINPUT95), .A2(KEYINPUT17), .ZN(new_n566));
  NAND2_X1  g365(.A1(KEYINPUT95), .A2(KEYINPUT17), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n566), .B(new_n567), .C1(new_n555), .C2(new_n556), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n528), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(new_n513), .A3(new_n560), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT18), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n561), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n571), .A2(KEYINPUT18), .A3(new_n513), .A4(new_n560), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n512), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n573), .ZN(new_n578));
  INV_X1    g377(.A(new_n561), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n578), .A2(new_n512), .A3(new_n575), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n506), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n282), .ZN(new_n584));
  AND2_X1   g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G57gat), .B(G64gat), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(G57gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(G64gat), .ZN(new_n592));
  INV_X1    g391(.A(G64gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(G57gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G71gat), .B(G78gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n589), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT97), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n603), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n532), .B1(new_n600), .B2(new_n599), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n612), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n617));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n620));
  NAND2_X1  g419(.A1(G99gat), .A2(G106gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT8), .ZN(new_n622));
  NAND2_X1  g421(.A1(G85gat), .A2(G92gat), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT7), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(G85gat), .ZN(new_n626));
  INV_X1    g425(.A(G92gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n622), .A2(new_n625), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G99gat), .B(G106gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g432(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI22_X1  g435(.A1(KEYINPUT8), .A2(new_n621), .B1(new_n626), .B2(new_n627), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n631), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n620), .B1(new_n558), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(new_n569), .B2(new_n640), .ZN(new_n642));
  XOR2_X1   g441(.A(G190gat), .B(G218gat), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n644), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n619), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n647), .ZN(new_n649));
  INV_X1    g448(.A(new_n619), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n649), .A2(new_n645), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n615), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n599), .B1(new_n633), .B2(new_n638), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n630), .A2(new_n632), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n636), .A2(new_n631), .A3(new_n637), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n657), .A2(new_n590), .A3(new_n658), .A4(new_n598), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n655), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n639), .A2(KEYINPUT98), .A3(new_n590), .A4(new_n598), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT10), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT10), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n654), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n654), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n660), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n665), .A2(new_n667), .A3(new_n671), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n653), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n583), .A2(new_n584), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G1gat), .ZN(G1324gat));
  INV_X1    g479(.A(new_n503), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n677), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n583), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(G8gat), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT16), .B(G8gat), .Z(new_n686));
  NAND3_X1  g485(.A1(new_n583), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n688), .A3(new_n685), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n687), .B2(new_n685), .ZN(new_n691));
  OAI221_X1 g490(.A(new_n684), .B1(new_n685), .B2(new_n687), .C1(new_n690), .C2(new_n691), .ZN(G1325gat));
  NAND2_X1  g491(.A1(new_n583), .A2(new_n678), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n472), .A2(KEYINPUT100), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT100), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n470), .A2(new_n695), .A3(new_n471), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G15gat), .B1(new_n693), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n453), .A2(new_n519), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n693), .B2(new_n699), .ZN(G1326gat));
  NOR2_X1   g499(.A1(new_n693), .A2(new_n414), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT43), .B(G22gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  INV_X1    g502(.A(new_n615), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n704), .A2(new_n582), .A3(new_n675), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n652), .B(new_n705), .C1(new_n468), .C2(new_n505), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n706), .A2(G29gat), .A3(new_n282), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT45), .Z(new_n708));
  OAI211_X1 g507(.A(KEYINPUT44), .B(new_n652), .C1(new_n468), .C2(new_n505), .ZN(new_n709));
  INV_X1    g508(.A(new_n652), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n490), .A2(new_n486), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n488), .A2(new_n489), .A3(new_n487), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n504), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n375), .A2(new_n714), .A3(new_n473), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n375), .B2(new_n473), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n713), .A2(new_n697), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n460), .A2(new_n467), .ZN(new_n719));
  INV_X1    g518(.A(new_n445), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n720), .A2(new_n282), .A3(new_n370), .A4(new_n458), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n448), .B1(new_n721), .B2(KEYINPUT35), .ZN(new_n722));
  INV_X1    g521(.A(new_n449), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n719), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n710), .B1(new_n718), .B2(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n705), .B(new_n709), .C1(new_n725), .C2(KEYINPUT44), .ZN(new_n726));
  OAI21_X1  g525(.A(G29gat), .B1(new_n726), .B2(new_n282), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n708), .A2(new_n727), .ZN(G1328gat));
  NAND2_X1  g527(.A1(new_n503), .A2(new_n550), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n706), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT46), .ZN(new_n731));
  OAI21_X1  g530(.A(G36gat), .B1(new_n726), .B2(new_n681), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n731), .A2(KEYINPUT102), .A3(new_n732), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(G1329gat));
  INV_X1    g536(.A(new_n726), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n540), .A2(new_n542), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n694), .A2(new_n696), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  OR2_X1    g541(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n706), .A2(new_n454), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n744), .A2(new_n739), .B1(KEYINPUT103), .B2(KEYINPUT47), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n743), .B1(new_n742), .B2(new_n745), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(G1330gat));
  OAI21_X1  g548(.A(G50gat), .B1(new_n726), .B2(new_n414), .ZN(new_n750));
  OR3_X1    g549(.A1(new_n706), .A2(G50gat), .A3(new_n414), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT48), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1331gat));
  NAND2_X1  g553(.A1(new_n718), .A2(new_n724), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n615), .A2(new_n652), .A3(new_n581), .A4(new_n676), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n282), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(new_n591), .ZN(G1332gat));
  NOR2_X1   g558(.A1(new_n757), .A2(new_n681), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  AND2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n760), .B2(new_n761), .ZN(G1333gat));
  OR3_X1    g563(.A1(new_n757), .A2(G71gat), .A3(new_n454), .ZN(new_n765));
  OAI21_X1  g564(.A(G71gat), .B1(new_n757), .B2(new_n697), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g567(.A1(new_n757), .A2(new_n414), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g569(.A1(new_n704), .A2(new_n581), .A3(new_n676), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n709), .B(new_n771), .C1(new_n725), .C2(KEYINPUT44), .ZN(new_n772));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772), .B2(new_n282), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n584), .A2(new_n626), .A3(new_n675), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n704), .A2(new_n581), .ZN(new_n776));
  AND4_X1   g575(.A1(KEYINPUT51), .A2(new_n755), .A3(new_n652), .A4(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT51), .B1(new_n725), .B2(new_n776), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT104), .ZN(G1336gat));
  NOR2_X1   g580(.A1(KEYINPUT106), .A2(KEYINPUT52), .ZN(new_n782));
  AND2_X1   g581(.A1(KEYINPUT106), .A2(KEYINPUT52), .ZN(new_n783));
  OAI21_X1  g582(.A(G92gat), .B1(new_n772), .B2(new_n681), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n503), .A2(new_n627), .A3(new_n675), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n785), .B(KEYINPUT105), .Z(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n777), .B2(new_n778), .ZN(new_n787));
  AOI211_X1 g586(.A(new_n782), .B(new_n783), .C1(new_n784), .C2(new_n787), .ZN(new_n788));
  AND4_X1   g587(.A1(KEYINPUT106), .A2(new_n784), .A3(new_n787), .A4(KEYINPUT52), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(G1337gat));
  XOR2_X1   g589(.A(KEYINPUT108), .B(G99gat), .Z(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n454), .A2(new_n676), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n777), .B2(new_n778), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n772), .A2(new_n697), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT107), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n792), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n795), .A2(new_n796), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n794), .B1(new_n798), .B2(new_n799), .ZN(G1338gat));
  OAI21_X1  g599(.A(G106gat), .B1(new_n772), .B2(new_n414), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n414), .A2(G106gat), .A3(new_n676), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n777), .B2(new_n778), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g604(.A1(new_n677), .A2(new_n581), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n660), .A2(new_n661), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n663), .ZN(new_n808));
  INV_X1    g607(.A(new_n664), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n666), .A3(new_n809), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n810), .A2(KEYINPUT54), .A3(new_n665), .ZN(new_n811));
  XNOR2_X1  g610(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n654), .B(new_n812), .C1(new_n662), .C2(new_n664), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n672), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT110), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n813), .A2(KEYINPUT110), .A3(new_n672), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n811), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT111), .B1(new_n818), .B2(KEYINPUT55), .ZN(new_n819));
  INV_X1    g618(.A(new_n674), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n818), .B2(KEYINPUT55), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n810), .A2(KEYINPUT54), .A3(new_n665), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n813), .A2(KEYINPUT110), .A3(new_n672), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT110), .B1(new_n813), .B2(new_n672), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT111), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n819), .A2(new_n821), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT112), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n513), .B1(new_n571), .B2(new_n560), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n559), .A2(new_n560), .A3(new_n515), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n510), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT113), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n835), .B(new_n510), .C1(new_n831), .C2(new_n832), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n652), .A2(new_n837), .A3(new_n580), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n819), .A2(new_n821), .A3(new_n839), .A4(new_n828), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n830), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT114), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n830), .A2(new_n838), .A3(new_n843), .A4(new_n840), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n581), .A3(new_n840), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n834), .A2(new_n580), .A3(new_n675), .A4(new_n836), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n710), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n806), .B1(new_n850), .B2(new_n615), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n282), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n460), .ZN(new_n853));
  INV_X1    g652(.A(G113gat), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n853), .A2(new_n854), .A3(new_n582), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n503), .A2(new_n445), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n581), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n855), .B1(new_n854), .B2(new_n859), .ZN(G1340gat));
  INV_X1    g659(.A(G120gat), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n853), .A2(new_n861), .A3(new_n676), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n858), .A2(new_n675), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n861), .B2(new_n863), .ZN(G1341gat));
  OAI21_X1  g663(.A(G127gat), .B1(new_n853), .B2(new_n615), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n615), .A2(G127gat), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n857), .B2(new_n866), .ZN(G1342gat));
  OAI21_X1  g666(.A(G134gat), .B1(new_n853), .B2(new_n710), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n710), .A2(G134gat), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT56), .B1(new_n857), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT56), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n852), .A2(new_n872), .A3(new_n856), .A4(new_n869), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n868), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n868), .A2(new_n871), .A3(KEYINPUT115), .A4(new_n873), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1343gat));
  XNOR2_X1  g677(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n697), .A2(new_n584), .A3(new_n681), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n473), .A2(KEYINPUT57), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n847), .B(KEYINPUT116), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n825), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g684(.A(KEYINPUT117), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n827), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n581), .A3(new_n821), .ZN(new_n888));
  AOI211_X1 g687(.A(KEYINPUT118), .B(new_n652), .C1(new_n883), .C2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n837), .A2(KEYINPUT116), .A3(new_n580), .A4(new_n675), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n847), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n885), .A2(new_n827), .A3(new_n886), .ZN(new_n894));
  OAI211_X1 g693(.A(KEYINPUT55), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n895));
  INV_X1    g694(.A(new_n580), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n674), .B(new_n895), .C1(new_n896), .C2(new_n576), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n891), .B(new_n893), .C1(new_n894), .C2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n890), .B1(new_n898), .B2(new_n710), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n889), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n704), .B1(new_n900), .B2(new_n845), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n806), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n842), .A2(new_n844), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n898), .A2(new_n710), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT118), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n898), .A2(new_n890), .A3(new_n710), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n615), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT119), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n882), .B1(new_n903), .B2(new_n910), .ZN(new_n911));
  AOI22_X1  g710(.A1(new_n710), .A2(new_n848), .B1(new_n842), .B2(new_n844), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n912), .A2(new_n704), .B1(new_n581), .B2(new_n677), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT57), .B1(new_n913), .B2(new_n473), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n581), .B(new_n881), .C1(new_n911), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(G141gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(new_n473), .A3(new_n881), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n582), .A2(G141gat), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT120), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n879), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n879), .ZN(new_n923));
  AOI211_X1 g722(.A(new_n920), .B(new_n923), .C1(new_n915), .C2(G141gat), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n922), .A2(new_n924), .ZN(G1344gat));
  INV_X1    g724(.A(new_n917), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n204), .A3(new_n675), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT59), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G148gat), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n911), .A2(new_n914), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n930), .A2(new_n880), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n929), .B1(new_n931), .B2(new_n675), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n913), .A2(KEYINPUT57), .A3(new_n473), .ZN(new_n933));
  INV_X1    g732(.A(new_n829), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n838), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n704), .B1(new_n905), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n473), .B1(new_n936), .B2(new_n806), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT57), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n676), .B1(new_n933), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n881), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n928), .B1(new_n941), .B2(G148gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n927), .B1(new_n932), .B2(new_n942), .ZN(G1345gat));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n212), .A3(new_n704), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n930), .A2(new_n615), .A3(new_n880), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n212), .ZN(G1346gat));
  NAND3_X1  g745(.A1(new_n926), .A2(new_n213), .A3(new_n652), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n652), .B(new_n881), .C1(new_n911), .C2(new_n914), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G162gat), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n948), .A2(new_n949), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(G1347gat));
  NAND3_X1  g752(.A1(new_n503), .A2(new_n282), .A3(new_n414), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n851), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(new_n453), .ZN(new_n956));
  OAI21_X1  g755(.A(G169gat), .B1(new_n956), .B2(new_n582), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n503), .A2(new_n720), .ZN(new_n958));
  XOR2_X1   g757(.A(new_n958), .B(KEYINPUT123), .Z(new_n959));
  NAND3_X1  g758(.A1(new_n913), .A2(new_n282), .A3(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n292), .A3(new_n581), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n957), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT124), .ZN(G1348gat));
  AOI21_X1  g763(.A(G176gat), .B1(new_n961), .B2(new_n675), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n454), .A2(new_n293), .A3(new_n676), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n955), .B2(new_n966), .ZN(G1349gat));
  OAI21_X1  g766(.A(G183gat), .B1(new_n956), .B2(new_n615), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n961), .A2(new_n318), .A3(new_n704), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g770(.A1(new_n961), .A2(new_n317), .A3(new_n652), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n453), .A3(new_n652), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n973), .A2(new_n974), .A3(G190gat), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n974), .B1(new_n973), .B2(G190gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(G1351gat));
  NOR3_X1   g776(.A1(new_n741), .A2(new_n681), .A3(new_n414), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n913), .A2(new_n978), .A3(new_n282), .ZN(new_n979));
  XOR2_X1   g778(.A(new_n979), .B(KEYINPUT125), .Z(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(new_n581), .ZN(new_n981));
  INV_X1    g780(.A(G197gat), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n933), .A2(new_n939), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n697), .A2(new_n282), .A3(new_n503), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n984), .B(KEYINPUT126), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n582), .A2(new_n982), .ZN(new_n987));
  AOI22_X1  g786(.A1(new_n981), .A2(new_n982), .B1(new_n986), .B2(new_n987), .ZN(G1352gat));
  INV_X1    g787(.A(G204gat), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n989), .B1(new_n940), .B2(new_n985), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n676), .A2(G204gat), .ZN(new_n991));
  NAND4_X1  g790(.A1(new_n913), .A2(new_n978), .A3(new_n282), .A4(new_n991), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT62), .ZN(new_n993));
  OR3_X1    g792(.A1(new_n990), .A2(new_n993), .A3(KEYINPUT127), .ZN(new_n994));
  OAI21_X1  g793(.A(KEYINPUT127), .B1(new_n990), .B2(new_n993), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(G1353gat));
  OR2_X1    g795(.A1(new_n984), .A2(new_n615), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n332), .B1(new_n983), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT63), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n980), .A2(new_n332), .A3(new_n704), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1354gat));
  NAND2_X1  g801(.A1(new_n980), .A2(new_n652), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n710), .A2(new_n333), .ZN(new_n1004));
  AOI22_X1  g803(.A1(new_n1003), .A2(new_n333), .B1(new_n986), .B2(new_n1004), .ZN(G1355gat));
endmodule


