//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n571, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1224, new_n1225, new_n1226;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G219), .A3(G218), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT67), .B(G2105), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(G137), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n460), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT69), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(new_n470), .A3(new_n467), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT67), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT68), .Z(new_n478));
  NAND2_X1  g053(.A1(new_n463), .A2(G125), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n469), .A2(new_n471), .B1(new_n476), .B2(new_n480), .ZN(G160));
  AND2_X1   g056(.A1(new_n461), .A2(new_n462), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n464), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT70), .Z(new_n485));
  AOI21_X1  g060(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n464), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n485), .A2(new_n490), .ZN(G162));
  NAND3_X1  g066(.A1(new_n463), .A2(new_n464), .A3(G138), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n463), .A2(new_n464), .A3(G138), .A4(new_n496), .ZN(new_n497));
  AND2_X1   g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  OR2_X1    g073(.A1(new_n472), .A2(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n463), .A2(new_n498), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n494), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  OR2_X1    g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n507), .A2(new_n511), .A3(G88), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(G50), .A3(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT72), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n510), .B1(new_n516), .B2(new_n517), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n511), .A2(G51), .A3(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  OAI21_X1  g102(.A(G89), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n522), .A2(new_n530), .ZN(G168));
  NAND3_X1  g106(.A1(new_n507), .A2(new_n511), .A3(G90), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n511), .A2(G52), .A3(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(G64), .B1(new_n523), .B2(new_n524), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n509), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  AOI22_X1  g113(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n509), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n511), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n524), .A2(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n541), .A2(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT73), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  INV_X1    g127(.A(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(KEYINPUT6), .A2(G651), .ZN(new_n554));
  NAND2_X1  g129(.A1(KEYINPUT6), .A2(G651), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n556), .B(G53), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n511), .A2(G53), .A3(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n557), .A2(new_n558), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n525), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n505), .A2(new_n506), .B1(new_n554), .B2(new_n555), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n566), .A2(G651), .B1(new_n567), .B2(G91), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n563), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  AND2_X1   g145(.A1(new_n528), .A2(new_n529), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n521), .B(new_n520), .C1(new_n571), .C2(new_n525), .ZN(G286));
  INV_X1    g147(.A(new_n517), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT72), .B1(new_n512), .B2(new_n513), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n573), .A2(new_n574), .B1(new_n509), .B2(new_n508), .ZN(G303));
  INV_X1    g150(.A(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n505), .A2(new_n576), .A3(new_n506), .ZN(new_n577));
  AOI22_X1  g152(.A1(G49), .A2(new_n556), .B1(new_n577), .B2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n567), .A2(G87), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT75), .ZN(G288));
  NAND3_X1  g156(.A1(new_n511), .A2(G48), .A3(G543), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n556), .A2(KEYINPUT76), .A3(G48), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n525), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n567), .B2(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(G305));
  INV_X1    g166(.A(G47), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n541), .A2(new_n592), .B1(new_n543), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n507), .A2(G60), .ZN(new_n596));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n509), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n567), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n543), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n525), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(G54), .B2(new_n556), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n601), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n601), .B1(new_n612), .B2(G868), .ZN(G321));
  MUX2_X1   g189(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g190(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n612), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n612), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g197(.A1(new_n483), .A2(G123), .B1(G135), .B2(new_n486), .ZN(new_n623));
  OAI221_X1 g198(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n464), .C2(G111), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT79), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n463), .A2(new_n466), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT77), .B(G2100), .Z(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT78), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n631), .B(new_n634), .Z(new_n635));
  OAI211_X1 g210(.A(new_n628), .B(new_n635), .C1(KEYINPUT78), .C2(new_n633), .ZN(G156));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT14), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n646), .A2(new_n649), .ZN(new_n651));
  AND3_X1   g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n656), .B2(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT81), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2100), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n654), .A2(new_n655), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(G2096), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n659), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n671), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(KEYINPUT82), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n686), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n668), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(new_n667), .A3(new_n687), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G23), .ZN(new_n696));
  INV_X1    g271(.A(new_n580), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT33), .ZN(new_n699));
  INV_X1    g274(.A(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n695), .A2(G22), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n695), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1971), .ZN(new_n704));
  NOR2_X1   g279(.A1(G6), .A2(G16), .ZN(new_n705));
  INV_X1    g280(.A(G305), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G16), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT32), .B(G1981), .Z(new_n708));
  XOR2_X1   g283(.A(new_n707), .B(new_n708), .Z(new_n709));
  NOR3_X1   g284(.A1(new_n701), .A2(new_n704), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n486), .A2(G131), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT83), .ZN(new_n714));
  OAI21_X1  g289(.A(KEYINPUT84), .B1(G95), .B2(G2105), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NOR3_X1   g291(.A1(KEYINPUT84), .A2(G95), .A3(G2105), .ZN(new_n717));
  OAI221_X1 g292(.A(G2104), .B1(new_n716), .B2(new_n717), .C1(new_n464), .C2(G107), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n483), .A2(G119), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n714), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT85), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G25), .B2(new_n722), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT35), .B(G1991), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT86), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n724), .A2(new_n727), .ZN(new_n729));
  MUX2_X1   g304(.A(G24), .B(G290), .S(G16), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1986), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n710), .A2(new_n711), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n712), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n734), .B(new_n735), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n722), .A2(G35), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n722), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT29), .Z(new_n739));
  INV_X1    g314(.A(G2090), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n739), .B1(KEYINPUT99), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n740), .A2(KEYINPUT99), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n722), .A2(G33), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n486), .A2(G139), .ZN(new_n746));
  AND2_X1   g321(.A1(G103), .A2(G2104), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n473), .A2(new_n475), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT90), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n473), .A2(new_n475), .A3(new_n747), .A4(KEYINPUT90), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n752));
  AND3_X1   g327(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(new_n750), .B2(new_n751), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n746), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT91), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n752), .ZN(new_n758));
  AOI21_X1  g333(.A(KEYINPUT90), .B1(new_n464), .B2(new_n747), .ZN(new_n759));
  INV_X1    g334(.A(new_n751), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n763), .A2(KEYINPUT91), .A3(new_n746), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n757), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(G115), .A2(G2104), .ZN(new_n766));
  INV_X1    g341(.A(G127), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n482), .B2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT92), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI211_X1 g345(.A(KEYINPUT92), .B(new_n766), .C1(new_n482), .C2(new_n767), .ZN(new_n771));
  AND3_X1   g346(.A1(new_n770), .A2(new_n476), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n745), .B1(new_n765), .B2(new_n773), .ZN(new_n774));
  AOI211_X1 g349(.A(KEYINPUT93), .B(new_n772), .C1(new_n757), .C2(new_n764), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n744), .B1(new_n776), .B2(new_n722), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(G2072), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(G2072), .ZN(new_n779));
  NOR2_X1   g354(.A1(G16), .A2(G19), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n546), .B2(G16), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n781), .A2(G1341), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n625), .B(KEYINPUT79), .ZN(new_n783));
  OAI22_X1  g358(.A1(new_n783), .A2(new_n722), .B1(G1341), .B2(new_n781), .ZN(new_n784));
  INV_X1    g359(.A(G1961), .ZN(new_n785));
  NOR2_X1   g360(.A1(G171), .A2(new_n695), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G5), .B2(new_n695), .ZN(new_n787));
  AOI211_X1 g362(.A(new_n782), .B(new_n784), .C1(new_n785), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n695), .A2(G20), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT23), .Z(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G299), .B2(G16), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G1956), .Z(new_n792));
  INV_X1    g367(.A(G2084), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT24), .B(G34), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(new_n722), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT94), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n480), .A2(new_n476), .ZN(new_n797));
  INV_X1    g372(.A(new_n471), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n470), .B1(new_n465), .B2(new_n467), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n796), .B1(new_n800), .B2(new_n722), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n792), .B1(new_n793), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT31), .B(G11), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT98), .B(G28), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n804), .A2(KEYINPUT30), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(KEYINPUT30), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(new_n722), .ZN(new_n807));
  OAI221_X1 g382(.A(new_n803), .B1(new_n805), .B2(new_n807), .C1(new_n787), .C2(new_n785), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n612), .A2(new_n695), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G4), .B2(new_n695), .ZN(new_n810));
  INV_X1    g385(.A(G1348), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n788), .A2(new_n802), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n722), .A2(G32), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n486), .A2(G141), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n466), .A2(new_n816), .A3(G105), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(KEYINPUT95), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n476), .A2(new_n463), .A3(G129), .ZN(new_n822));
  NAND3_X1  g397(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT26), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT96), .B1(new_n821), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AOI22_X1  g403(.A1(G141), .A2(new_n486), .B1(new_n817), .B2(new_n819), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT96), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n829), .A2(new_n830), .A3(new_n822), .A4(new_n825), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n814), .B1(new_n833), .B2(new_n722), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT27), .B(G1996), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n722), .A2(G26), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT28), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n486), .A2(G140), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n464), .A2(G116), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n483), .A2(KEYINPUT88), .A3(G128), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n476), .A2(new_n463), .A3(G128), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT88), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n842), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n838), .B1(new_n847), .B2(new_n722), .ZN(new_n848));
  INV_X1    g423(.A(G2067), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n836), .B(new_n850), .C1(new_n793), .C2(new_n801), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n722), .A2(G27), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(G164), .B2(new_n722), .ZN(new_n853));
  INV_X1    g428(.A(G2078), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n695), .A2(G21), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(G168), .B2(new_n695), .ZN(new_n857));
  XOR2_X1   g432(.A(KEYINPUT97), .B(G1966), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n855), .B(new_n859), .C1(new_n810), .C2(new_n811), .ZN(new_n860));
  OR3_X1    g435(.A1(new_n813), .A2(new_n851), .A3(new_n860), .ZN(new_n861));
  NOR4_X1   g436(.A1(new_n743), .A2(new_n778), .A3(new_n779), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n736), .A2(new_n862), .ZN(G150));
  INV_X1    g438(.A(G150), .ZN(G311));
  NAND2_X1  g439(.A1(new_n612), .A2(G559), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT38), .ZN(new_n866));
  INV_X1    g441(.A(G55), .ZN(new_n867));
  XNOR2_X1  g442(.A(KEYINPUT100), .B(G93), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n541), .A2(new_n867), .B1(new_n543), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n507), .A2(G67), .ZN(new_n870));
  NAND2_X1  g445(.A1(G80), .A2(G543), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n509), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n546), .A2(new_n873), .ZN(new_n874));
  OAI22_X1  g449(.A1(new_n540), .A2(new_n545), .B1(new_n869), .B2(new_n872), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n866), .B(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n879));
  INV_X1    g454(.A(G860), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n873), .A2(new_n880), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT37), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(G145));
  NAND2_X1  g460(.A1(new_n783), .A2(G160), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n627), .A2(new_n800), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n886), .A2(new_n887), .A3(G162), .ZN(new_n888));
  AOI21_X1  g463(.A(G162), .B1(new_n886), .B2(new_n887), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT103), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n627), .A2(new_n800), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n783), .A2(G160), .ZN(new_n893));
  OAI22_X1  g468(.A1(new_n892), .A2(new_n893), .B1(new_n485), .B2(new_n490), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n886), .A2(new_n887), .A3(G162), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT101), .B1(new_n774), .B2(new_n775), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT91), .B1(new_n763), .B2(new_n746), .ZN(new_n899));
  INV_X1    g474(.A(new_n746), .ZN(new_n900));
  AOI211_X1 g475(.A(new_n756), .B(new_n900), .C1(new_n761), .C2(new_n762), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n773), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT93), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n765), .A2(new_n745), .A3(new_n773), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n847), .A2(new_n827), .A3(new_n831), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n843), .A2(new_n846), .ZN(new_n908));
  INV_X1    g483(.A(new_n842), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n827), .A2(new_n831), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n907), .A2(new_n910), .A3(new_n503), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n909), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(new_n828), .B2(new_n832), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n847), .A2(new_n827), .A3(new_n831), .ZN(new_n914));
  AOI21_X1  g489(.A(G164), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n898), .A2(new_n906), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n720), .B(new_n630), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n483), .A2(G130), .ZN(new_n919));
  OAI221_X1 g494(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n464), .C2(G118), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n486), .A2(G142), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n918), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n503), .B1(new_n907), .B2(new_n910), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n913), .A2(G164), .A3(new_n914), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n776), .A2(new_n905), .A3(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n917), .A2(new_n924), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n924), .B1(new_n917), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n897), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT104), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n897), .B(new_n933), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n917), .A2(new_n928), .ZN(new_n936));
  INV_X1    g511(.A(new_n924), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n917), .A2(new_n924), .A3(new_n928), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n888), .A2(new_n889), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n938), .A2(KEYINPUT102), .A3(new_n939), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G37), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n935), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g523(.A(new_n876), .B(new_n619), .Z(new_n949));
  NAND2_X1  g524(.A1(new_n611), .A2(G299), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n606), .A2(new_n563), .A3(new_n568), .A4(new_n610), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n950), .A2(KEYINPUT105), .A3(new_n951), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n949), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT41), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n950), .A2(new_n958), .A3(new_n951), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n952), .A2(KEYINPUT41), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n962), .A2(new_n960), .A3(new_n959), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n949), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n957), .A2(new_n964), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n965), .A2(KEYINPUT109), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n967));
  NAND2_X1  g542(.A1(G290), .A2(new_n580), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n697), .A2(new_n599), .A3(new_n595), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(G166), .A2(KEYINPUT107), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n972));
  AOI211_X1 g547(.A(new_n972), .B(new_n510), .C1(new_n516), .C2(new_n517), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n706), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(G303), .A2(new_n972), .ZN(new_n975));
  NAND2_X1  g550(.A1(G166), .A2(KEYINPUT107), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(new_n976), .A3(G305), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n970), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n971), .A2(new_n973), .A3(new_n706), .ZN(new_n979));
  AOI21_X1  g554(.A(G305), .B1(new_n975), .B2(new_n976), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n968), .A2(new_n969), .A3(new_n967), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n595), .A2(new_n599), .B1(new_n579), .B2(new_n578), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n580), .A2(new_n598), .A3(new_n594), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT108), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n978), .B1(new_n981), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT42), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n966), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n965), .A2(KEYINPUT109), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n988), .B1(new_n966), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(G868), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(G868), .B2(new_n873), .ZN(G295));
  OAI21_X1  g568(.A(new_n992), .B1(G868), .B2(new_n873), .ZN(G331));
  OAI21_X1  g569(.A(KEYINPUT110), .B1(new_n534), .B2(new_n537), .ZN(new_n995));
  INV_X1    g570(.A(G64), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n505), .B2(new_n506), .ZN(new_n997));
  INV_X1    g572(.A(new_n536), .ZN(new_n998));
  OAI21_X1  g573(.A(G651), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n999), .A2(new_n1000), .A3(new_n533), .A4(new_n532), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(G286), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(G171), .A2(G168), .A3(new_n1000), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n876), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n874), .A2(new_n1002), .A3(new_n1003), .A4(new_n875), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n877), .A2(KEYINPUT111), .A3(new_n1003), .A4(new_n1002), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n952), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n985), .B1(new_n979), .B2(new_n980), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n986), .A2(new_n977), .A3(new_n974), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n963), .A2(new_n961), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1012), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1018), .A2(new_n946), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n962), .A2(new_n959), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1008), .A2(new_n1020), .A3(new_n1009), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n954), .A2(new_n1005), .A3(new_n955), .A4(new_n1007), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n987), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1019), .A2(KEYINPUT43), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1017), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n952), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n987), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT43), .B1(new_n1019), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT44), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT43), .ZN(new_n1031));
  AND4_X1   g606(.A1(new_n1031), .A2(new_n1024), .A3(new_n1018), .A4(new_n946), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n946), .A3(new_n1018), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT43), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1034), .B2(KEYINPUT112), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT112), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n1036), .A3(KEYINPUT43), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1030), .B1(new_n1038), .B2(KEYINPUT44), .ZN(G397));
  OAI211_X1 g614(.A(new_n797), .B(G40), .C1(new_n798), .C2(new_n799), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G1384), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT45), .B1(new_n503), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1044), .A2(G1996), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1045), .B(KEYINPUT46), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1044), .B(KEYINPUT113), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n828), .B2(new_n832), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n912), .A2(G2067), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n847), .A2(new_n849), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT114), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n1047), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1046), .A2(new_n1048), .A3(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT47), .ZN(new_n1055));
  XOR2_X1   g630(.A(new_n1053), .B(KEYINPUT115), .Z(new_n1056));
  NOR2_X1   g631(.A1(new_n833), .A2(G1996), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1057), .B1(new_n1048), .B2(new_n1045), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n720), .B(new_n726), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1047), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1044), .A2(G1986), .A3(G290), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT48), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1055), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n721), .A2(new_n727), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(KEYINPUT125), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1050), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1065), .B1(new_n1047), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G8), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n503), .A2(new_n1042), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT45), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1971), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1040), .B1(KEYINPUT50), .B2(new_n1073), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n503), .A2(new_n1080), .A3(new_n1042), .ZN(new_n1081));
  XOR2_X1   g656(.A(KEYINPUT116), .B(G2090), .Z(new_n1082));
  NAND3_X1  g657(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1071), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G166), .A2(new_n1071), .ZN(new_n1085));
  XOR2_X1   g660(.A(new_n1085), .B(KEYINPUT55), .Z(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1076), .A2(new_n858), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1079), .A2(new_n793), .A3(new_n1081), .ZN(new_n1090));
  AOI211_X1 g665(.A(new_n1071), .B(G286), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1071), .B1(new_n1041), .B2(new_n1074), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(G288), .B2(new_n700), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n697), .A2(G1976), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT49), .ZN(new_n1096));
  INV_X1    g671(.A(G1981), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n586), .A2(new_n590), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1097), .B1(new_n586), .B2(new_n590), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1074), .A2(G40), .A3(G160), .ZN(new_n1102));
  NAND2_X1  g677(.A1(G305), .A2(G1981), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(KEYINPUT49), .A3(new_n1098), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .A4(G8), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1094), .B(G8), .C1(new_n1040), .C2(new_n1073), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT52), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1095), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1971), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1073), .A2(KEYINPUT50), .ZN(new_n1111));
  AND4_X1   g686(.A1(new_n1041), .A2(new_n1081), .A3(new_n1111), .A4(new_n1082), .ZN(new_n1112));
  OAI21_X1  g687(.A(G8), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n1086), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1088), .A2(new_n1091), .A3(new_n1109), .A4(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1108), .B1(new_n1086), .B2(new_n1113), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1118), .A2(KEYINPUT63), .A3(new_n1088), .A4(new_n1091), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(G288), .A2(G1976), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1099), .B1(new_n1105), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1092), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI211_X1 g699(.A(KEYINPUT117), .B(new_n1099), .C1(new_n1105), .C2(new_n1121), .ZN(new_n1125));
  OAI22_X1  g700(.A1(new_n1124), .A2(new_n1125), .B1(new_n1088), .B2(new_n1108), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT118), .B1(new_n1120), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n1129), .B(new_n1126), .C1(new_n1117), .C2(new_n1119), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1072), .A2(new_n1075), .A3(new_n854), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT53), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1079), .A2(KEYINPUT122), .A3(new_n1081), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1041), .A2(new_n1081), .A3(new_n1111), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1135), .A2(new_n1138), .A3(new_n785), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1134), .A2(G301), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(G301), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1132), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(G171), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1145), .A2(new_n1140), .A3(KEYINPUT54), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1089), .A2(G168), .A3(new_n1090), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(G8), .ZN(new_n1148));
  AOI21_X1  g723(.A(G168), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT51), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1147), .A2(new_n1151), .A3(G8), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1118), .A2(new_n1088), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1143), .A2(new_n1146), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1135), .A2(new_n1138), .A3(new_n811), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1074), .A2(new_n1157), .A3(G160), .A4(G40), .ZN(new_n1158));
  OAI21_X1  g733(.A(KEYINPUT121), .B1(new_n1040), .B2(new_n1073), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n849), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1156), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT124), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1156), .A2(new_n1165), .A3(KEYINPUT60), .A4(new_n1161), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n612), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT57), .ZN(new_n1173));
  OAI21_X1  g748(.A(G299), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1174), .B(new_n1175), .Z(new_n1176));
  XOR2_X1   g751(.A(KEYINPUT119), .B(G1956), .Z(new_n1177));
  AOI21_X1  g752(.A(new_n1177), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1178));
  XNOR2_X1  g753(.A(KEYINPUT56), .B(G2072), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1072), .A2(new_n1075), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1176), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1174), .B(new_n1175), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1072), .A2(new_n1075), .A3(new_n1179), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1136), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1182), .B(new_n1183), .C1(new_n1184), .C2(new_n1177), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1181), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1171), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(KEYINPUT58), .B(G1341), .ZN(new_n1189));
  OAI22_X1  g764(.A1(new_n1160), .A2(new_n1189), .B1(new_n1076), .B2(G1996), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n546), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1190), .A2(KEYINPUT59), .A3(new_n546), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1188), .A2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1164), .A2(new_n612), .A3(new_n1168), .A4(new_n1166), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1186), .A2(new_n1187), .A3(new_n1171), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1170), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1181), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n1185), .A2(new_n612), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1200), .B1(new_n1201), .B2(new_n1162), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1155), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1153), .A2(KEYINPUT62), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1153), .A2(KEYINPUT62), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1154), .A2(new_n1142), .ZN(new_n1206));
  NOR3_X1   g781(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1131), .A2(new_n1203), .A3(new_n1207), .ZN(new_n1208));
  XOR2_X1   g783(.A(G290), .B(G1986), .Z(new_n1209));
  OAI211_X1 g784(.A(new_n1059), .B(new_n1061), .C1(new_n1044), .C2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1070), .B1(new_n1208), .B2(new_n1210), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n1213));
  NAND2_X1  g787(.A1(new_n665), .A2(G319), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n1214), .A2(KEYINPUT126), .ZN(new_n1215));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n1216));
  NAND3_X1  g790(.A1(new_n665), .A2(new_n1216), .A3(G319), .ZN(new_n1217));
  AOI21_X1  g791(.A(G401), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n693), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g793(.A(new_n1219), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1220));
  AND3_X1   g794(.A1(new_n947), .A2(new_n1213), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g795(.A(new_n1213), .B1(new_n947), .B2(new_n1220), .ZN(new_n1222));
  NOR2_X1   g796(.A1(new_n1221), .A2(new_n1222), .ZN(G308));
  NAND2_X1  g797(.A1(new_n947), .A2(new_n1220), .ZN(new_n1224));
  NAND2_X1  g798(.A1(new_n1224), .A2(KEYINPUT127), .ZN(new_n1225));
  NAND3_X1  g799(.A1(new_n947), .A2(new_n1220), .A3(new_n1213), .ZN(new_n1226));
  NAND2_X1  g800(.A1(new_n1225), .A2(new_n1226), .ZN(G225));
endmodule


