//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT0), .A2(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  OR2_X1    g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n192), .A2(new_n190), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n191), .B1(new_n193), .B2(new_n189), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G125), .ZN(new_n195));
  INV_X1    g009(.A(new_n189), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n197), .B(KEYINPUT1), .C1(new_n198), .C2(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G128), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n197), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n196), .B1(new_n200), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n198), .A2(G146), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n202), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n195), .B1(new_n210), .B2(G125), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n212));
  INV_X1    g026(.A(G224), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G953), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n211), .B(new_n216), .C1(new_n215), .C2(new_n214), .ZN(new_n217));
  INV_X1    g031(.A(G119), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G116), .ZN(new_n219));
  INV_X1    g033(.A(G116), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G119), .ZN(new_n221));
  INV_X1    g035(.A(G113), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n219), .B(new_n221), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n219), .A2(new_n221), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT2), .B(G113), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G104), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G107), .ZN(new_n231));
  INV_X1    g045(.A(G107), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n232), .A2(KEYINPUT3), .A3(G104), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT3), .B1(new_n232), .B2(G104), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n231), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(G101), .ZN(new_n237));
  INV_X1    g051(.A(G101), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n238), .B(new_n231), .C1(new_n233), .C2(new_n234), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT4), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(new_n230), .B2(G107), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n232), .A2(KEYINPUT3), .A3(G104), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n238), .B1(new_n244), .B2(new_n231), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n229), .B(new_n237), .C1(new_n240), .C2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G110), .B(G122), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT74), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n248), .B1(new_n232), .B2(G104), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT73), .B1(new_n230), .B2(G107), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT73), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n232), .A3(G104), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n230), .A2(KEYINPUT74), .A3(G107), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n249), .A2(new_n250), .A3(new_n252), .A4(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G101), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT76), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n256), .B1(new_n219), .B2(KEYINPUT5), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT5), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n259), .A2(new_n218), .A3(KEYINPUT76), .A4(G116), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n257), .A2(new_n258), .A3(G113), .A4(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n255), .A2(new_n261), .A3(new_n225), .A4(new_n239), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n246), .A2(new_n247), .A3(new_n262), .ZN(new_n263));
  OAI221_X1 g077(.A(new_n195), .B1(new_n212), .B2(new_n214), .C1(new_n210), .C2(G125), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n217), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n247), .B(KEYINPUT8), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n255), .A2(new_n239), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n261), .A2(new_n225), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT80), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n255), .A2(new_n225), .A3(new_n239), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n257), .A2(G113), .A3(new_n260), .ZN(new_n272));
  OR2_X1    g086(.A1(new_n272), .A2(KEYINPUT79), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(KEYINPUT79), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n258), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n270), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT80), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n267), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n188), .B1(new_n265), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G210), .B1(G237), .B2(G902), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(KEYINPUT82), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n246), .A2(new_n262), .ZN(new_n282));
  INV_X1    g096(.A(new_n247), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(KEYINPUT6), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(KEYINPUT77), .A3(new_n283), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT6), .A3(new_n263), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT77), .B1(new_n282), .B2(new_n283), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT78), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n245), .A2(new_n236), .B1(new_n228), .B2(new_n225), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n232), .A2(G104), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n242), .B2(new_n243), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n236), .B1(new_n293), .B2(new_n238), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n235), .A2(G101), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n271), .A2(new_n261), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n290), .B1(new_n297), .B2(new_n247), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n263), .A2(KEYINPUT6), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT78), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .A4(new_n286), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n285), .B1(new_n289), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n211), .B(new_n214), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  AOI211_X1 g118(.A(new_n279), .B(new_n281), .C1(new_n302), .C2(new_n304), .ZN(new_n305));
  XOR2_X1   g119(.A(new_n281), .B(KEYINPUT83), .Z(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n285), .ZN(new_n308));
  AOI211_X1 g122(.A(new_n290), .B(new_n247), .C1(new_n246), .C2(new_n262), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n263), .A2(KEYINPUT6), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n300), .B1(new_n311), .B2(new_n298), .ZN(new_n312));
  AND4_X1   g126(.A1(new_n300), .A2(new_n298), .A3(new_n299), .A4(new_n286), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n308), .B(new_n304), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n279), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n307), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n187), .B1(new_n305), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT84), .ZN(new_n318));
  AOI211_X1 g132(.A(new_n285), .B(new_n303), .C1(new_n289), .C2(new_n301), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n306), .B1(new_n319), .B2(new_n279), .ZN(new_n320));
  INV_X1    g134(.A(new_n281), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n314), .A2(new_n315), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT84), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(new_n187), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT16), .ZN(new_n327));
  INV_X1    g141(.A(G140), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(G125), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n329), .B1(new_n333), .B2(new_n327), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n201), .ZN(new_n335));
  OAI211_X1 g149(.A(G146), .B(new_n329), .C1(new_n333), .C2(new_n327), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n218), .B2(G128), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n205), .A2(KEYINPUT23), .A3(G119), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n339), .B(new_n340), .C1(G119), .C2(new_n205), .ZN(new_n341));
  XNOR2_X1  g155(.A(G119), .B(G128), .ZN(new_n342));
  XOR2_X1   g156(.A(KEYINPUT24), .B(G110), .Z(new_n343));
  AOI22_X1  g157(.A1(new_n341), .A2(G110), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n337), .A2(new_n344), .ZN(new_n345));
  OAI22_X1  g159(.A1(new_n341), .A2(G110), .B1(new_n342), .B2(new_n343), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n346), .B(new_n336), .C1(G146), .C2(new_n333), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G137), .ZN(new_n349));
  INV_X1    g163(.A(G953), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(G221), .A3(G234), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n349), .B(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n345), .A2(new_n347), .A3(new_n352), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT72), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT25), .ZN(new_n357));
  AOI21_X1  g171(.A(G902), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n354), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n356), .A2(new_n357), .ZN(new_n360));
  OR2_X1    g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G217), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(G234), .B2(new_n188), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT71), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n359), .B2(new_n360), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n354), .A2(new_n355), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n363), .A2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(KEYINPUT67), .A2(G237), .ZN(new_n371));
  NOR2_X1   g185(.A1(KEYINPUT67), .A2(G237), .ZN(new_n372));
  OAI211_X1 g186(.A(G210), .B(new_n350), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n374));
  XNOR2_X1  g188(.A(new_n373), .B(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT26), .B(G101), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G131), .ZN(new_n379));
  INV_X1    g193(.A(G137), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n380), .A2(G134), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT11), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(G134), .B2(new_n380), .ZN(new_n384));
  INV_X1    g198(.A(G134), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n385), .A2(KEYINPUT11), .A3(G137), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n379), .B(new_n382), .C1(new_n384), .C2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT64), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT11), .B1(new_n385), .B2(G137), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n383), .A2(new_n380), .A3(G134), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n381), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(KEYINPUT64), .A3(new_n379), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n381), .A2(KEYINPUT65), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n380), .A2(G134), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n396), .B1(new_n381), .B2(KEYINPUT65), .ZN(new_n397));
  OAI21_X1  g211(.A(G131), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n394), .A2(new_n209), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n194), .ZN(new_n400));
  INV_X1    g214(.A(new_n392), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G131), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n394), .B2(new_n402), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n399), .A2(new_n403), .A3(new_n229), .ZN(new_n404));
  INV_X1    g218(.A(new_n229), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n387), .A2(new_n388), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT64), .B1(new_n392), .B2(new_n379), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n402), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n194), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n394), .A2(new_n209), .A3(new_n398), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n405), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT28), .B1(new_n404), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n409), .A2(new_n405), .A3(new_n410), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT28), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n378), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n399), .A2(new_n403), .A3(KEYINPUT30), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT30), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n418), .B1(new_n409), .B2(new_n410), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n229), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(new_n378), .A3(new_n413), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT31), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT30), .B1(new_n399), .B2(new_n403), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n409), .A2(new_n418), .A3(new_n410), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n404), .B1(new_n426), .B2(new_n229), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT31), .A3(new_n378), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n416), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(G472), .A2(G902), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT32), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n416), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT31), .B1(new_n427), .B2(new_n378), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n405), .B1(new_n424), .B2(new_n425), .ZN(new_n435));
  NOR4_X1   g249(.A1(new_n435), .A2(new_n422), .A3(new_n377), .A4(new_n404), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n433), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT32), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n430), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n412), .A2(new_n378), .A3(new_n415), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT29), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(G902), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT69), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n412), .A2(KEYINPUT69), .A3(new_n378), .A4(new_n415), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n442), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT70), .B1(new_n427), .B2(new_n378), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT70), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n450), .B(new_n377), .C1(new_n435), .C2(new_n404), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n444), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G472), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n370), .B1(new_n440), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n220), .A2(G122), .ZN(new_n456));
  INV_X1    g270(.A(G122), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(G116), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(new_n232), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n198), .A2(G128), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT13), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n205), .A2(G143), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n461), .A2(new_n462), .ZN(new_n466));
  OAI21_X1  g280(.A(G134), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n461), .A2(new_n464), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n385), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n460), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT14), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n458), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT90), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n456), .B1(new_n471), .B2(new_n458), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n232), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n468), .B(new_n385), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n459), .A2(new_n232), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n470), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT9), .B(G234), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n480), .A2(new_n362), .A3(G953), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n470), .B(new_n481), .C1(new_n475), .C2(new_n478), .ZN(new_n484));
  AOI21_X1  g298(.A(G902), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G478), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(KEYINPUT15), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n485), .B(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G952), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n489), .A2(KEYINPUT91), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(KEYINPUT91), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n350), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n492), .B1(G234), .B2(G237), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT21), .B(G898), .ZN(new_n494));
  AOI211_X1 g308(.A(new_n188), .B(new_n350), .C1(G234), .C2(G237), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n488), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G469), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n209), .A2(KEYINPUT10), .A3(new_n239), .A4(new_n255), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n205), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n208), .B1(new_n501), .B2(new_n189), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n255), .A2(new_n502), .A3(new_n239), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT10), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n194), .B(new_n237), .C1(new_n240), .C2(new_n245), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n389), .A2(new_n393), .B1(G131), .B2(new_n401), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n500), .A2(new_n505), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(G110), .B(G140), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n350), .A2(G227), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n509), .B(new_n510), .Z(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n255), .A2(new_n239), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n503), .B1(new_n514), .B2(new_n209), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT75), .B1(new_n394), .B2(new_n402), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT12), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n517), .B1(new_n515), .B2(new_n516), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n513), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n500), .A2(new_n506), .A3(new_n505), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n408), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n512), .B1(new_n522), .B2(new_n508), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n499), .B(new_n188), .C1(new_n520), .C2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n513), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n522), .ZN(new_n526));
  INV_X1    g340(.A(new_n508), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n518), .A2(new_n527), .A3(new_n519), .ZN(new_n528));
  OAI211_X1 g342(.A(G469), .B(new_n526), .C1(new_n528), .C2(new_n512), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n499), .A2(new_n188), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n524), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(G221), .B1(new_n480), .B2(G902), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT89), .ZN(new_n535));
  NOR2_X1   g349(.A1(G475), .A2(G902), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G113), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(new_n230), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n333), .B(KEYINPUT19), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n336), .B1(new_n541), .B2(G146), .ZN(new_n542));
  OAI211_X1 g356(.A(G214), .B(new_n350), .C1(new_n371), .C2(new_n372), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n198), .ZN(new_n544));
  AND2_X1   g358(.A1(G143), .A2(G214), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n350), .B(new_n545), .C1(new_n371), .C2(new_n372), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n379), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n379), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n198), .B2(new_n543), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT86), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n544), .A2(new_n379), .A3(new_n546), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT86), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n542), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n333), .B(new_n201), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n544), .A2(KEYINPUT85), .A3(new_n546), .ZN(new_n556));
  NAND2_X1  g370(.A1(KEYINPUT18), .A2(G131), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n555), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n544), .A2(KEYINPUT85), .A3(new_n557), .A4(new_n546), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n540), .B1(new_n554), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n544), .A2(new_n546), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G131), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT17), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n544), .A2(new_n550), .A3(new_n379), .A4(new_n546), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n553), .A2(new_n564), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n337), .B1(KEYINPUT17), .B2(new_n547), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n559), .A2(new_n560), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n539), .B(KEYINPUT87), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n537), .B1(new_n562), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT88), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT20), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI211_X1 g389(.A(KEYINPUT88), .B(new_n537), .C1(new_n562), .C2(new_n572), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT20), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n553), .A2(new_n564), .A3(new_n566), .ZN(new_n579));
  INV_X1    g393(.A(new_n542), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n570), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n567), .A2(new_n568), .B1(new_n560), .B2(new_n559), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n540), .A2(new_n582), .B1(new_n583), .B2(new_n571), .ZN(new_n584));
  OAI211_X1 g398(.A(KEYINPUT88), .B(new_n578), .C1(new_n584), .C2(new_n537), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n539), .B1(new_n569), .B2(new_n570), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n188), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G475), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n535), .B1(new_n577), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT88), .B1(new_n584), .B2(new_n537), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n573), .A2(new_n574), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(KEYINPUT20), .A3(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n594), .A2(KEYINPUT89), .A3(new_n585), .A4(new_n589), .ZN(new_n595));
  AOI211_X1 g409(.A(new_n498), .B(new_n534), .C1(new_n591), .C2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n326), .A2(new_n455), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  AOI21_X1  g412(.A(new_n321), .B1(new_n314), .B2(new_n315), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n187), .B(new_n497), .C1(new_n305), .C2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n486), .A2(new_n188), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n485), .A2(new_n486), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n483), .A2(new_n484), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(new_n605));
  AOI211_X1 g419(.A(new_n601), .B(new_n602), .C1(new_n605), .C2(G478), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n591), .A2(new_n595), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G472), .B1(new_n429), .B2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n437), .A2(new_n430), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n533), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n515), .A2(new_n516), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT12), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n508), .A3(new_n616), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n617), .A2(new_n511), .B1(new_n522), .B2(new_n525), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n530), .B1(new_n618), .B2(G469), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n613), .B1(new_n619), .B2(new_n524), .ZN(new_n620));
  INV_X1    g434(.A(new_n370), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n612), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n609), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT34), .B(G104), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  NOR2_X1   g440(.A1(new_n577), .A2(new_n590), .ZN(new_n627));
  INV_X1    g441(.A(new_n488), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n600), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n623), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT35), .B(G107), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NOR3_X1   g448(.A1(new_n348), .A2(KEYINPUT36), .A3(new_n353), .ZN(new_n635));
  INV_X1    g449(.A(new_n368), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT36), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n345), .A2(new_n347), .B1(new_n637), .B2(new_n352), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n361), .B2(new_n365), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n610), .A2(new_n611), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n317), .A2(KEYINPUT84), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n324), .B1(new_n323), .B2(new_n187), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n596), .B(new_n642), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT37), .B(G110), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G12));
  AOI21_X1  g461(.A(new_n640), .B1(new_n440), .B2(new_n454), .ZN(new_n648));
  INV_X1    g462(.A(new_n187), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n281), .B1(new_n319), .B2(new_n279), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n649), .B1(new_n650), .B2(new_n322), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n620), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n573), .A2(new_n574), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n655), .A2(new_n578), .B1(G475), .B2(new_n588), .ZN(new_n656));
  INV_X1    g470(.A(new_n493), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT92), .B(G900), .Z(new_n658));
  NAND2_X1  g472(.A1(new_n495), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n656), .A2(new_n594), .A3(new_n628), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT93), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n654), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  NOR2_X1   g478(.A1(new_n305), .A2(new_n316), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n427), .A2(new_n377), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n229), .B1(new_n399), .B2(new_n403), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n377), .A3(new_n413), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n188), .ZN(new_n673));
  OAI21_X1  g487(.A(G472), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n440), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n591), .A2(new_n595), .A3(new_n628), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n669), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n660), .B(KEYINPUT39), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n620), .A2(new_n678), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n187), .B(new_n640), .C1(new_n679), .C2(KEYINPUT40), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(KEYINPUT40), .B2(new_n679), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  AND4_X1   g497(.A1(new_n591), .A2(new_n595), .A3(new_n606), .A4(new_n660), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n654), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  OAI21_X1  g500(.A(new_n188), .B1(new_n520), .B2(new_n523), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G469), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n533), .A3(new_n524), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(KEYINPUT95), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT95), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n688), .A2(new_n691), .A3(new_n533), .A4(new_n524), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n455), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n694), .A2(new_n609), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT41), .B(G113), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NOR2_X1   g511(.A1(new_n694), .A2(new_n631), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(new_n220), .ZN(G18));
  AOI21_X1  g513(.A(new_n498), .B1(new_n591), .B2(new_n595), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n187), .B1(new_n305), .B2(new_n599), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n701), .A2(KEYINPUT96), .A3(new_n689), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT96), .ZN(new_n703));
  INV_X1    g517(.A(new_n689), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n703), .B1(new_n651), .B2(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n700), .B(new_n648), .C1(new_n702), .C2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G119), .ZN(G21));
  AOI21_X1  g521(.A(new_n414), .B1(new_n671), .B2(new_n413), .ZN(new_n708));
  INV_X1    g522(.A(new_n415), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT97), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n377), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n708), .A2(new_n709), .A3(KEYINPUT97), .ZN(new_n712));
  OAI22_X1  g526(.A1(new_n711), .A2(new_n712), .B1(new_n434), .B2(new_n436), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n430), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n610), .A2(new_n714), .A3(new_n621), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n690), .A2(new_n497), .A3(new_n692), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT98), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n701), .B1(new_n676), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n591), .A2(new_n595), .A3(KEYINPUT98), .A4(new_n628), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n717), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NAND3_X1  g536(.A1(new_n610), .A2(new_n714), .A3(new_n641), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n591), .A2(new_n595), .A3(new_n606), .A4(new_n660), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n702), .B2(new_n705), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT99), .B(G125), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G27));
  NAND2_X1  g542(.A1(new_n440), .A2(new_n454), .ZN(new_n729));
  AND4_X1   g543(.A1(new_n187), .A2(new_n320), .A3(new_n620), .A4(new_n322), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n729), .A2(new_n684), .A3(new_n730), .A4(new_n621), .ZN(new_n731));
  NOR2_X1   g545(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n732), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n455), .A2(new_n684), .A3(new_n730), .A4(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G131), .ZN(G33));
  AND3_X1   g551(.A1(new_n455), .A2(new_n662), .A3(new_n730), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n385), .ZN(G36));
  AND2_X1   g553(.A1(new_n618), .A2(KEYINPUT45), .ZN(new_n740));
  OAI21_X1  g554(.A(G469), .B1(new_n618), .B2(KEYINPUT45), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT101), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n530), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n744), .A2(KEYINPUT46), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n524), .B1(new_n744), .B2(KEYINPUT46), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n533), .B(new_n678), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n612), .A2(new_n641), .ZN(new_n749));
  XOR2_X1   g563(.A(new_n749), .B(KEYINPUT103), .Z(new_n750));
  NAND2_X1  g564(.A1(new_n591), .A2(new_n595), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n606), .ZN(new_n752));
  NOR2_X1   g566(.A1(KEYINPUT102), .A2(KEYINPUT43), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(KEYINPUT102), .A2(KEYINPUT43), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n752), .B1(new_n755), .B2(new_n753), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n750), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n747), .B1(new_n748), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n665), .A2(new_n187), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT104), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n759), .B(new_n761), .C1(new_n748), .C2(new_n758), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  OAI21_X1  g577(.A(new_n533), .B1(new_n745), .B2(new_n746), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI211_X1 g580(.A(KEYINPUT47), .B(new_n533), .C1(new_n745), .C2(new_n746), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n729), .A2(new_n621), .A3(new_n760), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n684), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  NAND3_X1  g585(.A1(new_n621), .A2(new_n187), .A3(new_n533), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n688), .A2(new_n524), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n772), .B1(new_n773), .B2(KEYINPUT49), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n751), .A3(new_n606), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT105), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n773), .A2(KEYINPUT49), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n776), .A2(new_n669), .A3(new_n675), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n492), .B(KEYINPUT115), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n760), .A2(new_n689), .ZN(new_n780));
  AND4_X1   g594(.A1(new_n621), .A2(new_n780), .A3(new_n675), .A4(new_n493), .ZN(new_n781));
  INV_X1    g595(.A(new_n607), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n657), .B1(new_n754), .B2(new_n756), .ZN(new_n784));
  INV_X1    g598(.A(new_n715), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n702), .A2(new_n705), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT116), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT48), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n784), .A2(new_n780), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT113), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n784), .A2(new_n793), .A3(new_n780), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n790), .B1(new_n795), .B2(new_n455), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n795), .A2(new_n790), .A3(new_n455), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n789), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n689), .A2(new_n187), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n669), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n669), .A2(KEYINPUT112), .A3(new_n800), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n799), .B1(new_n805), .B2(new_n786), .ZN(new_n806));
  INV_X1    g620(.A(new_n786), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n807), .A2(KEYINPUT50), .A3(new_n804), .A4(new_n803), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n606), .B1(new_n591), .B2(new_n595), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n781), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n723), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT114), .B1(new_n795), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n814), .B(new_n723), .C1(new_n792), .C2(new_n794), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n809), .B(new_n811), .C1(new_n813), .C2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n688), .A2(new_n613), .A3(new_n524), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n766), .A2(new_n767), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n761), .ZN(new_n820));
  OR3_X1    g634(.A1(new_n786), .A2(KEYINPUT110), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT110), .B1(new_n786), .B2(new_n820), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n823), .A2(KEYINPUT51), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n798), .B1(new_n817), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(KEYINPUT109), .B(KEYINPUT51), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n823), .A2(KEYINPUT111), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n819), .A2(new_n828), .A3(new_n821), .A4(new_n822), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n826), .B1(new_n830), .B2(new_n816), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n825), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n738), .B1(new_n733), .B2(new_n735), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n455), .B(new_n693), .C1(new_n608), .C2(new_n630), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n488), .B(KEYINPUT106), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n751), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n607), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n612), .A2(new_n496), .A3(new_n622), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n326), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n834), .A2(new_n706), .A3(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n597), .A2(new_n721), .A3(new_n645), .ZN(new_n841));
  INV_X1    g655(.A(new_n730), .ZN(new_n842));
  INV_X1    g656(.A(new_n660), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n835), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n729), .A2(new_n627), .A3(new_n641), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n725), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n833), .A2(new_n840), .A3(new_n841), .A4(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n648), .B(new_n653), .C1(new_n662), .C2(new_n684), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n843), .B(new_n639), .C1(new_n361), .C2(new_n365), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n620), .A2(KEYINPUT107), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n532), .A2(new_n851), .A3(new_n533), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT107), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n440), .A2(new_n674), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n719), .A3(new_n720), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n850), .A2(new_n726), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n850), .A2(new_n726), .A3(new_n857), .A4(KEYINPUT52), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT53), .B1(new_n849), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n834), .A2(new_n706), .A3(new_n839), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n597), .A2(new_n721), .A3(new_n645), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n864), .A2(new_n865), .A3(new_n847), .ZN(new_n866));
  AND4_X1   g680(.A1(KEYINPUT53), .A2(new_n862), .A3(new_n866), .A4(new_n833), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT54), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n860), .A2(new_n861), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n840), .A2(new_n833), .A3(new_n841), .A4(new_n848), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n862), .A2(new_n866), .A3(KEYINPUT53), .A4(new_n833), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n868), .A2(KEYINPUT108), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT108), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n832), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(G952), .A2(G953), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n778), .B1(new_n881), .B2(new_n882), .ZN(G75));
  NOR2_X1   g697(.A1(new_n350), .A2(G952), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT119), .Z(new_n885));
  AOI21_X1  g699(.A(new_n188), .B1(new_n872), .B2(new_n874), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT56), .B1(new_n886), .B2(new_n281), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n302), .A2(new_n304), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n319), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT55), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n885), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n890), .B(KEYINPUT117), .Z(new_n892));
  AOI211_X1 g706(.A(KEYINPUT56), .B(new_n892), .C1(new_n886), .C2(new_n306), .ZN(new_n893));
  OR2_X1    g707(.A1(new_n893), .A2(KEYINPUT118), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(KEYINPUT118), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(G51));
  NAND2_X1  g710(.A1(new_n872), .A2(new_n874), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT120), .B1(new_n897), .B2(KEYINPUT54), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n868), .A2(new_n875), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n899), .B2(KEYINPUT120), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n530), .B(KEYINPUT57), .Z(new_n901));
  OAI22_X1  g715(.A1(new_n900), .A2(new_n901), .B1(new_n523), .B2(new_n520), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n886), .A2(new_n743), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n884), .B1(new_n902), .B2(new_n903), .ZN(G54));
  INV_X1    g718(.A(new_n584), .ZN(new_n905));
  AND2_X1   g719(.A1(KEYINPUT58), .A2(G475), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n886), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n905), .B1(new_n886), .B2(new_n906), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n907), .A2(new_n908), .A3(new_n884), .ZN(G60));
  XOR2_X1   g723(.A(new_n601), .B(KEYINPUT59), .Z(new_n910));
  NAND3_X1  g724(.A1(new_n880), .A2(new_n876), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n605), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT122), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n911), .A2(new_n914), .A3(new_n605), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n916));
  INV_X1    g730(.A(new_n605), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n910), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT120), .B1(new_n878), .B2(new_n879), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n868), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n918), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n885), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n916), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(KEYINPUT121), .B(new_n885), .C1(new_n900), .C2(new_n918), .ZN(new_n925));
  AOI22_X1  g739(.A1(new_n913), .A2(new_n915), .B1(new_n924), .B2(new_n925), .ZN(G63));
  NOR2_X1   g740(.A1(new_n635), .A2(new_n638), .ZN(new_n927));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT123), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT60), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n897), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n897), .A2(new_n930), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n885), .B(new_n931), .C1(new_n932), .C2(new_n367), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g748(.A(G953), .B1(new_n494), .B2(new_n213), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n840), .A2(new_n841), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n936), .A2(KEYINPUT124), .A3(new_n350), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT124), .B1(new_n936), .B2(new_n350), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n302), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(G898), .B2(new_n350), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n940), .B(new_n942), .ZN(G69));
  XOR2_X1   g757(.A(new_n541), .B(KEYINPUT125), .Z(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT126), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(new_n426), .ZN(new_n946));
  NAND2_X1  g760(.A1(G900), .A2(G953), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n719), .A2(new_n455), .A3(new_n720), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n747), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n850), .A2(new_n726), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n762), .A2(new_n770), .A3(new_n833), .A4(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n946), .B(new_n947), .C1(new_n952), .C2(G953), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n837), .A2(new_n455), .A3(new_n678), .A4(new_n730), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n762), .A2(new_n770), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n950), .B1(new_n677), .B2(new_n681), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT62), .ZN(new_n957));
  AOI21_X1  g771(.A(G953), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n953), .B1(new_n958), .B2(new_n946), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n350), .B1(G227), .B2(G900), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n960), .B1(new_n953), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n959), .A2(new_n962), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(G72));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n952), .B2(new_n936), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n435), .A2(new_n378), .A3(new_n404), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n884), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n449), .A2(new_n451), .A3(new_n421), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n897), .A2(new_n967), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n955), .A2(new_n957), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n967), .B1(new_n974), .B2(new_n936), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n973), .B1(new_n670), .B2(new_n975), .ZN(G57));
endmodule


