//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n450, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1139;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  INV_X1    g024(.A(G567), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT67), .Z(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT68), .Z(new_n455));
  NOR4_X1   g030(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT2), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G325));
  XOR2_X1   g034(.A(new_n458), .B(KEYINPUT69), .Z(G261));
  OR2_X1    g035(.A1(new_n455), .A2(new_n450), .ZN(new_n461));
  INV_X1    g036(.A(new_n457), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2106), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n466), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OR2_X1    g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n466), .A2(G137), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n472), .A2(new_n470), .B1(G101), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  INV_X1    g052(.A(new_n466), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n470), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(G124), .A2(new_n479), .B1(new_n480), .B2(G136), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n470), .C2(G112), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND3_X1  g059(.A1(new_n466), .A2(G126), .A3(G2105), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n486));
  OR2_X1    g061(.A1(new_n486), .A2(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(G114), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n473), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(new_n491), .A2(KEYINPUT72), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n470), .A2(new_n466), .A3(G138), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n470), .A2(new_n466), .A3(new_n495), .A4(G138), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n491), .A2(KEYINPUT72), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n492), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  XNOR2_X1  g075(.A(KEYINPUT73), .B(G651), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT75), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n507), .A2(G62), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  XOR2_X1   g084(.A(new_n509), .B(KEYINPUT78), .Z(new_n510));
  OAI21_X1  g085(.A(new_n502), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n505), .A2(new_n506), .B1(new_n512), .B2(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n514), .B1(new_n501), .B2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  AND4_X1   g094(.A1(new_n514), .A2(new_n517), .A3(new_n519), .A4(KEYINPUT6), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n513), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT76), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n517), .A2(new_n519), .A3(KEYINPUT6), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT74), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n501), .A2(new_n514), .A3(KEYINPUT6), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT76), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n526), .A2(new_n527), .A3(new_n513), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n522), .A2(G88), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT77), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n504), .B1(new_n512), .B2(G651), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G50), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n529), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n530), .B1(new_n529), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n511), .B1(new_n534), .B2(new_n535), .ZN(G303));
  INV_X1    g111(.A(G303), .ZN(G166));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n526), .A2(new_n531), .ZN(new_n541));
  INV_X1    g116(.A(G51), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n522), .A2(new_n528), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n543), .B1(new_n544), .B2(G89), .ZN(G168));
  NAND2_X1  g120(.A1(new_n544), .A2(G90), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(new_n507), .ZN(new_n548));
  INV_X1    g123(.A(G64), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n532), .A2(G52), .B1(new_n502), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n546), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND3_X1  g128(.A1(new_n522), .A2(G81), .A3(new_n528), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n532), .A2(G43), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n554), .A2(KEYINPUT79), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n501), .ZN(new_n562));
  AOI21_X1  g137(.A(KEYINPUT80), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  AND3_X1   g138(.A1(new_n554), .A2(KEYINPUT79), .A3(new_n555), .ZN(new_n564));
  AOI21_X1  g139(.A(KEYINPUT79), .B1(new_n554), .B2(new_n555), .ZN(new_n565));
  OAI211_X1 g140(.A(KEYINPUT80), .B(new_n562), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n548), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n544), .A2(G91), .B1(G651), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(G53), .ZN(new_n578));
  OR3_X1    g153(.A1(new_n541), .A2(KEYINPUT9), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT9), .B1(new_n541), .B2(new_n578), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G168), .ZN(G286));
  NAND2_X1  g158(.A1(new_n544), .A2(G87), .ZN(new_n584));
  INV_X1    g159(.A(G74), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n516), .B1(new_n548), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n532), .B2(G49), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(new_n544), .A2(G86), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n507), .A2(G61), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT81), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n501), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n595), .A2(new_n596), .B1(new_n532), .B2(G48), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n589), .A2(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n532), .A2(G47), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n522), .A2(new_n528), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI221_X1 g177(.A(new_n599), .B1(new_n501), .B2(new_n600), .C1(new_n601), .C2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n522), .A2(G92), .A3(new_n528), .ZN(new_n605));
  XNOR2_X1  g180(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT84), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n516), .B1(new_n609), .B2(new_n610), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n532), .A2(G54), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n607), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n604), .B1(new_n615), .B2(G868), .ZN(G321));
  XNOR2_X1  g191(.A(G321), .B(KEYINPUT85), .ZN(G284));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(G299), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G297));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G280));
  INV_X1    g196(.A(G860), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n614), .B1(G559), .B2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT86), .Z(G148));
  NOR2_X1   g199(.A1(new_n614), .A2(G559), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n568), .B2(G868), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n470), .A2(G111), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(KEYINPUT88), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(KEYINPUT88), .B2(new_n631), .ZN(new_n633));
  AOI22_X1  g208(.A1(G123), .A2(new_n479), .B1(new_n480), .B2(G135), .ZN(new_n634));
  AND2_X1   g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n466), .A2(new_n474), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT87), .B(KEYINPUT13), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n636), .A2(G2096), .B1(G2100), .B2(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(G2100), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n641), .B(new_n642), .C1(G2096), .C2(new_n636), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT89), .Z(G156));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n650), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  AND3_X1   g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(G401));
  NOR2_X1   g234(.A1(G2072), .A2(G2078), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n442), .A2(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n661), .A2(KEYINPUT90), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(KEYINPUT90), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n661), .B(KEYINPUT17), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n666), .B(new_n668), .C1(new_n665), .C2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT91), .Z(new_n671));
  NOR3_X1   g246(.A1(new_n668), .A2(new_n661), .A3(new_n665), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT18), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n665), .A3(new_n667), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2096), .B(G2100), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n679), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(new_n682), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT20), .Z(new_n686));
  AOI211_X1 g261(.A(new_n684), .B(new_n686), .C1(new_n679), .C2(new_n683), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT92), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G229));
  INV_X1    g269(.A(KEYINPUT101), .ZN(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G23), .ZN(new_n697));
  INV_X1    g272(.A(G288), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT33), .B(G1976), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n589), .A2(new_n597), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G16), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G6), .B2(G16), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(KEYINPUT32), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(KEYINPUT32), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G1981), .ZN(new_n708));
  INV_X1    g283(.A(G1981), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n705), .A2(new_n709), .A3(new_n706), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n701), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(G16), .A2(G22), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G166), .B2(G16), .ZN(new_n713));
  INV_X1    g288(.A(G1971), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT34), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n711), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  MUX2_X1   g292(.A(G24), .B(G290), .S(G16), .Z(new_n718));
  AND2_X1   g293(.A1(new_n718), .A2(G1986), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(G1986), .ZN(new_n720));
  AOI22_X1  g295(.A1(G119), .A2(new_n479), .B1(new_n480), .B2(G131), .ZN(new_n721));
  OAI221_X1 g296(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n470), .C2(G107), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G25), .B(new_n723), .S(G29), .Z(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n724), .B(new_n726), .ZN(new_n727));
  NOR3_X1   g302(.A1(new_n719), .A2(new_n720), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n717), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n716), .B1(new_n711), .B2(new_n715), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT93), .B(KEYINPUT36), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OR3_X1    g307(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n729), .B2(new_n730), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G32), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n480), .A2(G141), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT96), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n479), .A2(G129), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT26), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n743), .A2(new_n744), .B1(G105), .B2(new_n474), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n739), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n737), .B1(new_n748), .B2(new_n736), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT97), .ZN(new_n753));
  INV_X1    g328(.A(G2078), .ZN(new_n754));
  NOR2_X1   g329(.A1(G164), .A2(new_n736), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G27), .B2(new_n736), .ZN(new_n756));
  OAI22_X1  g331(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT31), .B(G11), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n736), .B1(new_n759), .B2(G28), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n760), .A2(KEYINPUT98), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(G28), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n760), .B2(KEYINPUT98), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n758), .B1(new_n761), .B2(new_n763), .C1(new_n636), .C2(new_n736), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT99), .Z(new_n765));
  AOI211_X1 g340(.A(new_n757), .B(new_n765), .C1(new_n753), .C2(new_n752), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n756), .A2(new_n754), .ZN(new_n767));
  INV_X1    g342(.A(G34), .ZN(new_n768));
  AOI21_X1  g343(.A(G29), .B1(new_n768), .B2(KEYINPUT24), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(KEYINPUT24), .B2(new_n768), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n476), .B2(new_n736), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2084), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n767), .B(new_n772), .C1(new_n750), .C2(new_n751), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT25), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n480), .A2(G139), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n775), .B(new_n776), .C1(new_n470), .C2(new_n777), .ZN(new_n778));
  MUX2_X1   g353(.A(G33), .B(new_n778), .S(G29), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2072), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n736), .A2(G35), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G162), .B2(new_n736), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT29), .B(G2090), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n736), .A2(G26), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT28), .Z(new_n786));
  AOI22_X1  g361(.A1(G128), .A2(new_n479), .B1(new_n480), .B2(G140), .ZN(new_n787));
  OAI221_X1 g362(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n470), .C2(G116), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n786), .B1(new_n789), .B2(G29), .ZN(new_n790));
  INV_X1    g365(.A(G2067), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR4_X1   g367(.A1(new_n773), .A2(new_n780), .A3(new_n784), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n696), .A2(G20), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT23), .Z(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G299), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT100), .B(G1956), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n766), .A2(new_n793), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n568), .A2(new_n696), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n696), .A2(G19), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT95), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G1341), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n615), .A2(G16), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G4), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT94), .B(G1348), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n807), .A2(new_n809), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n696), .A2(G5), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G171), .B2(new_n696), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G1961), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n696), .A2(G21), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G168), .B2(new_n696), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n814), .A2(new_n815), .B1(G1966), .B2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n817), .ZN(new_n819));
  INV_X1    g394(.A(G1966), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n813), .A2(G1961), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n810), .A2(new_n811), .A3(new_n818), .A4(new_n821), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n800), .A2(new_n805), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n695), .B1(new_n735), .B2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n823), .ZN(new_n825));
  AOI211_X1 g400(.A(KEYINPUT101), .B(new_n825), .C1(new_n733), .C2(new_n734), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n824), .A2(new_n826), .ZN(G311));
  NAND2_X1  g402(.A1(new_n735), .A2(new_n823), .ZN(G150));
  NAND2_X1  g403(.A1(new_n615), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n829), .B(new_n830), .Z(new_n831));
  AOI22_X1  g406(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n501), .B1(new_n832), .B2(KEYINPUT102), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(KEYINPUT102), .B2(new_n832), .ZN(new_n834));
  INV_X1    g409(.A(G55), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n541), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G93), .B2(new_n544), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n563), .B2(new_n567), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n560), .A2(new_n562), .A3(new_n837), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n831), .B(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n843), .A2(new_n622), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n838), .A2(G860), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT104), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n848), .ZN(G145));
  XNOR2_X1  g424(.A(new_n483), .B(new_n476), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n635), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT106), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n778), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n748), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n789), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n491), .B1(new_n497), .B2(KEYINPUT105), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(KEYINPUT105), .B2(new_n497), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n855), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n723), .B(new_n638), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n470), .A2(G118), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT107), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  AOI22_X1  g439(.A1(G130), .A2(new_n479), .B1(new_n480), .B2(G142), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n859), .B(new_n866), .Z(new_n867));
  AOI21_X1  g442(.A(new_n851), .B1(new_n858), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n858), .B2(new_n867), .ZN(new_n869));
  INV_X1    g444(.A(G37), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT108), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n858), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n858), .A2(new_n872), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n851), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n869), .B(new_n870), .C1(new_n873), .C2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g452(.A(new_n841), .B(new_n626), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n614), .A2(G299), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n608), .A2(new_n613), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n880), .A2(new_n581), .A3(new_n577), .A4(new_n607), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n879), .A2(new_n881), .A3(KEYINPUT41), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(new_n879), .B2(new_n881), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n883), .B1(new_n886), .B2(new_n878), .ZN(new_n887));
  XNOR2_X1  g462(.A(G305), .B(G290), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(G303), .A2(new_n698), .ZN(new_n890));
  OAI211_X1 g465(.A(G288), .B(new_n511), .C1(new_n534), .C2(new_n535), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT42), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT109), .ZN(new_n896));
  INV_X1    g471(.A(new_n894), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n893), .A2(KEYINPUT109), .A3(new_n894), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n895), .B1(new_n901), .B2(KEYINPUT42), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n887), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(G868), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(G868), .B2(new_n837), .ZN(G295));
  OAI21_X1  g480(.A(new_n904), .B1(G868), .B2(new_n837), .ZN(G331));
  INV_X1    g481(.A(new_n882), .ZN(new_n907));
  XNOR2_X1  g482(.A(G301), .B(G168), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n909), .B1(new_n839), .B2(new_n840), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT80), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n837), .B1(new_n913), .B2(new_n566), .ZN(new_n914));
  INV_X1    g489(.A(new_n840), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n914), .A2(new_n915), .A3(new_n908), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n907), .B1(new_n910), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n839), .A2(new_n840), .A3(new_n909), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n908), .B1(new_n914), .B2(new_n915), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n886), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT110), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(KEYINPUT110), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n901), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n918), .A2(new_n919), .A3(new_n886), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n882), .B1(new_n918), .B2(new_n919), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n901), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n929), .A3(new_n922), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(new_n930), .A3(new_n870), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT111), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n931), .A2(new_n934), .A3(KEYINPUT43), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n901), .B1(new_n926), .B2(new_n927), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n901), .B(KEYINPUT112), .C1(new_n926), .C2(new_n927), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n930), .A2(new_n938), .A3(new_n870), .A4(new_n939), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n933), .A2(new_n935), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  INV_X1    g520(.A(new_n939), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n917), .A2(new_n920), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT112), .B1(new_n947), .B2(new_n901), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT113), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n949), .A2(new_n950), .A3(new_n870), .A4(new_n930), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n940), .A2(KEYINPUT113), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n945), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n931), .A2(new_n945), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT44), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n944), .A2(new_n955), .ZN(G397));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n857), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g534(.A1(G160), .A2(G40), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT114), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n958), .A2(KEYINPUT114), .A3(new_n959), .A4(new_n961), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n789), .B(new_n791), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n966), .B1(new_n748), .B2(new_n967), .ZN(new_n968));
  OR3_X1    g543(.A1(new_n966), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT46), .B1(new_n966), .B2(G1996), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT47), .ZN(new_n972));
  INV_X1    g547(.A(new_n966), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(G1996), .A3(new_n747), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT115), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n967), .B1(G1996), .B2(new_n747), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n723), .A2(new_n726), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n787), .A2(new_n791), .A3(new_n788), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n966), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n725), .B1(new_n721), .B2(new_n722), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n973), .B1(new_n982), .B2(new_n978), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n977), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n966), .A2(G1986), .A3(G290), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n986), .B(KEYINPUT48), .Z(new_n987));
  AOI211_X1 g562(.A(new_n972), .B(new_n981), .C1(new_n985), .C2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n702), .A2(new_n709), .ZN(new_n989));
  NAND2_X1  g564(.A1(G305), .A2(G1981), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT49), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(KEYINPUT49), .A3(new_n990), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n958), .A2(new_n960), .ZN(new_n995));
  INV_X1    g570(.A(G8), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n993), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n698), .A2(G1976), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT52), .ZN(new_n1001));
  INV_X1    g576(.A(G1976), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT52), .B1(G288), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n997), .A2(new_n999), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n998), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT116), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n998), .B2(new_n1005), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G303), .A2(G8), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT55), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n499), .A2(new_n957), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1015), .B(new_n961), .C1(KEYINPUT50), .C2(new_n958), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1016), .A2(G2090), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n959), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1018), .B(new_n961), .C1(new_n958), .C2(new_n959), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n714), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n996), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1013), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT63), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1015), .A2(new_n961), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n958), .A2(KEYINPUT50), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G2084), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n960), .B1(new_n958), .B2(new_n959), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n957), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n820), .ZN(new_n1034));
  AOI211_X1 g609(.A(new_n996), .B(G286), .C1(new_n1030), .C2(new_n1034), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1013), .A2(new_n1021), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1010), .A2(new_n1025), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n958), .A2(KEYINPUT50), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(new_n961), .C1(KEYINPUT50), .C2(new_n1014), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1020), .B1(G2090), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G8), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n1012), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1006), .A2(new_n1022), .A3(new_n1042), .A4(new_n1035), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1043), .A2(KEYINPUT118), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1024), .B1(new_n1043), .B2(KEYINPUT118), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1037), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n1019), .B2(G2078), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1016), .A2(new_n815), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n857), .A2(new_n957), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT45), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1052), .A2(new_n1031), .A3(KEYINPUT53), .A4(new_n754), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1047), .B1(new_n1054), .B2(G171), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1031), .A2(KEYINPUT53), .A3(new_n754), .A4(new_n1032), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1049), .A2(new_n1056), .A3(new_n1050), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1055), .B1(G171), .B2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1058), .A2(new_n1022), .A3(new_n1042), .A4(new_n1006), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1060), .A2(new_n996), .A3(G168), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1030), .A2(new_n1034), .A3(G168), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT124), .B(KEYINPUT51), .Z(new_n1063));
  AND3_X1   g638(.A1(new_n1062), .A2(G8), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n1062), .B2(G8), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1061), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n619), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(G299), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT121), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1076), .A3(new_n1073), .ZN(new_n1077));
  INV_X1    g652(.A(G1956), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1039), .A2(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT56), .B(G2072), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1052), .A2(new_n1018), .A3(new_n961), .A4(new_n1080), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1075), .A2(new_n1077), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  AND4_X1   g657(.A1(new_n1079), .A2(new_n1081), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(new_n614), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n995), .A2(new_n791), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT120), .ZN(new_n1086));
  INV_X1    g661(.A(G1348), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1016), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n995), .A2(new_n1089), .A3(new_n791), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1086), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1082), .B1(new_n1084), .B2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1079), .A2(new_n1081), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1083), .B2(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT58), .B(G1341), .ZN(new_n1096));
  OAI22_X1  g671(.A1(new_n1019), .A2(G1996), .B1(new_n995), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n568), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1086), .A2(new_n1088), .A3(KEYINPUT60), .A4(new_n1090), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1101), .A2(new_n615), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1095), .A2(new_n1100), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT60), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1091), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1106), .A2(new_n615), .A3(new_n1101), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT61), .B1(new_n1108), .B2(new_n1074), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1107), .B1(new_n1082), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1092), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1057), .A2(G171), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1112), .B(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT126), .ZN(new_n1115));
  OR3_X1    g690(.A1(new_n1054), .A2(new_n1115), .A3(G171), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(new_n1054), .B2(G171), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1047), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1068), .A2(new_n1111), .A3(new_n1119), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1061), .A2(new_n1066), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT62), .B1(new_n1121), .B2(new_n1064), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1006), .A2(new_n1022), .A3(new_n1042), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1067), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .A4(new_n1114), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n997), .B(KEYINPUT117), .ZN(new_n1127));
  OR3_X1    g702(.A1(new_n998), .A2(G1976), .A3(G288), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1127), .B1(new_n1128), .B2(new_n989), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1010), .B2(new_n1023), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1046), .A2(new_n1120), .A3(new_n1126), .A4(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT127), .ZN(new_n1132));
  XNOR2_X1  g707(.A(G290), .B(G1986), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n984), .B1(new_n973), .B2(new_n1133), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1132), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n988), .B1(new_n1135), .B2(new_n1136), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g712(.A1(G229), .A2(new_n464), .A3(G401), .A4(G227), .ZN(new_n1139));
  NAND3_X1  g713(.A1(new_n942), .A2(new_n876), .A3(new_n1139), .ZN(G225));
  INV_X1    g714(.A(G225), .ZN(G308));
endmodule


