//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n208), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  INV_X1    g0016(.A(new_n201), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(KEYINPUT64), .ZN(new_n219));
  AND3_X1   g0019(.A1(new_n218), .A2(G50), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n208), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n216), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n215), .ZN(G361));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT65), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n233), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G58), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G1698), .ZN(new_n247));
  AND2_X1   g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NOR2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  OAI211_X1 g0049(.A(G223), .B(new_n247), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT77), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n252), .A2(new_n253), .A3(G223), .A4(new_n247), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G87), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n252), .A2(G226), .A3(G1698), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n251), .A2(new_n254), .A3(new_n255), .A4(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT67), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  AND4_X1   g0059(.A1(new_n258), .A2(new_n259), .A3(G1), .A4(G13), .ZN(new_n260));
  AND2_X1   g0060(.A1(G1), .A2(G13), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n258), .B1(new_n261), .B2(new_n259), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G179), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(new_n269), .A3(G274), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n267), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(new_n235), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n264), .A2(new_n265), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT78), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT8), .B(G58), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n276), .B1(new_n266), .B2(G20), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n221), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n277), .A2(new_n282), .B1(new_n279), .B2(new_n276), .ZN(new_n283));
  XNOR2_X1  g0083(.A(G58), .B(G68), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n284), .A2(G20), .B1(G159), .B2(new_n285), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n248), .A2(new_n249), .A3(G20), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT7), .ZN(new_n288));
  OAI21_X1  g0088(.A(G68), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OR2_X1    g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n222), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n288), .A2(KEYINPUT76), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT76), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT7), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(KEYINPUT16), .B(new_n286), .C1(new_n289), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n281), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n290), .A2(KEYINPUT7), .A3(new_n222), .A4(new_n291), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n287), .B2(new_n296), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G68), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT16), .B1(new_n302), .B2(new_n286), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n283), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n264), .A2(new_n273), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n272), .B1(new_n257), .B2(new_n263), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT78), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(new_n309), .A3(new_n265), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n275), .A2(new_n304), .A3(new_n307), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT18), .ZN(new_n312));
  AOI211_X1 g0112(.A(G179), .B(new_n272), .C1(new_n257), .C2(new_n263), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n313), .A2(new_n309), .B1(new_n305), .B2(new_n306), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT18), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n314), .A2(new_n315), .A3(new_n304), .A4(new_n275), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT17), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT79), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n264), .A2(G190), .A3(new_n273), .ZN(new_n320));
  INV_X1    g0120(.A(G200), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n308), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n319), .B1(new_n322), .B2(new_n304), .ZN(new_n323));
  INV_X1    g0123(.A(new_n283), .ZN(new_n324));
  INV_X1    g0124(.A(new_n281), .ZN(new_n325));
  INV_X1    g0125(.A(G58), .ZN(new_n326));
  INV_X1    g0126(.A(G68), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(G20), .B1(new_n328), .B2(new_n201), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n285), .A2(G159), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n293), .A2(new_n295), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n287), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n327), .B1(new_n292), .B2(KEYINPUT7), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n325), .B1(new_n335), .B2(KEYINPUT16), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT16), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n332), .A2(new_n292), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n327), .B1(new_n338), .B2(new_n300), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n337), .B1(new_n339), .B2(new_n331), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n324), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n305), .A2(G200), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n341), .A2(KEYINPUT79), .A3(new_n320), .A4(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n318), .B1(new_n323), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n322), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT17), .B1(new_n345), .B2(new_n341), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n317), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n325), .A2(new_n278), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n266), .A2(G20), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G50), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n348), .A2(new_n350), .B1(G50), .B2(new_n278), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT70), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n276), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n222), .A2(G33), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT68), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G33), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(G20), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT68), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n354), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n285), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n325), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(KEYINPUT69), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n363), .A2(KEYINPUT69), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n353), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n252), .A2(G222), .A3(new_n247), .ZN(new_n367));
  INV_X1    g0167(.A(G77), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n252), .A2(G1698), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT66), .B(G223), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n367), .B1(new_n368), .B2(new_n252), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n263), .ZN(new_n372));
  INV_X1    g0172(.A(new_n270), .ZN(new_n373));
  INV_X1    g0173(.A(new_n271), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n373), .B1(G226), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(new_n265), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n372), .A2(new_n375), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n306), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n366), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT9), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n366), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT72), .ZN(new_n382));
  INV_X1    g0182(.A(G190), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n372), .A2(KEYINPUT72), .A3(G190), .A4(new_n375), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n353), .B(KEYINPUT9), .C1(new_n364), .C2(new_n365), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n377), .A2(G200), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n381), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT10), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n387), .A2(new_n388), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT10), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n391), .A2(new_n392), .A3(new_n386), .A4(new_n381), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n379), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n360), .A2(G77), .A3(new_n357), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n285), .A2(G50), .B1(G20), .B2(new_n327), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n281), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT11), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT11), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(new_n400), .A3(new_n281), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n266), .A2(new_n327), .A3(G13), .A4(G20), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT12), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n325), .A2(G68), .A3(new_n278), .A4(new_n349), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT75), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT75), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n399), .A2(new_n401), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n270), .A2(KEYINPUT74), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G97), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT73), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(G226), .A2(G1698), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n235), .B2(G1698), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n415), .B1(new_n252), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n269), .A2(KEYINPUT67), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n261), .A2(new_n258), .A3(new_n259), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n410), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT74), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n268), .A2(new_n269), .A3(new_n423), .A4(G274), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n269), .A2(G238), .A3(new_n267), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT13), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(KEYINPUT73), .A2(G33), .A3(G97), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT73), .B1(G33), .B2(G97), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n235), .A2(G1698), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(G226), .B2(G1698), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n248), .A2(new_n249), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n434), .A2(new_n263), .B1(KEYINPUT74), .B2(new_n270), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT13), .ZN(new_n436));
  INV_X1    g0236(.A(new_n426), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n427), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n409), .B1(new_n439), .B2(new_n383), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n321), .B1(new_n427), .B2(new_n438), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n422), .A2(KEYINPUT13), .A3(new_n426), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n436), .B1(new_n435), .B2(new_n437), .ZN(new_n444));
  OAI21_X1  g0244(.A(G169), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT14), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n427), .A2(G179), .A3(new_n438), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT14), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n448), .B(G169), .C1(new_n443), .C2(new_n444), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n409), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n442), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT71), .ZN(new_n453));
  INV_X1    g0253(.A(G244), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n270), .B1(new_n454), .B2(new_n271), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n252), .A2(G232), .A3(new_n247), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n252), .A2(G238), .A3(G1698), .ZN(new_n457));
  INV_X1    g0257(.A(G107), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n252), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n455), .B1(new_n459), .B2(new_n263), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(G169), .ZN(new_n461));
  INV_X1    g0261(.A(new_n285), .ZN(new_n462));
  OAI22_X1  g0262(.A1(new_n276), .A2(new_n462), .B1(new_n222), .B2(new_n368), .ZN(new_n463));
  XNOR2_X1  g0263(.A(KEYINPUT15), .B(G87), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(new_n355), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n281), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n279), .A2(new_n368), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n282), .A2(G77), .A3(new_n349), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n453), .B1(new_n461), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n460), .A2(new_n265), .ZN(new_n472));
  OAI211_X1 g0272(.A(KEYINPUT71), .B(new_n469), .C1(new_n460), .C2(G169), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n459), .A2(new_n263), .ZN(new_n475));
  INV_X1    g0275(.A(new_n455), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n469), .B1(new_n477), .B2(G200), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n383), .B2(new_n477), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  AND4_X1   g0280(.A1(new_n347), .A2(new_n394), .A3(new_n452), .A4(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT82), .ZN(new_n482));
  AOI21_X1  g0282(.A(G20), .B1(new_n290), .B2(new_n291), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G68), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT19), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n485), .B1(new_n355), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT19), .B1(new_n428), .B2(new_n429), .ZN(new_n489));
  INV_X1    g0289(.A(G87), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n489), .A2(new_n222), .B1(new_n490), .B2(new_n205), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n482), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n485), .B1(new_n413), .B2(new_n414), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n493), .A2(G20), .B1(G87), .B2(new_n206), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n494), .A2(KEYINPUT82), .A3(new_n484), .A4(new_n487), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n492), .A2(new_n495), .A3(new_n281), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n464), .A2(new_n279), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n348), .B1(new_n266), .B2(G33), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G87), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G45), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(G1), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n269), .A2(G274), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n266), .A2(G45), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n269), .A2(G250), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(G244), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n507));
  OAI211_X1 g0307(.A(G238), .B(new_n247), .C1(new_n248), .C2(new_n249), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G116), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n506), .B1(new_n263), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n383), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(G200), .B2(new_n511), .ZN(new_n513));
  INV_X1    g0313(.A(new_n464), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n498), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n496), .A2(new_n515), .A3(new_n497), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n511), .A2(G179), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n306), .B2(new_n511), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n500), .A2(new_n513), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT6), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n520), .A2(new_n486), .A3(G107), .ZN(new_n521));
  XNOR2_X1  g0321(.A(G97), .B(G107), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n521), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  OAI22_X1  g0323(.A1(new_n523), .A2(new_n222), .B1(new_n368), .B2(new_n462), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n458), .B1(new_n338), .B2(new_n300), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n281), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n278), .A2(G97), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(new_n498), .B2(G97), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G244), .B(new_n247), .C1(new_n248), .C2(new_n249), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT4), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G250), .A2(G1698), .ZN(new_n533));
  NAND2_X1  g0333(.A1(KEYINPUT4), .A2(G244), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(G1698), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n252), .A2(new_n535), .B1(G33), .B2(G283), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n263), .ZN(new_n538));
  AND2_X1   g0338(.A1(KEYINPUT5), .A2(G41), .ZN(new_n539));
  NOR2_X1   g0339(.A1(KEYINPUT5), .A2(G41), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n502), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(G257), .A3(new_n269), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n269), .A2(G274), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n540), .ZN(new_n545));
  NAND2_X1  g0345(.A1(KEYINPUT5), .A2(G41), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n504), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n542), .A2(KEYINPUT80), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT80), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n541), .A2(new_n549), .A3(G257), .A4(new_n269), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n538), .A2(new_n265), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n542), .A2(KEYINPUT80), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n544), .A2(new_n547), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n421), .B1(new_n532), .B2(new_n536), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n306), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n529), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n321), .B1(new_n554), .B2(new_n555), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n538), .A2(new_n548), .A3(new_n383), .A4(new_n550), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n526), .A2(new_n528), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT81), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n562), .B1(new_n560), .B2(new_n561), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n519), .B(new_n557), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n282), .B(G116), .C1(G1), .C2(new_n358), .ZN(new_n567));
  INV_X1    g0367(.A(G116), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n279), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n280), .A2(new_n221), .B1(G20), .B2(new_n568), .ZN(new_n570));
  AOI21_X1  g0370(.A(G20), .B1(G33), .B2(G283), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(G33), .B2(new_n486), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT20), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n570), .A2(new_n572), .A3(KEYINPUT20), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n567), .B(new_n569), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT21), .ZN(new_n576));
  XNOR2_X1  g0376(.A(KEYINPUT5), .B(G41), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(new_n502), .B1(new_n261), .B2(new_n259), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(G270), .B1(new_n544), .B2(new_n547), .ZN(new_n579));
  OAI211_X1 g0379(.A(G264), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n580));
  OAI211_X1 g0380(.A(G257), .B(new_n247), .C1(new_n248), .C2(new_n249), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n290), .A2(G303), .A3(new_n291), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n263), .ZN(new_n584));
  AOI211_X1 g0384(.A(new_n576), .B(new_n306), .C1(new_n579), .C2(new_n584), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n579), .A2(G179), .A3(new_n584), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n575), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n579), .A2(new_n584), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n575), .A2(new_n588), .A3(G169), .ZN(new_n589));
  XOR2_X1   g0389(.A(KEYINPUT83), .B(KEYINPUT21), .Z(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(G200), .ZN(new_n594));
  INV_X1    g0394(.A(new_n575), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n594), .B(new_n595), .C1(new_n383), .C2(new_n588), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(G257), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n598));
  OAI211_X1 g0398(.A(G250), .B(new_n247), .C1(new_n248), .C2(new_n249), .ZN(new_n599));
  AND2_X1   g0399(.A1(KEYINPUT87), .A2(G294), .ZN(new_n600));
  NOR2_X1   g0400(.A1(KEYINPUT87), .A2(G294), .ZN(new_n601));
  OAI21_X1  g0401(.A(G33), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n598), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n603), .A2(new_n263), .B1(new_n578), .B2(G264), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n553), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT88), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT88), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n604), .A2(new_n607), .A3(new_n553), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(G169), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT89), .B1(new_n605), .B2(new_n265), .ZN(new_n610));
  INV_X1    g0410(.A(new_n605), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT89), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n612), .A3(G179), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT24), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n222), .B(G87), .C1(new_n248), .C2(new_n249), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT22), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT84), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT85), .B1(new_n616), .B2(KEYINPUT22), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT22), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n483), .A2(new_n622), .A3(new_n623), .A4(G87), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n619), .A2(new_n620), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n458), .A2(KEYINPUT23), .A3(G20), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT23), .B1(new_n458), .B2(G20), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n627), .A2(new_n628), .B1(G20), .B2(new_n509), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n615), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n629), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n621), .A2(new_n624), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n616), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT84), .B1(new_n616), .B2(KEYINPUT22), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(KEYINPUT24), .B(new_n631), .C1(new_n632), .C2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n630), .A2(new_n636), .A3(new_n281), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n279), .A2(new_n458), .ZN(new_n638));
  NOR2_X1   g0438(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n638), .B2(new_n639), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n498), .A2(G107), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n614), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(G190), .B1(new_n606), .B2(new_n608), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n611), .A2(G200), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n637), .B(new_n643), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n481), .A2(new_n566), .A3(new_n597), .A4(new_n649), .ZN(G372));
  NAND4_X1  g0450(.A1(new_n513), .A2(new_n497), .A3(new_n496), .A4(new_n499), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n511), .A2(new_n306), .ZN(new_n652));
  AOI211_X1 g0452(.A(new_n265), .B(new_n506), .C1(new_n263), .C2(new_n510), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT90), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT90), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n517), .B(new_n655), .C1(new_n306), .C2(new_n511), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n654), .A2(new_n516), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n648), .A2(new_n651), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n592), .B1(new_n644), .B2(new_n614), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n557), .B1(new_n563), .B2(new_n564), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n557), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n516), .A2(new_n518), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n663), .A3(new_n651), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT26), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n657), .A2(new_n662), .A3(new_n666), .A4(new_n651), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n665), .A2(new_n657), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n481), .B1(new_n661), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n669), .B(KEYINPUT91), .Z(new_n670));
  NAND2_X1  g0470(.A1(new_n449), .A2(new_n447), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n448), .B1(new_n439), .B2(G169), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n451), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n477), .A2(new_n306), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT71), .B1(new_n674), .B2(new_n469), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n473), .A2(new_n472), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT92), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT92), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n471), .A2(new_n678), .A3(new_n472), .A4(new_n473), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n673), .B1(new_n680), .B2(new_n442), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n323), .A2(new_n343), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n346), .B1(new_n682), .B2(KEYINPUT17), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n312), .A2(new_n316), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n390), .A2(new_n393), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n379), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n670), .A2(new_n688), .ZN(G369));
  NAND3_X1  g0489(.A1(new_n266), .A2(new_n222), .A3(G13), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G213), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(KEYINPUT27), .B2(new_n690), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n595), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT93), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n597), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n593), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n694), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n644), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n649), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n645), .B2(new_n694), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n645), .A2(new_n701), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n592), .A2(new_n694), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT94), .Z(new_n708));
  AOI21_X1  g0508(.A(new_n706), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n705), .A2(new_n709), .ZN(G399));
  NOR3_X1   g0510(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n711));
  INV_X1    g0511(.A(G41), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n225), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(new_n713), .A3(G1), .ZN(new_n714));
  INV_X1    g0514(.A(new_n220), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT95), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n660), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n659), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n648), .A2(new_n651), .A3(new_n657), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT95), .B(new_n557), .C1(new_n563), .C2(new_n564), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n719), .A2(new_n720), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n657), .A2(new_n651), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n666), .B1(new_n724), .B2(new_n662), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n657), .B1(new_n664), .B2(KEYINPUT26), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .A3(new_n694), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n661), .A2(new_n668), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n730), .B1(new_n731), .B2(new_n701), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n511), .A2(new_n604), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n554), .A2(new_n555), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(new_n586), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n734), .A2(new_n735), .A3(new_n586), .A4(KEYINPUT30), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n538), .A2(new_n550), .A3(new_n548), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n511), .A2(G179), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(new_n741), .A3(new_n588), .A4(new_n605), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n738), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n744));
  AND4_X1   g0544(.A1(new_n587), .A2(new_n596), .A3(new_n591), .A4(new_n694), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(new_n645), .A3(new_n648), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n744), .B1(new_n746), .B2(new_n565), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT31), .B1(new_n743), .B2(new_n701), .ZN(new_n748));
  OAI21_X1  g0548(.A(G330), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n733), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n717), .B1(new_n751), .B2(G1), .ZN(G364));
  AND2_X1   g0552(.A1(new_n222), .A2(G13), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n266), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n713), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n700), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G330), .B2(new_n698), .ZN(new_n759));
  INV_X1    g0559(.A(G355), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n252), .A2(new_n225), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n761), .B1(G116), .B2(new_n225), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n242), .A2(new_n501), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n433), .A2(new_n225), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n220), .B2(new_n501), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n221), .B1(G20), .B2(new_n306), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n757), .B1(new_n766), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n222), .A2(new_n265), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G190), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n222), .A2(G179), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(new_n383), .A3(G200), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n777), .A2(new_n327), .B1(new_n458), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n775), .A2(new_n383), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n782), .A2(new_n202), .B1(new_n490), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n774), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n774), .A2(G190), .A3(new_n321), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n252), .B1(new_n786), .B2(new_n368), .C1(new_n326), .C2(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n780), .A2(new_n784), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n265), .A2(new_n321), .A3(G190), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n486), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n778), .A2(new_n785), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G159), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n793), .B1(KEYINPUT32), .B2(new_n796), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n789), .B(new_n797), .C1(KEYINPUT32), .C2(new_n796), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n783), .B(KEYINPUT96), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G303), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n781), .A2(G326), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n600), .A2(new_n601), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n804), .B2(new_n792), .ZN(new_n805));
  INV_X1    g0605(.A(new_n779), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(G283), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(KEYINPUT33), .B(G317), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n809), .A2(KEYINPUT97), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(KEYINPUT97), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n810), .A2(new_n776), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n786), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n252), .B1(new_n813), .B2(G311), .ZN(new_n814));
  INV_X1    g0614(.A(new_n787), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(G322), .B1(new_n795), .B2(G329), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n807), .A2(new_n812), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n798), .B1(new_n802), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT98), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n770), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n818), .B2(new_n819), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n773), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n769), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n698), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n759), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  NAND4_X1  g0627(.A1(new_n677), .A2(new_n679), .A3(new_n469), .A4(new_n701), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n474), .B(new_n479), .C1(new_n470), .C2(new_n694), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n731), .B2(new_n701), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n694), .B(new_n830), .C1(new_n661), .C2(new_n668), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n757), .B1(new_n834), .B2(new_n749), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n749), .B2(new_n834), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n770), .A2(new_n767), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n757), .B1(G77), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n815), .A2(G143), .B1(new_n813), .B2(G159), .ZN(new_n840));
  INV_X1    g0640(.A(G137), .ZN(new_n841));
  INV_X1    g0641(.A(G150), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n840), .B1(new_n782), .B2(new_n841), .C1(new_n842), .C2(new_n777), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT34), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n799), .A2(G50), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n252), .B1(new_n794), .B2(new_n848), .C1(new_n779), .C2(new_n327), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G58), .B2(new_n791), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n850), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n782), .A2(new_n801), .B1(new_n786), .B2(new_n568), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n776), .A2(KEYINPUT99), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n776), .A2(KEYINPUT99), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n852), .B1(new_n856), .B2(G283), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT100), .Z(new_n858));
  AOI211_X1 g0658(.A(new_n252), .B(new_n793), .C1(G294), .C2(new_n815), .ZN(new_n859));
  INV_X1    g0659(.A(G311), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n779), .A2(new_n490), .B1(new_n794), .B2(new_n860), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT101), .Z(new_n862));
  OAI211_X1 g0662(.A(new_n859), .B(new_n862), .C1(new_n458), .C2(new_n800), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n851), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n839), .B1(new_n864), .B2(new_n770), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n768), .B2(new_n830), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n836), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(G384));
  XNOR2_X1  g0668(.A(new_n523), .B(KEYINPUT102), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT35), .ZN(new_n870));
  OAI211_X1 g0670(.A(G116), .B(new_n223), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n870), .B2(new_n869), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT36), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n715), .A2(new_n368), .A3(new_n328), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n874), .A2(KEYINPUT103), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n874), .A2(KEYINPUT103), .B1(new_n202), .B2(G68), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n266), .B(G13), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n451), .B(new_n701), .C1(new_n450), .C2(new_n442), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n440), .A2(new_n441), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n451), .A2(new_n701), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n673), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n879), .A2(new_n882), .B1(new_n828), .B2(new_n829), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT105), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n743), .A2(new_n884), .A3(new_n701), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n884), .B1(new_n743), .B2(new_n701), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT31), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n883), .B1(new_n887), .B2(new_n747), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT106), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n334), .A2(new_n333), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT16), .B1(new_n892), .B2(new_n286), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n283), .B1(new_n299), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n693), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n683), .B2(new_n685), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n275), .A2(new_n894), .A3(new_n307), .A4(new_n310), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n323), .A2(new_n343), .A3(new_n897), .A4(new_n895), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n323), .A2(new_n343), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT37), .B1(new_n304), .B2(new_n693), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n311), .A2(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(KEYINPUT37), .A2(new_n898), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n891), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n898), .A2(KEYINPUT37), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n899), .A2(new_n901), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n906), .B(KEYINPUT38), .C1(new_n347), .C2(new_n895), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n883), .B(KEYINPUT106), .C1(new_n887), .C2(new_n747), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n890), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n304), .A2(new_n693), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n683), .B2(new_n685), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n311), .B(new_n913), .C1(new_n304), .C2(new_n322), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n901), .A2(new_n899), .B1(new_n915), .B2(KEYINPUT37), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n891), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n917), .A2(new_n907), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n883), .B(KEYINPUT40), .C1(new_n887), .C2(new_n747), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n912), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n887), .A2(new_n747), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n481), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(G330), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n920), .B2(new_n922), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n450), .A2(new_n451), .A3(new_n694), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n927));
  AND3_X1   g0727(.A1(new_n917), .A2(new_n907), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT39), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n903), .B2(new_n907), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n926), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n879), .A2(new_n882), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n474), .A2(new_n701), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n932), .B1(new_n833), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n908), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n685), .A2(new_n693), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n931), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n729), .A2(new_n732), .A3(new_n481), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n940), .A2(new_n688), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n939), .B(new_n941), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n924), .A2(new_n942), .B1(new_n266), .B2(new_n753), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n924), .A2(new_n942), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n878), .B1(new_n943), .B2(new_n944), .ZN(G367));
  AND3_X1   g0745(.A1(new_n233), .A2(new_n225), .A3(new_n433), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n771), .B1(new_n225), .B2(new_n464), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n757), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n856), .A2(G159), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n787), .A2(new_n842), .B1(new_n794), .B2(new_n841), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n433), .B(new_n950), .C1(G50), .C2(new_n813), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n781), .A2(G143), .B1(G68), .B2(new_n791), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n779), .A2(new_n368), .ZN(new_n953));
  INV_X1    g0753(.A(new_n783), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n953), .B1(G58), .B2(new_n954), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n949), .A2(new_n951), .A3(new_n952), .A4(new_n955), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n782), .A2(new_n860), .B1(new_n779), .B2(new_n486), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(G107), .B2(new_n791), .ZN(new_n958));
  INV_X1    g0758(.A(G317), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n787), .A2(new_n801), .B1(new_n794), .B2(new_n959), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n252), .B(new_n960), .C1(G283), .C2(new_n813), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n783), .A2(new_n568), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n958), .B(new_n961), .C1(KEYINPUT46), .C2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n799), .A2(KEYINPUT46), .A3(G116), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n855), .B2(new_n804), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n956), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT47), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n948), .B1(new_n967), .B2(new_n770), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n500), .A2(new_n694), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n724), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n657), .B2(new_n969), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n968), .B1(new_n824), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n719), .B(new_n722), .C1(new_n561), .C2(new_n694), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n662), .A2(new_n701), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT107), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n709), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(KEYINPUT110), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT110), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n709), .A2(new_n979), .A3(new_n976), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n709), .A2(new_n976), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT44), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n978), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT111), .ZN(new_n988));
  INV_X1    g0788(.A(new_n705), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n983), .A2(new_n985), .A3(new_n705), .A4(new_n986), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n704), .A2(new_n708), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(KEYINPUT112), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n700), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(KEYINPUT112), .A3(new_n699), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n704), .B2(new_n708), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n704), .A2(new_n708), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n995), .A2(new_n999), .A3(new_n996), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n750), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n705), .A2(KEYINPUT111), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n992), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n751), .B1(new_n991), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n713), .B(KEYINPUT41), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n755), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n989), .A2(new_n976), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT109), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n973), .A2(new_n975), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n557), .B1(new_n1010), .B2(new_n645), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n694), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT42), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n993), .A2(new_n1010), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT108), .ZN(new_n1015));
  NOR4_X1   g0815(.A1(new_n993), .A2(new_n1010), .A3(new_n1015), .A4(KEYINPUT42), .ZN(new_n1016));
  AOI21_X1  g0816(.A(KEYINPUT108), .B1(new_n1014), .B2(new_n1013), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1009), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1009), .A2(new_n1019), .A3(new_n1018), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1023), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1025), .A2(new_n1020), .B1(KEYINPUT43), .B2(new_n971), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n972), .B1(new_n1007), .B2(new_n1027), .ZN(G387));
  NOR2_X1   g0828(.A1(new_n1001), .A2(new_n713), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n998), .A2(new_n1000), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1029), .B1(new_n751), .B2(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n704), .A2(new_n824), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n711), .A2(new_n761), .B1(G107), .B2(new_n225), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n711), .ZN(new_n1034));
  AOI211_X1 g0834(.A(G45), .B(new_n1034), .C1(G68), .C2(G77), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n276), .A2(G50), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT50), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n764), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n238), .A2(G45), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1033), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n757), .B1(new_n1040), .B2(new_n772), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n786), .A2(new_n327), .B1(new_n794), .B2(new_n842), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n433), .B(new_n1042), .C1(G50), .C2(new_n815), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n954), .A2(G77), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n792), .A2(new_n464), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n354), .B2(new_n776), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n781), .A2(G159), .B1(new_n806), .B2(G97), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n252), .B1(new_n795), .B2(G326), .ZN(new_n1049));
  INV_X1    g0849(.A(G283), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n792), .A2(new_n1050), .B1(new_n804), .B2(new_n783), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT113), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n787), .A2(new_n959), .B1(new_n786), .B2(new_n801), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G322), .B2(new_n781), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n855), .B2(new_n860), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT48), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1052), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT49), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1049), .B1(new_n568), .B2(new_n779), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1048), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT114), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n821), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1041), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1030), .A2(new_n755), .B1(new_n1032), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1031), .A2(new_n1067), .ZN(G393));
  NAND2_X1  g0868(.A1(new_n987), .A2(new_n989), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1069), .A2(new_n992), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1070), .A2(new_n1001), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1003), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n713), .B1(new_n1072), .B2(new_n990), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1069), .A2(new_n755), .A3(new_n992), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n771), .B1(new_n486), .B2(new_n225), .C1(new_n245), .C2(new_n764), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n757), .ZN(new_n1077));
  INV_X1    g0877(.A(G159), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n782), .A2(new_n842), .B1(new_n1078), .B2(new_n787), .ZN(new_n1079));
  XOR2_X1   g0879(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n856), .A2(G50), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n792), .A2(new_n368), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n327), .B2(new_n783), .C1(new_n490), .C2(new_n779), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n433), .B1(new_n795), .B2(G143), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n276), .B2(new_n786), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1082), .B(new_n1088), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G317), .A2(new_n781), .B1(new_n815), .B2(G311), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n795), .A2(G322), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n252), .B(new_n1092), .C1(G294), .C2(new_n813), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n458), .A2(new_n779), .B1(new_n783), .B2(new_n1050), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G116), .B2(new_n791), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(new_n855), .C2(new_n801), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1089), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1077), .B1(new_n1097), .B2(new_n770), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n976), .B2(new_n824), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1075), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT116), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1075), .A2(KEYINPUT116), .A3(new_n1099), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1074), .A2(new_n1104), .ZN(G390));
  NAND3_X1  g0905(.A1(new_n481), .A2(new_n921), .A3(G330), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n940), .A2(new_n688), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n833), .A2(new_n934), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n921), .A2(G330), .A3(new_n883), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(G330), .B(new_n830), .C1(new_n747), .C2(new_n748), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1111), .A2(new_n932), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1108), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1111), .A2(new_n932), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n701), .B1(new_n723), .B2(new_n727), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n933), .B1(new_n1115), .B2(new_n830), .ZN(new_n1116));
  OAI211_X1 g0916(.A(G330), .B(new_n830), .C1(new_n887), .C2(new_n747), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n932), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1107), .B1(new_n1113), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n908), .A2(KEYINPUT39), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n917), .A2(new_n907), .A3(new_n927), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1122), .B(new_n1123), .C1(new_n935), .C2(new_n926), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n926), .B1(new_n917), .B2(new_n907), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n1116), .B2(new_n932), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1124), .A2(new_n1126), .A3(new_n1114), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1109), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1121), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n935), .A2(new_n926), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1126), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1110), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1124), .A2(new_n1126), .A3(new_n1114), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n1120), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1129), .A2(new_n756), .A3(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1122), .A2(new_n767), .A3(new_n1123), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n757), .B1(new_n354), .B2(new_n838), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT117), .Z(new_n1140));
  OAI221_X1 g0940(.A(new_n1084), .B1(new_n327), .B2(new_n779), .C1(new_n1050), .C2(new_n782), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(G97), .A2(new_n813), .B1(new_n795), .B2(G294), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1142), .B(new_n433), .C1(new_n568), .C2(new_n787), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n855), .A2(new_n458), .B1(new_n490), .B2(new_n800), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n781), .A2(G128), .B1(new_n806), .B2(G50), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n1078), .B2(new_n792), .C1(new_n855), .C2(new_n841), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n783), .A2(new_n842), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT53), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n252), .B1(new_n787), .B2(new_n848), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G125), .B2(new_n795), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT54), .B(G143), .Z(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT118), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1149), .B(new_n1151), .C1(new_n1154), .C2(new_n786), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1144), .A2(new_n1145), .B1(new_n1147), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1140), .B1(new_n1156), .B2(new_n770), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT119), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1137), .A2(new_n755), .B1(new_n1138), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1136), .A2(new_n1159), .ZN(G378));
  NAND2_X1  g0960(.A1(new_n1113), .A2(new_n1119), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1107), .B1(new_n1137), .B2(new_n1161), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n931), .A2(new_n936), .A3(new_n938), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1163), .A2(KEYINPUT122), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n889), .A2(new_n888), .B1(new_n903), .B2(new_n907), .ZN(new_n1166));
  AOI21_X1  g0966(.A(KEYINPUT40), .B1(new_n1166), .B2(new_n909), .ZN(new_n1167));
  OAI21_X1  g0967(.A(G330), .B1(new_n918), .B2(new_n919), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n366), .A2(new_n693), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n394), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n394), .A2(new_n1171), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1170), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n394), .A2(new_n1171), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1176), .A2(new_n1172), .A3(new_n1169), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1167), .A2(new_n1168), .A3(new_n1178), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1180));
  INV_X1    g0980(.A(G330), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n919), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n917), .A2(new_n907), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1180), .B1(new_n912), .B2(new_n1184), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1179), .A2(new_n1185), .A3(KEYINPUT123), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT123), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1178), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n912), .A2(new_n1184), .A3(new_n1180), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1165), .B1(new_n1186), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(KEYINPUT123), .B1(new_n1179), .B2(new_n1185), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1188), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1192), .A2(new_n1164), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1162), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(KEYINPUT125), .B1(new_n1195), .B2(KEYINPUT57), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n939), .B1(new_n1179), .B2(new_n1185), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1163), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1197), .A2(KEYINPUT57), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(KEYINPUT124), .B1(new_n1162), .B2(new_n1199), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1179), .A2(new_n1185), .A3(new_n939), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n937), .B1(new_n1130), .B2(new_n926), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1188), .A2(new_n1189), .B1(new_n1202), .B2(new_n936), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT124), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1107), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1135), .A2(new_n1206), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1207), .A4(KEYINPUT57), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n713), .B1(new_n1200), .B2(new_n1208), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1192), .A2(new_n1164), .A3(new_n1193), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1164), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1207), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT125), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT57), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1196), .A2(new_n1209), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n754), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1180), .A2(new_n767), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n757), .B1(G50), .B2(new_n838), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT121), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(G33), .A2(G41), .ZN(new_n1221));
  AOI211_X1 g1021(.A(G50), .B(new_n1221), .C1(new_n433), .C2(new_n712), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n779), .A2(new_n326), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G116), .B2(new_n781), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n486), .B2(new_n777), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n433), .B(new_n712), .C1(new_n794), .C2(new_n1050), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n787), .A2(new_n458), .B1(new_n786), .B2(new_n464), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1044), .B1(new_n327), .B2(new_n792), .ZN(new_n1228));
  OR4_X1    g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT58), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1222), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(G128), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n787), .A2(new_n1232), .B1(new_n786), .B2(new_n841), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G132), .B2(new_n776), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n781), .A2(G125), .B1(G150), .B2(new_n791), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(new_n1154), .C2(new_n783), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(KEYINPUT59), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(KEYINPUT59), .ZN(new_n1238));
  INV_X1    g1038(.A(G124), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1221), .B1(new_n794), .B2(new_n1239), .C1(new_n779), .C2(new_n1078), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT120), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1238), .A2(new_n1241), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1231), .B1(new_n1230), .B2(new_n1229), .C1(new_n1237), .C2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1220), .B1(new_n1243), .B2(new_n770), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1217), .B1(new_n1218), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1216), .A2(new_n1245), .ZN(G375));
  NAND3_X1  g1046(.A1(new_n1113), .A2(new_n1107), .A3(new_n1119), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1121), .A2(new_n1006), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n932), .A2(new_n767), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n757), .B1(G68), .B2(new_n838), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n856), .A2(G116), .B1(G97), .B2(new_n799), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n786), .A2(new_n458), .B1(new_n794), .B2(new_n801), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n252), .B(new_n1252), .C1(G283), .C2(new_n815), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n953), .B(new_n1045), .C1(G294), .C2(new_n781), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1251), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n856), .A2(new_n1153), .B1(G159), .B2(new_n799), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n786), .A2(new_n842), .B1(new_n794), .B2(new_n1232), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n433), .B(new_n1257), .C1(G137), .C2(new_n815), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n792), .A2(new_n202), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1223), .B(new_n1259), .C1(G132), .C2(new_n781), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1256), .A2(new_n1258), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1255), .A2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1250), .B1(new_n1262), .B2(new_n770), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1161), .A2(new_n755), .B1(new_n1249), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1248), .A2(new_n1264), .ZN(G381));
  NAND3_X1  g1065(.A1(new_n1031), .A2(new_n826), .A3(new_n1067), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n867), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1264), .B(new_n1248), .C1(new_n1268), .C2(KEYINPUT126), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(KEYINPUT126), .B2(new_n1268), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1071), .A2(new_n1073), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1271));
  INV_X1    g1071(.A(G378), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  OR3_X1    g1073(.A1(new_n1273), .A2(G387), .A3(G375), .ZN(G407));
  INV_X1    g1074(.A(G343), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(G213), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1272), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G407), .B(G213), .C1(G375), .C2(new_n1278), .ZN(G409));
  INV_X1    g1079(.A(KEYINPUT63), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1216), .A2(G378), .A3(new_n1245), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1218), .A2(new_n1244), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1204), .A2(new_n755), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1282), .B(new_n1283), .C1(new_n1212), .C2(new_n1005), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1272), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1276), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT60), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1247), .B1(new_n1120), .B2(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1113), .A2(new_n1107), .A3(KEYINPUT60), .A4(new_n1119), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1289), .A2(new_n756), .A3(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(G384), .A3(new_n1264), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(G384), .B1(new_n1291), .B2(new_n1264), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1280), .B1(new_n1287), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1277), .A2(G2897), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT61), .B1(new_n1287), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G393), .A2(G396), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT127), .B1(new_n1303), .B2(new_n1266), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(G387), .B2(G390), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1271), .B(new_n972), .C1(new_n1007), .C2(new_n1027), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1303), .A2(KEYINPUT127), .A3(new_n1266), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1305), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1307), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1277), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1311), .A2(KEYINPUT63), .A3(new_n1295), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1297), .A2(new_n1302), .A3(new_n1310), .A4(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1311), .A2(new_n1314), .A3(new_n1295), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1301), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1316), .B1(new_n1311), .B2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1314), .B1(new_n1311), .B2(new_n1295), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1315), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1313), .B1(new_n1320), .B2(new_n1310), .ZN(G405));
  INV_X1    g1121(.A(new_n1310), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(G375), .A2(new_n1272), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1281), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1295), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1323), .A2(new_n1296), .A3(new_n1281), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1322), .B(new_n1327), .ZN(G402));
endmodule


